--Copyright (C)2014-2024 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--Tool Version: V1.9.9.01 (64-bit)
--Part Number: GW2AR-LV18QN88C8/I7
--Device: GW2AR-18
--Device Version: C
--Created Time: Wed Feb 28 23:50:26 2024

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM_basic is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(12 downto 0)
    );
end Gowin_pROM_basic;

architecture Behavioral of Gowin_pROM_basic is

    signal prom_inst_0_dout_w: std_logic_vector(29 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(29 downto 0);
    signal prom_inst_2_dout_w: std_logic_vector(29 downto 0);
    signal prom_inst_3_dout_w: std_logic_vector(29 downto 0);
    signal gw_gnd: std_logic;
    signal prom_inst_0_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_2_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_2_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_3_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_3_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 1;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    gw_gnd <= '0';

    prom_inst_0_AD_i <= ad(12 downto 0) & gw_gnd;
    dout(1 downto 0) <= prom_inst_0_DO_o(1 downto 0) ;
    prom_inst_0_dout_w(29 downto 0) <= prom_inst_0_DO_o(31 downto 2) ;
    prom_inst_1_AD_i <= ad(12 downto 0) & gw_gnd;
    dout(3 downto 2) <= prom_inst_1_DO_o(1 downto 0) ;
    prom_inst_1_dout_w(29 downto 0) <= prom_inst_1_DO_o(31 downto 2) ;
    prom_inst_2_AD_i <= ad(12 downto 0) & gw_gnd;
    dout(5 downto 4) <= prom_inst_2_DO_o(1 downto 0) ;
    prom_inst_2_dout_w(29 downto 0) <= prom_inst_2_DO_o(31 downto 2) ;
    prom_inst_3_AD_i <= ad(12 downto 0) & gw_gnd;
    dout(7 downto 6) <= prom_inst_3_DO_o(1 downto 0) ;
    prom_inst_3_dout_w(29 downto 0) <= prom_inst_3_DO_o(31 downto 2) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"FCC8FD1C1F989D60DED00019E76699B2BB3E5640626120703410EC35D0DD9B3C",
            INIT_RAM_01 => X"87C919999C705ECCD6A469FDB3699B3C4165049C494406B8912EF76C3BDEB245",
            INIT_RAM_02 => X"393521927FC1F0A9FC6ADE49BC6B26E7133A40CEB09361DF393DC78CD0BC98C9",
            INIT_RAM_03 => X"5181070E460490E2760387642783846930E11A4C46D18653C3C140D82423F462",
            INIT_RAM_04 => X"5B54B07F29B44950741442C1E7F0707291849EE070701A658764074156118E7D",
            INIT_RAM_05 => X"107CF045B91046EC3C398CC5D4443640741E618B7645A435181BE7062544C392",
            INIT_RAM_06 => X"99169090BA447DFCEEC9898AA98BAAABB998746465461C666B4E60E49592F0E7",
            INIT_RAM_07 => X"49889B8650190601913B2649C08749D921400292C6571D97559894554020D6A4",
            INIT_RAM_08 => X"C078C96308E316800F3490D2CD1C37D9E6AC084D48002053988B4188D0002229",
            INIT_RAM_09 => X"7654085C9226E4064EC918C17486764554D3546577502CC51CD148AE08CCA438",
            INIT_RAM_0A => X"0AC28339108515C2136A41D90A432404943243407240351321615C6507041320",
            INIT_RAM_0B => X"6053A8074C1C84714D850921D741340509210A8C044101450D4C891C1023721C",
            INIT_RAM_0C => X"0A6121436143437C41A244564DD34140CD2D20341430354334B50B49DE562102",
            INIT_RAM_0D => X"DDD89F35054408005D2D2C03371147614421C323404B1C4D08374677406440A8",
            INIT_RAM_0E => X"99D9614B045241D2418F142B64E14114F209120902C4B4CCCDCE0041ED2D0350",
            INIT_RAM_0F => X"0414B350438D0CC3A2649916433098C90850A324014526031832144E106CC9CD",
            INIT_RAM_10 => X"824C3010850DC953322B001331403616140AC90134214405D00B04C4DC225430",
            INIT_RAM_11 => X"6418D24914303182C5B89D434465762C2D033A431645451CE0010514924DF34C",
            INIT_RAM_12 => X"41657771888205C33C0191414E340304C5116CD451184C900424B7840388A3A2",
            INIT_RAM_13 => X"80911A89121012680C83015451070C8010860526C98531431A07458956446AA8",
            INIT_RAM_14 => X"144511442C4105A0350441081071450212344CC1186360C027C5C2328C812484",
            INIT_RAM_15 => X"130085D0D0C037C94CF14353A11CF3431484623707090DC413480538B0538D28",
            INIT_RAM_16 => X"DE0C985E104C24DC2143430114D5345073709314F24202A0C8F28322245A045F",
            INIT_RAM_17 => X"D234C63362103489F13747478D2CD9324E2C37873AC1E0CE306518673AC1E0C0",
            INIT_RAM_18 => X"1041C91076727434684444332B4D335013A1501004CA0E0DC98530394418643C",
            INIT_RAM_19 => X"073801CDCD033183440C843049364091A218124413243437274C1C1189304638",
            INIT_RAM_1A => X"1296E355966515771521130321655B84064128CA4E214CC00124C7A31B11BB46",
            INIT_RAM_1B => X"C2014C04269D931737019C31515565CDC50451B3C5202AE8A3290CC401840C41",
            INIT_RAM_1C => X"D991413491498C53070C20524D0453034A900A70516C05094007172BA2A9B22C",
            INIT_RAM_1D => X"041158A3CC1C3174D1355CC0C1E0C1072725243625B633881CDC31C330C51E05",
            INIT_RAM_1E => X"8C1130130D20484120320048423004000C046161904C17474054446010CE3324",
            INIT_RAM_1F => X"301D5DD17300C5009F579093820E081161C918A030C8B84103C808C20170B830",
            INIT_RAM_20 => X"403626868EC91032B20C9D60505242A1072968651123016676710D37744D1D57",
            INIT_RAM_21 => X"35634034A94014C1128C86559101C505D818730CB1C43298B0C704521080100A",
            INIT_RAM_22 => X"34D341D935403441C1044D32614343500370C4C4C1853352405351404DD04D24",
            INIT_RAM_23 => X"556445466091460524005244C8311505525460C105C0004110356D034409374D",
            INIT_RAM_24 => X"5AA3649355A000428CD0D43078CA2B074B4D236614D044091E1E1D914B320441",
            INIT_RAM_25 => X"8D5060951DD207449D8D51929B0444A185020C185450E896C36341250001ED03",
            INIT_RAM_26 => X"14C6C1486329808A80945741D83415346D04AA2645698E65821B08164124CD88",
            INIT_RAM_27 => X"9093745324811B14C00934D04B26C50C11A38D0CE180AC1C000B258A445D18A3",
            INIT_RAM_28 => X"01090A0341C050909090909034930C134918341D92649370080D0524B6634914",
            INIT_RAM_29 => X"40D34E280E401082756454C648A80384324068425D1049C10D0D332434BA85CA",
            INIT_RAM_2A => X"A68C5C861DD61C513403A697771C49E9252DA58C01E1E034588D20A143714120",
            INIT_RAM_2B => X"A264D5DE9E91E0C0818C881929324091271C8104EE89958240B0559046424A43",
            INIT_RAM_2C => X"0D0408A0360A106810CE413404D1CB01158915A9113C612DD119D9521549D03B",
            INIT_RAM_2D => X"20240114B4037643400CA0A37433303009290902CC94170A8550016420CA0D2D",
            INIT_RAM_2E => X"38200154120140B1151760482B34E248511778D1342203A26402841108210074",
            INIT_RAM_2F => X"15527893C60CA86100C10404184EE192AA1B28CCE04602418320E0900E018ACE",
            INIT_RAM_30 => X"014815A8B0C8014217667660331405910AD30426F010BCE141010F0114504133",
            INIT_RAM_31 => X"925440441889B8ABA2801CC95176491D3544119D1211331061314001A0076212",
            INIT_RAM_32 => X"E2A3A0A1A08745754747776766764262EA86855DC522B898958999DDD1115551",
            INIT_RAM_33 => X"2544D58320C39000314C438AC83F1EBC010022EA66686010600502132030018C",
            INIT_RAM_34 => X"AA667774445554406733CA264D9064590547646CB320456031040450107C4D31",
            INIT_RAM_35 => X"0000C6338A2408060C04D9274CC510040531455924676664D9064590C922098B",
            INIT_RAM_36 => X"A81F0999DDD1115552222B89A05085121100023302214A1AC5504C8838E38A14",
            INIT_RAM_37 => X"99025499D927491254328C8600E0805924664D9064590C93154477664C2F01AA",
            INIT_RAM_38 => X"8D11244512244204104A22458546D92D193058DA51508730B14248468C092116",
            INIT_RAM_39 => X"5CC9280147648D55186240C01501099A19005215A50764812144D890511D3044",
            INIT_RAM_3A => X"061810A1A30C04D4AA312A84895273394906000C2C0D09858DC3016270C4D0E0",
            INIT_RAM_3B => X"4801C318449356205387040BA5A58C50E9FA72D091240A4A6100526486D99000",
            INIT_RAM_3C => X"DF747115D4520434188D2532269926D8D49158C101A886A220C4D88310576045",
            INIT_RAM_3D => X"4599D9C90E91555690422B449010D48000876C43498637613003674288802799",
            INIT_RAM_3E => X"1438C502AAAAAAAAAAAAAAB001F203F3C2FFF803F300F2413203A00041444D04",
            INIT_RAM_3F => X"24CC11833401092D6872067BFE8A077849D98588D20096038C30C09032700A13"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_0_AD_i
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"57476757B2020FA1C330EFE4A0219769BB80001BABA88B98B9D0B99F48203052",
            INIT_RAM_01 => X"06C56615413D87CD34C541353446D375744E54E14E116735D172CF5E3B8AA8AA",
            INIT_RAM_02 => X"4DE534C783097DC00C44101ED3F373EE147F660376057553CD321C312DF1E01E",
            INIT_RAM_03 => X"DE45171F7914E1F74407C4957747C79D31F1E74C791E4B33D356D66157480314",
            INIT_RAM_04 => X"63DC7177D1799C4317E111C5C4D179931521E0D179919C4DC495317E731E4782",
            INIT_RAM_05 => X"9CF0F4373444797F3D1E12132C49449317EC620F8998005E5120041077510557",
            INIT_RAM_06 => X"BE44B0E0304CEF0133031122230302232110300001334F985F935155D5E7C170",
            INIT_RAM_07 => X"4E80A6622288498919A424690A8661D98458222A40E50390E4389020EAA0842C",
            INIT_RAM_08 => X"C0AC06C029B02984A93A0092412F04711EA0C001445AA21914896A2014853061",
            INIT_RAM_09 => X"667680D0602518902101960B76877B5776CB544747011096284D849C08099403",
            INIT_RAM_0A => X"491EB5D0220F38C030442210086A024C008476534188B0EA77444F3D54898276",
            INIT_RAM_0B => X"A0EA6422A89C0E71AD0A4A90A2A864090E83AA6901CE424A4ECD429424B3903D",
            INIT_RAM_0C => X"A58B044777546574C2734B74A98A22C24CACA3325882316B30743649E93B0343",
            INIT_RAM_0D => X"DED4293A4BC9C0545CACA4B03341579156928032B084288A4427B67A6074AAA2",
            INIT_RAM_0E => X"11E5E3CF1A9A629A6A422AABA4224124900E920EA2C9BACD0E41D741DCAC8302",
            INIT_RAM_0F => X"3A3A9080B1F7002E426698A62AC280080DD48266C8A9A78E3801288823B3114A",
            INIT_RAM_10 => X"41B0B02899D999D5C361176C00AB6667772999C8300460D29A3F1808AED2A70E",
            INIT_RAM_11 => X"66A49A69A6BB5C3C8E889EC24864B714D949266A16566A287E022EA69A6920A7",
            INIT_RAM_12 => X"52855791540B3A801F914293A71F8C088A107C64A23C80292622556641438242",
            INIT_RAM_13 => X"BCB0460B05443194CC9A32168503380A30AF2DB7C29922301415555554554619",
            INIT_RAM_14 => X"20280A00181102607445440AD55357235705244540FF8B0003B515E20C486CA4",
            INIT_RAM_15 => X"270A42ECAAC23A4A419380430320A2053CCDF3293A2602042208E106F391C9E4",
            INIT_RAM_16 => X"21099DDB3397841EE647531004E23BEC806B903A9032825140A23012A49928A6",
            INIT_RAM_17 => X"9106B900703AE442D30683F8483CAF20810F06C207CE7001F083200207CE7000",
            INIT_RAM_18 => X"7202999B96909714A6810D026689005303030304089951D9999921444BA114E8",
            INIT_RAM_19 => X"672FCE418009C05473C088A068B62C8B02A4DFCC2267654666F0E4220DC33A10",
            INIT_RAM_1A => X"228A7E4390E4393D0BAF02092654BA0095A6A9784226480043410F1353353D80",
            INIT_RAM_1B => X"9B0BC40A861E7C351A337B034374A2024288D2C082A9099095D3000D9BCD000E",
            INIT_RAM_1C => X"D5DB6DA69A61A9F0182C0E1861965E28611A0D7BEF70828288093626426B7124",
            INIT_RAM_1D => X"3BAEBCE37061C183E5B94C880A4D480A67082A2B38B80E0CACEEC00CC00D22C1",
            INIT_RAM_1E => X"2D12213340E92903347F84D41B744884CD04935555481495A09496EE91780C20",
            INIT_RAM_1F => X"2C9955953243CFC45E97AAC37AA72A596BCF3CE0300AA355FF44480041457CFC",
            INIT_RAM_20 => X"CFF806A00CC0CCB152AC5E14281ADD63744454DD20EE02A67B4300E565699953",
            INIT_RAM_21 => X"314350747744030A19408A55D201060DE4640200A00403743B00085D2004200B",
            INIT_RAM_22 => X"B2CB22C5B1407699226606A64447475110BB08C886553092A86A90B206DACC96",
            INIT_RAM_23 => X"350D60E0EA5960259682DB77B8E01A08717CF00154C000998075A9256012B72C",
            INIT_RAM_24 => X"4683168315041810B4C49113417CC1072B6C931516C081411D1DDEDB6D243888",
            INIT_RAM_25 => X"CC596A1129C837061C0D1A50662241121160209A9C9C9111332B22A2A8D28CAA",
            INIT_RAM_26 => X"340D0A6A6A0452AA8034A729C1169996610A6816054189151A58C88465C74CA4",
            INIT_RAM_27 => X"C2DB40FF74012F19FA29A65A6F0B4F0812E040178D02982C2DC0474056119450",
            INIT_RAM_28 => X"50455403ABC0F0CACACACAC8269BB0236DB89699CA729A6498A4A63297036DBC",
            INIT_RAM_29 => X"051BAD16A5D855404444457840560754A09046011D86020945CCB04476540111",
            INIT_RAM_2A => X"457014199129907135044774591445110A1D11DD051950B4944D029554605006",
            INIT_RAM_2B => X"4046151DD111D0D44181C450A0A0200900148949110116802082990A64282800",
            INIT_RAM_2C => X"AC0ED86075C60458517444B006DBCC2595BCA66C994C99519219DC5A654DD004",
            INIT_RAM_2D => X"6E80270A900149617241194046A07142A0A0A00981155F05055A8902A211ACAC",
            INIT_RAM_2E => X"D020A9461AA96AD314179002AA1073C4A21797E0906DC84046A981172AA04810",
            INIT_RAM_2F => X"08715FF14E0991140B0212901609151A4446667040B50523800B0E00840B4100",
            INIT_RAM_30 => X"106CA6146F0B328AC775796C9F088994094008096040980D65A40525945555E1",
            INIT_RAM_31 => X"514490A85455454460682401108442510954615EA020136011928410140B9744",
            INIT_RAM_32 => X"C04051617047857957947847857941551101C12E418045544A71911915D55D51",
            INIT_RAM_33 => X"184AE12C03890000451142A1246829F0002CA5111110141A9228644445445517",
            INIT_RAM_34 => X"5565565676676688A8C2FB0681A1685A066554A4AC2C86F29208082823AC8A92",
            INIT_RAM_35 => X"C0044193400A0BCBE7A4E5176B0124EC41B24190A4B7574290B42D0411128665",
            INIT_RAM_36 => X"AC2BE919919D5DD5D8312677722409A2975176064064B2064118B84B2383422B",
            INIT_RAM_37 => X"5D040601E580605815047899404F01108494210942504119D6564545574BE1AA",
            INIT_RAM_38 => X"014A04900415129015458D44554AE18121E020E9606B0B1060418A4538062194",
            INIT_RAM_39 => X"EC8B60095446355128954780212601112589A1282B27A852A073E058541EA152",
            INIT_RAM_3A => X"2EFC2A83436DC058D81236C80DDB4377BD8B0700144A8A8ECA4001B3A004A454",
            INIT_RAM_3B => X"8002DC04A153B81482FF388046678022BF6FFFB3D2A02B6ABC05A2B6B1D5DF2F",
            INIT_RAM_3C => X"1D857A55EA50013A248EB8402DD28AE4A8AB438A336CCD83038C20CE32B5A8CE",
            INIT_RAM_3D => X"88282A8AAC8260BAD8A336A0E828E14C448BA513AE4D3BA856ABAB9280C48761",
            INIT_RAM_3E => X"2420C2F2AAAAAAAAAAAAAABC0BF300F202FFF80FF802F1033183A00002088E81",
            INIT_RAM_3F => X"170021A3380020177A8EDE4F635791AA05E5418AF280EA2AC58380EF33640CAC"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_1_AD_i
        );

    prom_inst_2: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"7646466748BAA6697570547038BA01111367A9A60231012312043231030400AB",
            INIT_RAM_01 => X"50101044440104114115114045101441001015095010504005857C825F5DB5DB",
            INIT_RAM_02 => X"50004404141400155111541007F401AA45400614060504040045404141010590",
            INIT_RAM_03 => X"0025549000950904116420100424200049080012004024081020240640901019",
            INIT_RAM_04 => X"5402094404451058000108250509411854511509411941012010800000802014",
            INIT_RAM_05 => X"4102060440420000818054104215410800011920110452200544458040116200",
            INIT_RAM_06 => X"0901020845200002100221032113321033213321032100411010488011040980",
            INIT_RAM_07 => X"FE2D1115F4571434A6D0D2B6B6A9A866F302966430484100C0312900EAB80100",
            INIT_RAM_08 => X"D8862E48CE18A8ED80B8B208642CA0B82E009A3C11CABE9B9AD1C489C19CA6B8",
            INIT_RAM_09 => X"0929308E1B4AAD26D81A623A9BAA3AA22971A2A2A1C846038A20E1CEF8ECC282",
            INIT_RAM_0A => X"2E08031B5A04C222962242A92A936C27B2622A80386D14F0A23B8C3198E40529",
            INIT_RAM_0B => X"F470BB6347070C15B0103EFCF34B8343C7C383002C5C1C961CB2780F8DBF0430",
            INIT_RAM_0C => X"A461B3322AB33BBA920A0AA09A9262D977270C54610D5581DE10AAACEC3743D1",
            INIT_RAM_0D => X"0C2180B8A920B36147270628DC0913851A84A3860CE18A9831B3AB3A9930847A",
            INIT_RAM_0E => X"8ACA0823A8E382E394238A988108A42D0BC73F470CE0BB327C508CD8472795DC",
            INIT_RAM_0F => X"0C0E1E14BC828E0B8739CF33C005F21F2CC383B8A08208E6823860E69B808822",
            INIT_RAM_10 => X"2841B622CCEECCE307994C2048AB33BB30EEEED4FA8003A2AC83A8ED001F0830",
            INIT_RAM_11 => X"3942CB2CB28031A230420EDB0AB09946AA387BB4DB9BB08A20A38238E38E3884",
            INIT_RAM_12 => X"9D2182BD10AAE0A38886140C058820CEF0868EA30386BD82C2FC0088080AEB87",
            INIT_RAM_13 => X"921BB9A1B220B41A142948681A27965946A18208EE0048C3985099911A91A8A1",
            INIT_RAM_14 => X"85C1705C96442A7B2199EB222A8E28462872C15CB2729010AF4AAA59A5039A23",
            INIT_RAM_15 => X"83EC52CF2DFBB0221608958B812538A4967219F3E0D8783F38A229903A8D6302",
            INIT_RAM_16 => X"86ACCEE1888C6360330B878DDAE8BA6A8D882B400AFC8A692D388384A1206585",
            INIT_RAM_17 => X"0858C0A594230E32F8D8E329A28EE386242C982990EA5A560880222990EA58E5",
            INIT_RAM_18 => X"4812EE06838E00C0B216D23B30E085BC4B80A85A4ECC2200EE0048010A62220E",
            INIT_RAM_19 => X"53842E163322058884528E380F33CBF0960210EB3B308803B80383382278419A",
            INIT_RAM_1A => X"39982307C1F07C0DC3F5896688A03DA2A08244C2308012321051604807004021",
            INIT_RAM_1B => X"28A02B06A88E704B4BE48C38240020705ECE0208E2022CC1E31BE332E4628ED8",
            INIT_RAM_1C => X"888A28A28A242008E2EE28A28A28A5862A8A0E80208E0303530541B307A015E5",
            INIT_RAM_1D => X"AAAA863881C70614CAB29ED65861204BB861E1E1E24031A2A1C205670CE020AA",
            INIT_RAM_1E => X"90A415A4650ACAC84A61AA42C102505651B0AC88A212AAA884A8AB3298C23074",
            INIT_RAM_1F => X"9E00A00A780AE0064ED3BA3840A580A2A823863A48E818AA73E1416A0A223642",
            INIT_RAM_20 => X"E738DA223EB9B14E842E8EA123AE886AAA221A0026258AA2B29C650082A020A7",
            INIT_RAM_21 => X"54AE07922A90941A4C0E800002565850E18F5B4E8561380080358E0038AD3968",
            INIT_RAM_22 => X"14514252148B2066391012513BA13ABD050010B0142299860AAD84169264F508",
            INIT_RAM_23 => X"1A0680C0FA082782084820094D59A8528E8218EAA9E006440698828001A25945",
            INIT_RAM_24 => X"B005480548B08259895225B498C29969C9971D484072FE1C84EA0E082381E0E0",
            INIT_RAM_25 => X"158A28CC20724968E526EDB713543EE2CC09C16247650ACC494142A261222500",
            INIT_RAM_26 => X"CA947A9A847B2E980891A1C8788A0641858A0048122C10CAA6A1237383101501",
            INIT_RAM_27 => X"38209A00016403A9038E382083B8E0924239A68C69A6EB2FB41A200BBAEEDA68",
            INIT_RAM_28 => X"7912A9CBA9620A1212121218B2C803382082082C330CE3962D0301CC80C82082",
            INIT_RAM_29 => X"3EEF0092A4032208686868C61A64BA9E440FB21ECA6138D0303B3A232002A888",
            INIT_RAM_2A => X"2101C1E664244F78E07A22A90BD234882684EE002CCEE5809AF26AB333070570",
            INIT_RAM_2B => X"862964600AA84561587E51CB2B2ECDB3EFD2F416AA18A20AC71646B11AC2CACA",
            INIT_RAM_2C => X"0B23126BA926999E78C61B6CB288208A298119A1618E44EE42A4634826F028AA",
            INIT_RAM_2D => X"42A4A7881A89090505288B8739078716AB2B0B21688AA0AE1CE6D76C0E88AB2B",
            INIT_RAM_2E => X"128211924AA92A3AEB633DC900DA58E383A390C75A41268629A9A6678067155A",
            INIT_RAM_2F => X"D29E9439E0ACCEE929E3A52CA21CA8A72B33B9C148CADA78239062B234A809A6",
            INIT_RAM_30 => X"6EB3AA939C14B5662A223292619AF2072078CE206A521A6124A727861A44AA59",
            INIT_RAM_31 => X"6A20A60B23A2A2A28694923830E0C3830E0C3C6CE8EA969E1E8F3086908B22A1",
            INIT_RAM_32 => X"2A86868687B33A32A32A32A32A32AEAAAA3A182C3AF6AAAB09C8AA8AA8AA8AAC",
            INIT_RAM_33 => X"9A08EA404DADF000F33CCBB17C85317000992333333117E8AEC8684C4C4F0E8C",
            INIT_RAM_34 => X"AA2AA2AA2AA2A958040505A96A5A96A5BA22209E40526A7A69AA26259B926669",
            INIT_RAM_35 => X"2022BA7A0BC979271CA3CAA29C1825971A5EAA8B202A222C8B22C8B288947AAA",
            INIT_RAM_36 => X"012418AA8AA8AA8AAA4EEAAA0E2DF986228628629628BBE9E8AC96F4946A09B9",
            INIT_RAM_37 => X"8AB2689ACA2689A268A216223269AC8B2022C8B22C8B288522A2A2A28C642C00",
            INIT_RAM_38 => X"58B1602E68E2CE2CA2285232220ACA28286A23EA8E9CD6B73EACD26C96B349B2",
            INIT_RAM_39 => X"81D148AA222140A8A822B16B8AA1E8882AA8587284A3A1AACE9CC1ABABCE062C",
            INIT_RAM_3A => X"841EEE69858723AD468F59E1746D859906C8694EA13838383853B42E14E18381",
            INIT_RAM_3B => X"3322406B8C83686A884592DA23B962E2A7A9DF5C4EFC919071EA84198A88A7A4",
            INIT_RAM_3C => X"85EA17A85DA22C34E30D2B94C442CAE303258964959E94684D66E5759B939A6E",
            INIT_RAM_3D => X"48101EF2BA01206A6C86DA838FC0FE9C388B02C34A1437A380028B047353A17A",
            INIT_RAM_3E => X"6BDA664AAAAAAAAAAAAAAABC0BF40BF0007FF007F80DF803F141300222048D30",
            INIT_RAM_3F => X"91A16E69B8005F0BF16E472ADF777CBB28CA3A1269A22685E245622486962270"
        )
        port map (
            DO => prom_inst_2_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_2_AD_i
        );

    prom_inst_3: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"CCCFEEDDCCEDDFFEDED0DFCDDFECEDEDEDCEDDDCDCCFECCDEECEEEFCDC5555DD",
            INIT_RAM_01 => X"5D5D75575757577575D55D57555DD7575D5D755955D5D5D75C7DE7DF75C71D75",
            INIT_RAM_02 => X"5D7575D75D75D75D75D75D75D6ADD7AAD5D7565776575D755D5D75D757575595",
            INIT_RAM_03 => X"75455515D515515D55454555D545455D5151575455D54551536565565595D759",
            INIT_RAM_04 => X"7554515D555D5551555D514575515551557557515551575545551555D5154555",
            INIT_RAM_05 => X"D5545455575455D5151557555455D551555D5145555D544557555515D5554455",
            INIT_RAM_06 => X"01550050554014ECCCCFFFFEEEEDDDDDCCCCFFFFFEEED5D55D5551155D555115",
            INIT_RAM_07 => X"211FDDD9BE662726361C98C63B9DA27608B07E1230D8C360982363B0BFE85540",
            INIT_RAM_08 => X"E2B0E6F0F2C39B4C7D1122D3C22F0B22CA20492332367367B0CD9892332348E2",
            INIT_RAM_09 => X"8588B0B0D3F33FC883210F28D89CB488847989888989B02D34F7422EF8466D01",
            INIT_RAM_0A => X"2607DC4B9F08CF027888B122286FCB23220888B9C34C98E888888E388B86C989",
            INIT_RAM_0B => X"B3ACDBF3BF3F08ADC237330CE3BD80EFFB02FDA22623233A331073233FCFC022",
            INIT_RAM_0C => X"922C0888888888BC32E08488422CA2F4E6A68C9E238C9CBCD9988896E73A02BE",
            INIT_RAM_0D => X"2D233D118BC6233336E6FCC1D8888B8C096F412ECC4C34FB325B49B4848899B9",
            INIT_RAM_0E => X"6446E38F29249165630F096863E382AFD23AF33ACFE69CC0FFC075B666E68D8F",
            INIT_RAM_0F => X"C9CA08CACF9F0405C99626C9BD4C62762223CD9B06965B0C3810EC4E3AB522EA",
            INIT_RAM_10 => X"D35338212222662C4C88F5D4BA94888888F26630BC59A223239F284F7C7CF915",
            INIT_RAM_11 => X"94B065924971C4823BB86EF58D98D8B0222C99488C8C8C34E7811A492596F0B9",
            INIT_RAM_12 => X"B8C888F88897CF413D4DEECEDE3DE484BC0DBCA3B138FF3FCFD88888888825C9",
            INIT_RAM_13 => X"B0C19FCC19988CF87F67D59B662E3004F81E124BCA66E3510C88480084884000",
            INIT_RAM_14 => X"59B66D98BC6626D1999B462D5988D8C8D88DA32362D4F5220BD666E3CF3DBCB3",
            INIT_RAM_15 => X"0BC031DE32F0774200D08C8B822FC30E3CC0E1CCCDCB7B73130E4C08F08F8E78",
            INIT_RAM_16 => X"3E16622C38B1232C48988F80C9CC08208CB1F3CFD0AFCAE38FC3910FE238873E",
            INIT_RAM_17 => X"D0CBDC3C8C2F7830E0CBC38B8C3C2E0CD22F0BCC0BC2E132C182222C0BC2E043",
            INIT_RAM_18 => X"E3216620888CC8C89B1000119BCD0C90CB82C040C46666666666E19888A66D70",
            INIT_RAM_19 => X"5471EE32362C4099B5FB84F1B6C9B76C8EF0C7C3119999999B533313C2F39F3C",
            INIT_RAM_1A => X"1286E58260882208C32D0BCD19982B8248512B123E19B8323055455154055545",
            INIT_RAM_1B => X"670786ED842DC4C5858DB91199D443232B0462E3C26427736C4B9200038C04F3",
            INIT_RAM_1C => X"65659659659256E0DCDE056596596C189326E9B1E5B07A7AE6EFD89DCD885DE0",
            INIT_RAM_1D => X"8820B8F392BF4EF9D6B5B8323BF78C8598CFEDEFCEC6178EA3FC4B0F48422056",
            INIT_RAM_1E => X"AE0DCDCB0E69B98801D7426269B83F372C188C9999B85F9E8BD8D8F54B1214DC",
            INIT_RAM_1F => X"3C216216E088EE446B9AE9F3D69E1965A78F38F0AC493966C78373758999BCD6",
            INIT_RAM_20 => X"CC78C0B22EF762018FFE6E62237266E19999B8722D6D0999118B8E4405A1016E",
            INIT_RAM_21 => X"DD8CCCD98888BD330184A2642AF23332E33EC3848B021088B12C0462109F138B",
            INIT_RAM_22 => X"DB6DB266D9888B66E19B2119889988BDCDF137FF3766788CD5B1C9FFE16277D8",
            INIT_RAM_23 => X"26099090A9659E165989240B97D3A8AD81B8E0459B802966C9944259B26119B6",
            INIT_RAM_24 => X"9BC19BC19898B0E3DF722E3C8B120B95B946CDD8DF623333662224249F0BCC4C",
            INIT_RAM_25 => X"2765A766226DC99F262721FDDFDA367222C1F25A665F3266D1ADB161110226FC",
            INIT_RAM_26 => X"C9F7A86860912A28889889A2625A65996D08BC1B0626F3652A5B4311BC7527B3",
            INIT_RAM_27 => X"F165BCE59B828F2B5F1659659F2BCE382AF38F3120AF2F2F0D699888CA3230E0",
            INIT_RAM_28 => X"F19998CB97C2E16D6D6D6D6499671311967859666D9965BC6C96DADB99899678",
            INIT_RAM_29 => X"2213514BF229998898989B12332E19B48CCD9B26659833F33336F99998889666",
            INIT_RAM_2A => X"8B13333666266FE0CCCC88898BFC33222266226622222F4AB08225888888CC8E",
            INIT_RAM_2B => X"C88466666226627327233232E2CCB02C0BFCB73723221108BCB0652D94B0B888",
            INIT_RAM_2C => X"D62E7CE19B8E19B4D312251899678E165B16D9E66DB866226166566906F46488",
            INIT_RAM_2D => X"F5589D09B8488C8CCCD224C8844CCCCC62E2D223C2266E132211F88A4E2266E6",
            INIT_RAM_2E => X"78626599665599F29A9F69C86DF4E3C3311BB1D734F788C88467866D19A629F4",
            INIT_RAM_2F => X"ADA1B9F3CE16666227C10A488B26221189999BD3E056F6E38135E6223E188B8E",
            INIT_RAM_30 => X"8DCF9999BD3E0B8D5995B5B8D789F45226F0C426F122BCE492622F12492266E2",
            INIT_RAM_31 => X"5598BCC5999999999D88B4263098C263098C265D18DD913816B3D88D98875998",
            INIT_RAM_32 => X"25CDCDCDCDDB59B59B59B59B59B595555577261DE73111110716566566566566",
            INIT_RAM_33 => X"B9A976D40F0C480A308C208886489D50024FD11111320268FF049888888988B1",
            INIT_RAM_34 => X"449489489489482A1E4F9D1B46D1B46D188888B8E4F8EED1D3BB4EED3AB0EED3",
            INIT_RAM_35 => X"0009F7D18B843B0D7D50D659BD369000250D96629A19958A6298A622227D9444",
            INIT_RAM_36 => X"0F6D6676676676676B339111082032C81D8DD8DD8DD8BADF8670B07E31E18BBB",
            INIT_RAM_37 => X"66589A244689A2689888B066326196629A18A6298A62222F58989898B12E4600",
            INIT_RAM_38 => X"372CDE08DF14BEC88895F5999988D6A626C122E18DB1FD393D96FD98B05BF662",
            INIT_RAM_39 => X"32CD8899999BD266A2599B82B65B86458696E03DAD1BA04B1DB1D2637276CDCB",
            INIT_RAM_3A => X"1C7431F1C11E506F7F0FDFC03671B5175708118453333B333B210DCCD8433363",
            INIT_RAM_3B => X"23B2C4D8B66388108B1F3429988BCE605B16C8B163148140D41188DB56656C1C",
            INIT_RAM_3C => X"6C59B166C46A263B238EC980E6630AD230118B8D3DFCF7F00F4EA03D3A9BB0EA",
            INIT_RAM_3D => X"882821E3C282608A7080D8B33F38E6B333A36663B237392D9BFC474AC0C2DB16",
            INIT_RAM_3E => X"D9F8E2C2AAAAAAAAAAAAAAA00BF005FD08FFF00BFC0FFA0EFA80300922088E30",
            INIT_RAM_3F => X"1B0256C3A80204BF515421BC4914440896D63625F3026F1BC28F426F01BC26F4"
        )
        port map (
            DO => prom_inst_3_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_3_AD_i
        );

end Behavioral; --Gowin_pROM_basic
