--
--Written by GowinSynthesis
--Tool Version "V1.9.10 (64-bit)"
--Thu Aug 15 21:37:18 2024

--Source file index table:
--file0 "\C:/Gowin/Gowin_V1.9.10_x64/IDE/ipcore/PSRAM_HS/data/PSRAM_TOP.v"
--file1 "\C:/Gowin/Gowin_V1.9.10_x64/IDE/ipcore/PSRAM_HS/data/psram_code.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
KbhsnglLlH06TXIaEjajkuO98HWcEpYnCimXSYp5b0UYsE9unK/gGFsQnY2T417BdPAUb+nK2Ok1
EJgwE9HPAW6sGiAHz4WfIpXyAKvlH62j7h7MingdULYidMG3pb/QzXZONWLF7RNoUwim7df/c0fJ
xiHbAtlcXH9F63RKPw2w07gOOedHdGjO5JMq6Rh/QRwq+C2AK7/xZAv3QHP43jtGAOfon1VOhZ4h
tlrhKGl/jK03463btxBJhTiYjrlkELnG6Q1Z75D3h8Wv0/kYlrumkeLCIYOwzhsU9O2UEaCVE56M
nfBLLVE5c45IUrar8c6LD7j3BbXjxgO37b3LJg==

`protect encoding=(enctype="base64", line_length=76, bytes=310448)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
UElGxFoVYTf3nep9xJz7VWtZu7wXcoYuqxwroET17USkkKlYEibCWlz9JLNxfkPM1sTNyNdrLGRg
2yiqjZ/oY3L7lHgFS3NR3TkLnjU/LG0BWXBK9FmL645OQHG6esKaapqKgsHPT8akRbCtFULBAB8s
Eu/+cyfUIyWHt37u3Aa9l+guNAKYhMaTvB4JLZMsLieBXPElTqHgL7peUBGdZ9X1sOFbwlG8PM/z
Hi+xipUxcC1K7eKkK8qOJDGsWdzBhEzG/+L2A6l90Jj+IqZwSJi+3cph+4vIAlzFMGsQLfMvXdFy
G9V+F2yryJ9j8x5MWcGSHp3dK1tWNKX8z7iSNS35Yj2tb+ZTM/xznumtiOCHTXSte3aOmvIeCMJP
1TdaWd69gyVVM3RSJoP1ZbAX1eyBrMYWm/bD5f7I0JYqBRVQIO3r9G8XqDmTNUnc76yoqJXQx6MQ
DKl8VbecFWzuLttg7B5moqdPFIpPZhxwcwBTAzFTek2PmiDlCc/IHSqlQNYV8BWvmzbjyITXQBFZ
caDaha6lXMhTPPntl9K6aWIrkcsHH+Fyo8nRZDaSKYqOFBhmyE7gH4bAasJR/V43+ZmORTU+cjg9
Wm/1Y4KlqxgDOjQDokD6XJm6pkgJN+KOJMnv4UKWvNjskIeDLdRpcMFrZDs8SCB3CsOJ8CA3v6LW
qKVVF/5RLCz3VXALBUNT2LQLFXl5+Ij/QBSnAp+Blwk6vclB4iUIgdZQ5TdxpGXo5q6rXRII8sVI
eBSXnJXj5qMtijtO6CSXmx7PkG903HL6Ug0D3rhUDsMCePHnMr81nSEXN9M2JBHyw3a5aqoM5RlY
RT8Ni5iWYo9NaYykeqXlyz0kr5BmJ4BJ2WgqAZsTFsV0SOhENJ2V6DplA5XIsXd6hKgLGDf+6+jI
oxqnDwn32R2A835A4cjbFXicw7uiVq0yzgilHdvX6cmmoG8OxxHW4zTxVXsP0zyPCWyFOJrOQKHY
KRlEAKYy82xvWYG/7NZWrVGpQr0a6a5RQ3yTU+nTD1OsqgLdbLxDZ/M9NyNr6U5BwTpKwhM5lyro
OF2BL+Ej5ElN3cU4cKPK/IqPWiaG3peHis9uxa6EQ+8OLEtmoqgqTyghcumOnSEz8ii2TrpT89vk
grlF5MWVuePOUgqdHmnjqY1qMfbnuMETiUt/Gpnc6QsRrzh/zG1mSYOqOYmebTeHjxTYo5rRwjmU
gfgRHvegi5X99T/Gx9tG8Pz+q6pAqiBuBXjWPTH8WbRI/sTAaa3QUYncdjV6Kp0vNUrHIABUuYIw
a+OyfQXXHYWZ1iPVCJHvoTBwbHSzWai5XSYYPBXSC573e+DXbyYmZRnr0naIsk6V/hf7gm5gxFoF
Pj2nlz5Lv4UzkiIMJHB/T7hqpozZrgLmfzSYJU2+SmEiILbPm397bH7n/6drXVYSTPL+Pohz9v2a
k3v1/ohFzSeY86wV26ntoxMGfJaa0K7dlj8xd5iFWhgvasAIO1AKYCeDyvZtWqUQz1Qq1aY4C1+A
MxojyUlDuX1TR7qAPVkmQZ/7l1E2QmrnJXdOa8f05qXh6Dh+FOSi9QMP/Q2YiosC61J15mfFUTff
w/UHXL4w7tgFqJ0Pyudi3YLxeZfelZ96Bu/lhe+k+NvLieFo9xvDewHUZuu/eczbSWJ5KvHc9Cug
RMgzbQdDIvI1Q6Jf0y3pDpaD5+zEEBLS6Q1FRh5o/3FrknVGUJ/7qrID3PgFQ+xCGG8t65KY0Vd1
uAHf9lsbdOUUAE2yXObGXM4ux420Oh1qgcdwIBQoLzRQHqDrdrjEc+xwuV6b0hkoUgYCOVxqR4Bg
by0QXZ6Y+2rvl00OjfNCJxTQ6WRVe2LO8Lx4W4tBLouO+y1pVUp0rCvSPmC+EUmn37WWdD3ljsuJ
aK86Oex31BnsNxR3BcD0d/chVHLIqyMNRcGWmtVQT1w0KsmF+8UZPBnvZsbWXFWFrpv5/qe64nm0
KpaBOZHXRkPhOrsSll6CSLLxeHbK5Kk0fbiUSi8d4TlqOLwySvknCpoAfYlUQErIz+x7lP7/96LA
z8AMIRe25WRJFjwfSgmd2eE11vbLBYmnvO3OG19IV2T9xaB9mHY6PJ+YiR1q0Z7MSRh/UJ9T+aFC
MaIn53VThqXT7GJjV8qm0pI7iACaF9ixJZXk3U46nsRVRI39cMXb5M5NNU5c0VJ/TNH9g+e+n0Lm
9ZQvQH4WuISGDgCEVbAwwlBULhMIPv0QGqOD58oOtxAZRWuY2H9ur2PqeNorMbpQPEAM3bt13+bh
YXo3k+vqXpIiw/bDz/9fgFL1GC8mcf6bbtL4ultxmuGPMBfjjHKUYlJWmkWQs+g7z7Jz/YVo61Tq
jPYWOJ98fN4XsQ5RZ/aAhfzbYl6hQBk2DjBe9XKeofzcHes6BwaURgG5GVGmrWf+Rjb9dKK0WVwB
mDOX/z0Yw4E4GJzoxsgNjXe+w+GiWGdq0zPda9DxITqo2VM3Ik6+CbFjlk4o2EI/epDqwTYPfgkq
ZV6EzFBBPsYVKDwJXwA7/2pJ4x5IgxOKgn6Nn7JyR8OZLb7f4ZhIyv5sFHDe0bHZUGf6D9ltfhWq
W26bD+hHTLy/IAz3UkZ0RIbbJxAlNwg7u4PhC4StEX7L99a70GBOsPDFI6T2ho927IttO3WM3pR7
+cSd8bjpzR8PSXyCy0nbuqyKSiqnDqiua4nKqpwOnS+7GfGpNKtaVrkMP2n+KVtpoS8PANjU8oxN
MlH/uNw4DRhBw2fb7adWyEa3D2ZI/43Wucr6Lq0ADpwhUuRwQU+KAZu2VLBDghyDZbRgD7Qa2JOG
m5YkTABdyOhb0RLdx1m2FryRmL8o+elR1hsVlQ83Vs2/TZ7u5qyfDm75sQnaThkexUqx3WyMBMhF
fmZ0sH76LfU3MQexsIjA8ZrL5P4JwLhgXYPyO9cgQItkc2tl9nDedwJC1yaxzMZbF6nzfh44cY//
aI6CmJYV1LbSoeCU78J10uLNhYqkDATrVGpMOCy6NueRbcFHCQ0JxhrMAJkCu9RxgGHS6FOpuiJx
ay80QY+q+RC7Z5i+XX7tfM7Fz4AX8Q4sSif85V5Fi0DJe8kUrYbHkZ4oD0+oTsppiJcWDwW83pml
XL/CTta5ju/z32wkujj3gTTUa1ThDrl8jUcDv19g1ysblRstRA2O0Ns/aa96leb1SSnd19F9D2Ok
Igfe28qdKsvIbzrgLoudp25RwjjnJNJEsanbT3H6h2t9KuXDrOIDJDm4jG80RdrY0MwGvNfVEjcw
O5K9FlipmsC7aE1h1TR0Az24AmxL1muZx74cMrmUqFbFvFIl+5lDpmEfAEKXlHgi0r1oSLrEQRwP
MGghLo2KwwC2dRa6gcRZufGJMiHZBkif+K3ZZFhApxtpPBZjQ59DKjBEeoQu0T/owVcxjgYRi27o
DTEjsHLkNpHoHDYvDs/C0iqtNeSf7WDl4nYSDiRXv4MUmvqp3ypLMpcUs8/9zl8rm9nThfHUugrV
KQh/aMlJ2zhoVAyTzv6msVONOZgMdr6Y1Gp7rMtPKIueEFj9C+LfkqQrEcS2ddBJYn61bOWazlUP
gjVlElwgAF19eraG70i09EBbXsBeB3MqD1ZR2t319vUQ/a9A/PKLx/yJCk+1+/Ko+IDCj1xkXIYx
ryV6Y/E86KKvhkWJd2rW8MZVU/70c2xajTBSCSxAryoYkthQdWgpzPXbKEves8tpbQu5Ya/T+TvG
x4vsoOaPz4YVQa1sTzLIsXX17kBC2kM2D+yd2+a9+h2l9J5pk76rOWBpCoaWqbqDAscZHtwrlRNe
CtoMt/K3UyOBAdRMbYe7pd4H/fH23z8QBTsX1T34pfgSplW97JHcDcEQynR0s6ar99mr0EniyOTS
g9Ykxp6EApe3TA3yVJhZ/B3L6TT4qfYxPMdwWw53CcnG+m1KJTOO94APjihGiH/QmyNbFf6JDmNg
4MbKApYYIa+cEJYRBdHp6GQP61Kb6rkcFl6tKAEJrJ8O1znBEXH2t1fts0vy96rTqWk2Zp2cMR9y
6y7xezGXnxtLnKhmWtQRAmS0cMilAEyW9Scia0o3REzuwa88Yy0yxbBZOfFBSCGpcsP2md/6WpcI
oZ4Q8xD/bZnsVzY8R2bCa0cd1f/jRFIT3Vw8//llpX40v9yFBe+7oCVP2pnvblJmf7/qM/BN1cQ/
qFlXPfysdHSnsNA8BdZgPVJHtwAlvv4Hb2Plw2yAVk8OYUfiYz28LqAdd/HLX5DFZJBiDVqeH0v5
Evi3KJsZ3fji+Nw4SoD3jyYg73on4brECjYFkWg1AO3pJ+BMPPQmjDrMyFokcB2CmtsmodQrM9R3
QINApiPhCf00XgPRnCuYQvd0Pp/0q32FoIBfV3E0iD2FW/vlEeGGsa9tdnPDqsR9wc+qJuwKHFTY
x78fp0+bR4VYRbFfhfXuviBdgBrEV1MKe6cmgQaTG5wbkUJLWXJXMu/6zyzdO+J354W/bJ0G9GDq
Nm3QP9ZnJLV9G1MZ1vME35fqBT1h6s9nUklwlahznRrI6MVxrGjQP2OeAhDfhonaoa1tC/vm9opX
ogot8apVJEMbA3zz2Rb54LWp0mMydESAz910IAxF2qqhT4ozLw3ZSSd8uRPnQI+wGruDDm5Vetlf
36PgxV1XgC4NfeaHnbn857Oxx8pnot6blRexkS0b4eGNHIdd8XXs4UP7mCMR24yYzQI8pvifEN72
789irSrIGzHqcTXufrqwHMAn8/l5+JO+jIsHW/9Wlc018BXrWn9Xz1mOBp4pxGbAvlQbB2TcRCIJ
7WSOSU1QyGWeVdMPOZfFoocC1H9bmcvOhtXgxNHVcM7h6YxBzVykrf9LJbHhQ0Vbp5UOA6BNz7u/
Z9Ht6A9ql5OCcnKUCoL6VuNrf9NWErS2c61yDDPQsTFYXVQDlJS3HCs6hsB1eruvuf1IxJbyhIC5
7njscZMvtScwCUIDcHbyfTUBPOMcw5j107q+deVKpO9mK2FtkqxCZNOCm6jxTaZV5Cq7Iq8XC6dp
2a9U8FohCqn/e7DbqacU01vAQSLz1aKCs7yUuiYgQhnJ+vSMp4Pi8mJpaN2HdPsxdo+qN2z9jMxm
uvcv0nY4PQ/F0Ui3eILj0Yrpp0SslUFC11oftofdldb/h7RsuMsK5TyeAvHQgaTcRT/qjzScwOKC
k+rbvNq/HcWDLiKz7MpQmIWT5nrueJcDc17VqITPGIpw5JNT9ZCQP2b1A/6IrsNaNIpMisCU1l1C
n9O6wisTuNTCSdpuKxcg4wdI2pKdT2REfsezVjjLxeCZVSQvuQfo1flSGO50FjxOTY5m/56bNZEV
sH/fN8Weqr03mXR2kUXb2uqsasKcF79y4uEbjHyWGW/msw/DtzX620vOYdfEHeI6pGYW1trpBK+Z
mWsl63wzYWdl83Xw/m2ooPytMjFEGjRKFGQ6Z/5YGUMKwWWkb2XEReUiJszB6ygUgZQdpBXkHG+l
Dk1FZQd0SKp0eoMb54TUU8U+TxdGZczqvuVALhB6GWTTdn0QYTYAMf+kpq/4wbN0N8N+cmDK+R2l
tFbvsIQ88bMta7eHsJ3LtPkQQ0q+hZ+A4iEcDhHd2Rs0LeC5KZTk3+AAeGmb+yjKRaNDuJo2CbTc
IKDu1/HQnBZ/6ldqyuGOfuwpzIU/sFiFZL9uSwQJGZ0bicOhAsiKMBnWXulTS4CzOyFsG6fAZfPk
+O5plDfX1NJ/Tq4HxriGYRuWDB9DYpwNaP1gnLwKSgVC/W9eb6T2pOhhERrXU1vNkFnmJQmvGX6Y
SxtFM/2w4Pj0xKpRZI8S5Vl4JkdAm3ODZLibKKarvwea3o37u2cnOYP/PVbeNdpXzy+4MaFDUPvX
DsbYpGaxv55oao1RcpNz8xh8WYSvA+gpZeMt30NTE0OlfJNe4rLaJutkeW6dF54GwHqyLwbxdHjf
TXS/5w28IiK/EYVtaRvjU5jUT+zrf6wMnB/B7UoZeniJIyuE3iud1egylcqXFi+hT9UN8NFMIpeJ
/mitamjmI9l7nc5B0x2c1LIyLHRCL6FlghJWB1kzZiOyRMMnurHaUQFo3qke5+8lmfyoJrD7midg
pCqrzOjaWTz8iJfPMUTPkvhMecam1UE5Q/JsYCDICDXVpEG16LS96TnMR0jYa6G0B8e/ohvwaEAm
Cu6KyqkCKyDW8ZXrhrjJYrQDTLYHVWWQx/pKZIsQYQY6V5hXYjFY3VKKak29rjZ5L9yeI0WEABqL
YoSb55mm1kXUJPxG5Q+bGaGl7cgiwzTWkCZY1/Na6uxU7DuwZBAYrv95x7TxdjvTEHBLJhq+9B8w
6f/Z4plrOhBRqNIFRzsAPqxtWLF3Clkj0ITqX9QJQG7a6ljVLyATzOdSYXb2NHjaIGVBse4NDuiu
L4QHYfOxvfLA3Q4QqH8+XGnaE9wZA/AdTij7xJOTz/LzSJ/4MPvNHpD9qQwAeIilzH4OcAUdjJeD
qlnnctZlMpuvg90lCtVEL5EzuC2B3lOepE+Haq7YrmUS7fSg3uLQ2v+FZ88iiQUi0pKBRSVfgZ5d
QkrIOdtNdGZyyIHVr9Pl5TVR1IJWt4DKPHaSjiu/6MPluGUMU+E4i2AHzb/OCko1orOBIM4BNgGT
bYQgZiTC7l9mnU1KWn42M4npMqOqkXroVP8xT0bZTOKd0kHlHyaozpI3TTZ1H2opp5cqGP93mSYS
fcQn3XWLPCZOohckGsjOp2aMNNMkmbp4uXlFDb2g1Jv/il2I/AiqrXWgwEgqFQhSufXA0pZYyivI
NZTs0jZ96M+N1v6Dwnq7aLSFIJ2Hw7t0UF/Rxi4gxVIyWd57JoxquOygUWZs5Fub8+Dk7jNT3QeG
Yd4Ylqh6FkwkbJQiT1BSmSqYSC/eMB0gtvifTGvS6YE5ihMQZOxe/j37kS1V1NcZlQMgYGUe0wKr
PoR/Dd1Y/ibaqHq96hT5dmEEzndLlE2wCxAmw9PXdE3oZf43AmzZNdb00M+hKnTdxIEh22pD/rTG
IF4z/YpTwMCrrMjXKBVFqDjtkmSiTj0C80Nuiv+V+6s3reuGC+yhprAT8/XaGPprP4Qv2xBHOGcD
yOjxKjyIGe19R/ptQw+cJWybJAavyJoPPEYxeLJ9EZsDOAyU7EybeC/0i0komiO08F+fkzDD1Yvz
7ycVdTrBKqeakjHlBTEXKYalIzgJ/Zw/PYFVfDA80IPihKn0Z/quuwmCggCB2RrmKH9iLz7iBtMI
stpgPI66iOIDoI0KzvpSKDdN2PmosHopeMNPC5jKhOa65txe4etsxmtDNdv3VJaStyrsD3loG/CP
/M34R6NyvUzGn1czr0czSA6vjVkuuwOn0F9cpoq+hQg/jMJ9AShm0hRiMTo7u5EhJfj2Non6/x2K
c/zq+yAQw0kRXqtqDvuD5OpHD/SV/gPw9U1bxcPNyRZac0y/PDUb1BBdC3A306339950Sc/cqAaM
vNuNxE7pvbrKWKl4AGXRBgySnTjxrl9bFDzA9idqigQW6oNvzUapKd3iC+5XCZ1JjizFJ/Hjd32+
OitV0mNKdLuBc/Wt2XPGTGLeZv5A6+pG1aDZTWxus0bRJunpKwrcMfelP06LAIN6iwVFoPvdX21Y
NELLh2mSFsa2sTcpgQBEhx+sXYF3qFb2qPMarpkvdwkqJXQM5iblGyIIxelQ699kyO6KpibfaN3l
MPh3DyD9w3+AbYpvxyswfI7vvl1oUO1NIbPH01bbT7tIg3kClMpvFBJytKlXKNnnYX5Jpx8u2Zuo
GPHxdfjwpQievcmfsflDy+g3wUJOZKog5rLidKsnOjAMy1oF2cdogZkx7Aj2M4C/ouDSx1ebORpp
DCbWvvvq0LC0W2caLUOeaWnre0n35nQziH0rHr3RaU1gFVHlASpWEZjPOt7KpJ2ho/Bgx+hMxw49
hJLdD5k9bjzzFquTiSDBT0M768IPIloMzxxnfv8aHzv5HqRCcY9az6ZVVtXp4Nv5R1qFodhgslUQ
qwW0XcfqpvtrDPXaTcYQPlZyuTwKxm6Fu1lLlXTxe5YVdbgoJDX/yv2LCDEIbC8wYevTBDRQbBxr
Yold1PmcQcBuHSzwkQs+Apv4uwcaLt4Rh2M1Iypai9O//uSf5JgM1rKKoG9b78cAf91ybN35BEiD
hOeAD98cO8ox9mHNB+7DWGd99tGyewSu+cM4UpQmn0sTGIkGSu8m5vWqGwZbCsR7p4pwfJcpx00H
SaVJMw5qhfRmAcHKY2IBAJqUlgDU7Xgu0Hm/60q/9Q6cjSPeusbNNHYhAG93G2NcW3j29jMfwD2L
WTrazByBq/YZFrX/CGk4TVWmVWfzks/xAOSCEKYpzWcriIF1mVkGjZgWmG4PkronfJ/SF7/E0PBs
inY+zThwOuZkLZsejit+5kmwQ2OG/0uBPCg9V7OU/FEVSdBUIXM59IkapY+ZwR4IZJ2Yx15ULoS2
TZb0I8bJZumYTxhHkkaUW3hffHWX/y2mcb1qVgmZ81jsGSrzp10t0iEStpYYCn3AqVEumxDjumLZ
Mu85cS4JT7PV1XYuOehjgR/MTpJpTAvgx+OhkFEgwso2jTVQzb+0BvYJYGc2N+NmUZm1xLJTvF6I
rClqmJ6FO1p1TKXjmihJlwnPKByxBVt7RG+5lEdoHuM3eZrDViWpF2zT84u9S72U41lUb5c2slcy
np6SJl6ogR/9pUZmJFpa4trezBc+UzRt1tW/RO181fCS6klQqZ9VxHl+Q/b6BosottlqUNSGFKDF
2CsmvoGM9Q3/r/9JEePismqr4Pd4pKZOYzHs4d/z5smTg1taHxhkxPpL2RFrhuv4bxKc90/fuyvl
0+vB7tqdL4RQLGc+haQZevv/W2VA/qCO+R291jWHY3MT0yZ8xkknZYu53mFbTDMF93TkVKGd6+fF
e31dbOlsaNZeLrquw9uxfn6hI6k3zl7EG1rdvBNCcGbdSyyLBx1JXtUqKwfExVl0NjsH3+hgmUZJ
i3IYBzGBxVHci81fRle0v8Nj9vQgASSKSRsbp947BaWjwz338RQ1A1YWl1rh+xZZUrhw9go8DGb4
0GFwoDnEUTgPpjCclezLBsNY+ttVMgdjuETSlGS2U0SQv9aT+MblSGJESaxIUAnnrZ/oVVLNfgTS
P1sZYo7rkdx7Dba/hfZxc7/JdkF76uXOHa21V5l7lH3VUA/BmKbTgKPWF1A+W86BILGlQnSCvvlb
/0xpPQWxB15DfB0OzQTeTbTE2rXSvzmR6wbcpD2fQRC0bi1SxXLWJ3nobEHlCxwXyu7r+M7U2fdt
LoYV+GnO0VoZyHCpwimHvZJbYtxXFkYJDwvcjoI1pXVL30sMxaWtNzLszcMMBU2y5vHZHHCpx3Ou
LYVTNIVvyTh/+ZFS50bbPsbdqfOruojpFdLLBdRviMxJmHfPz3ZpgBtvnBwPAL6vawClrPzOCke5
XN6eBK8pbT/IThLVx0bcynEkXwOzfT/cR0PR+g5sa5HAb446xuPAlCsojquDqiaItIT8mDx8yoHz
MNOVRzxn+1sb+wp22gjwpM1y8BfFEqeVJZ3YSctNBtRmDsvc3owshKlAcQrAKD0S7NFb2zEyVVsk
SjS8xmJTn+ClDBMWdwQdIyAABVw3Pq9SoCyxR+BhJDbV00e80j9cQrYrfElMbzJdfOtnlThqyF14
tYihn4JKhrG5y6quv0J09OKe7pdcWsjbLLY8TO5vJj6LwDpzaGGDa+mzp8wihK973eoQPk83HEW/
rsPl9MiJoETzaOekPcoPLWuWZcrCJcfM33rK2TQLmhoxnLXxEahWEo0e7Y9E/EDl4+JmDb+Hxx25
byn0+3AOEb9rg7P8G9/Zohm0iOPEFA8Qbtv8pQU8ZHJcw4sxzwoIbyCMSZBAKONRrzI/Xw78Eenw
MOCDjbc4e6oG50+Lgly1jLsxej1nqWQgAW3AoqCTC3E2vewrUYLxKKUIXl4Iit3NQFx3c8qwnea6
imZFSinO+HrWUeOrRPmcBWcgppe0Zof6yTebWPJGqqiHVVQ31i3IAbf6Xnv7ZnhJ26z15i9sxvsa
Bc9yIgr/mSusWQcyJlgNktWXARhOPNjACh10A7XgXFPF6DeT2cXNsRw1cKdWVVFElUPaPrJn+Ucz
fmuaUbXPhEro9MblVqEs4gntS9163II+THX1UJuCRxGCTFviYwOlTlnm68KnYkqdY6WPU8q+hHrm
xB4NGn1yrWvYln/N89LDG1by3Qy00EY+SAkvzRCKihRcIBehPc9Ph0+Qu3PKdTixY+IxXs/30ihk
w+yjCNDIIwVnt9wcUvQM/V+tvqzF8Io2m1h4Yry9Xz2lWK2tasEjRkm0KAPogWCvuFXUkFOeme8U
XVWW5BgyApMIL47p19AliEzrLcAE3EHprtu4f9A97zXxln03QmdLM+l68Z82hUAaNeuhvyEjwEFY
crzxrzoYZeSvyGYw7fSr4pn8souEL8xdGjkO9fFUVDBYlphxJbbWbKfih/A6gQKhCBUuPqwyojXn
Vv1nsz6Cc1irNKBotjjbSdK7PpDm0ox1uR/yhEwKi8AQmnfmApBFt3zJ7ogibgfZL8o5eOOyA0Bg
zB6EbG1R28/Tp+/Ic3N0fjp08UCSNm1KMNLq64xkkW8RVM7J8AZYmE09g172t6DTrwRHir0n5EtW
Nr8MbewfUS2P+D6s/CrtQM96ZnNE3So5SYdkE3RXDOF6H2fPLLeEEFjyIqBV7X/LAekYqvSrsBFl
1omWxCjKgbdm2C6BZ0ZSYQgztdNuC7lMOhfX1jl7MCgF13+WxuWWgl18yjEsrxqHpSb91OiMOc5l
mMZHVKdXE4G8XVkqSpyK2WKksnvvImAR3jOUz8JSmmi7LBSA0a62OMfh4B4zDDefOGzqM2glhs3l
8B+Rb+/6tGYOQ75dMUNWvf9evMbNGA0yoSJLTwvy/oaBW05Rl6jVEEYZCgLu7AWAyIh6RvIZT811
umoN06rM5BeymLgcHY1Wn4/MQ+RLTqzxiThGWk5gZZOrfA+b9trD00Xg0g9U9lRJsNqHA9VD4id8
kUVB0TIOirCHHSf3J9L3zRA6WbUN9UtsBLQKyYpkVfZE290SZ1B/XDQV9Mc3PnKgOcKUXL9CHYrP
jXHSwkBSo99z+gbh3n/vadW/rzVFCzgWzRy2PtzVs+/9WwzDig5f2O2n7bxrutOTMbinkcrBMR8r
rDpXmzUH9rrh8bbvmnuUl7pUlNdSOnbaykchepT10yHZwGtS1IHlc1XkXtrH/uE02qaPeBdxOIaD
KvwB/dgIbcgpObkY4Zlx2fX35bMILBLrf/cpO6ppPFalunoYYItn+sueVcxa2vjZAy25siKXC5R2
e0R2BY/8Lg6GfmV7TzbaM5YLtPhAH5nMr4aTsHGG2aXPrHXktmTv/MzcAvNzY3ynMdSMq4v2JTY1
qL+7S+rlQdMT1HZfYEBXIW7/25xGiEAkfYiATk7XkWgE2Yqxhh8lTkvq3sGuy4u1gdtR7hz+v4+R
QqWhXJNgaTRR9aUJkDaC/ypbamNHNjB9aXtSdCAzeG6LgWsWPilUnDWjyr7DaH77XIRIj/Jr5kfY
xmSLpeXl0aKK38uAb/tRmrl1lFImpTMw7H0vUgBK8BTqDwwUc3yUyt6t2fwIthTMphbrGiL4bGXt
o+qvtEfcwGpojW/s4R3ae8ThYpDYNH2Ceng2DDxjSfsEGjFla+N4xPrYwsieqYO8M7qBIBTi4NDK
gTl9CeJz/Kr3n3NzRjfHvroq4K3gaT7BddHFq1NsXBtxMAMeNh6+EephECgHpfNVFK9C6+EZeb09
A2rxCmA806ndeUbtpKTOhbcaK968x/XjrxTN184BkI5U3cx7HQid2HCyK40zKYDvD0NjDexE5Wpt
a6riHevok6JGZt1tDK80AnHvGG0uNXjs7VlzcE+HObrvNHbwhHs6dOAvYyLpWAEjy3Cl/crs2G5Y
jPfj07wZDphrAxaLWGdiXMTVtBhOaOB+d6vxrOAshlxLgGdMj3/NaqO1uKMINzEXqPl8cCGXtBPv
1006xhjN2rDwV6gMsOpnqra3oEpScZ9RUSKvDXdgYAWyqno+oiH41VgS5rVro+WClALey9LcqZCW
jjf3BbRyQocKxFDRf5w3stza67mn4KZXi6GjxImNLSklbli6mbIdTbZnSyl3jxE2RXM0/S+uC8dc
iw54sSheDtcccex2H7tMNJVixkmxueuUUCXXlyjPn3WIVHI/gCKZ1s4F/jow3WbLwQCPPBi8Se/C
aZZEJpOMOaDUyCCQQHO0Xb1mXGdMqAakxObSLG0KuWTZrOr4AILOrHPBOisS1SGcMOT71VZ+RVh3
L1TkiroExBCFvA1bW1yPksopwism6HFoD6kM18MgjgxhiUEoFvWAb14gPrdipTXoc4QsMZTbgE5N
DzgAdAZDPi54n6rpeHP70qYBDPImuC+rHAEaPfOzn5/fVW6HHbKo0iLqEvj9bYt7lTpb6zQRiI9q
AtI39s52qdNM6C25uVT3ev5OJnwqhiMBOc5iwY+E0OqmW+RKhIfleCEWkzEjrqd1woA2u3z3EiyK
ZmBA1jyjqeSOIE9HYp2Vay+RgkW64pSJCxhBn0z3WRIaL48yjr+xrr84IBx/pVDoulddxPO50III
2l+GSDytZgJUY4T0X/KsSxIFXBMcfOpipH/LErWqAhAE4QJCzTlWmF/N9oyELTFAuKGNvGI81TKu
2qmmvZevs2x959T51US7oIxyKOe0IzYlpk1+5qBs53cVQO03Msv+PDesq4B/S/WpgTul/sUDUntf
/gejqRhaNSagDk3p+BZrlSrvnP/JJ9MsmgjOw+tFWF6Usu0PrvhwWk4WHv8IW5qnzPx+po5H8DBY
0GiPtTqZgqtSX3GaEktPZhi99AOxTp6WEusT+CYm6TG7YT/A455kQSD7pjxgSwhVJOYFhLLrj9CC
JHI/awnzrbRgawhYIdE0My2pnrOTXC3fh6hOODLqygar7WoxtpUAxL2VdYTEKKgKfMfgZ6q2c1JC
39AHxsMw/MGhfWuVeQiRiVCf9Uv/qSBEgk3FSl3pbDNq/xHZXdffkCQq01muFuloXYUcELwb+YRz
ANA/SKOKbOEWwa6RHAPr0TONgUFka36TMOaXyOEJit5rgFlDlXjkovKFI/zdbrufqFNrSMAKECzq
VKh7IwAhCfYgGST0e8hV9UJvVC+zLt9jZjNCOaLkK5N/elFDGdK/qfFSpPjxd3TkDyN0KEhlqelV
GnlF6KjZl+TuF3wGnCJeFgu+J2C4mW6FzE/esiy0woneeVBlLB2UQ/hH/YbXVmnKlEQNbJvIwifV
8cTfbxQ9zhLo3onxggfXokw37DGdC9RVqkEu1gir3EcSrcOYJRgNJYCYw8VUhKOqGTalNjEXBHIJ
e1eFV3UWUwOAAM8ti4z6Dn0f+imsdNn6YznO0bNuaOp3T/7VSaxyCpIN8pk26fxVIMZksuUVhOYP
1OwV6m8sc15s8LUE+C7kFEv22UTHiG8d7x+DmWNQ4Ybn09PQUMwvAKB7oEvtMZC2Uc/Wnp29djgV
c6EsovQAFsZ1/UgmJgSJD27MWnJozNl28T6RUFsNiW0kw46sPEMRxpNTAtAsMCO5Dt3bDx2oywca
mFOqhvnRAyHGS3bOKtjMD7ngm/yCoZQ4lFQkNQOuaMVFDsODxGjgPANFlQRDN642q7g9nllFeBXO
5TWC2UgDN+fWOrJdiF21E8j+nf9Bm9UuymB5fn9/uWdNVdrbTXDVjqQfYGxX+z81p2wh8tMvcAdA
Fqonx8CxCKorDnB8HLy6MKOFimsMKnmgJ4Jo03geOTw9YoBCcKE+xFa8DuL9EOxZSrxy+Q6ocN45
Ko05XJj5Od4SKwoWhyZbtwIAWjZGOgdeE26BDzs0nfhhoUgV/lNYY87Q1LX4h1mWulxDTYwueeMo
Cv1q192PuAYXt0u1X6X6v7DhLFihg1+KXgz3ZWxiVuBdOJEgrxsfJ6w0PTc69OxU+A7epSRyjF3c
icu6+5Y+Y1bj54Fza1ZrVam2ffLjXUvqqJoeHwJlfwGP7SOWs+K2f3iJ5AtJkGxZvOO0iXwwq6Zs
wP4dmTMbywYWG95JyLIc8ztOCSDf+89VpswwF1zDHeUMNiX0qmTkVAzOghHvANCz6uOQltz3g5I/
tRdVinwUrOwQnVWgr+OvPv77RGUmQ0Px+TqlqbqBKg4O9EnU3nS3l/DY7knmblr5qJnKbu0k1k6L
MNeG9AzwZqwlhkoBLDi/jDZNaPLnCceKq178Oi1eiUqW1pu417uyLVDVaD7LPEtfjFLdg44Ca8lg
ZpwWCOi7v0FBLGXaUXit8quZPUpaSRqJXpIsEgHG6sSfgX2zeveZr9y/Ju6CT5JSObt7qX76CLJ2
XMYHQuN0zY2fbgfstzmVfbTHL6Wk0TVOZb4dnEidFEj6gSHM0uEOjH68BLGYy+JpNJxfSYKaYFGv
xKyTB5sSXxiqvxVuTxpqfK9Xb0crIH9GDgQtYOr1KmAzZ3VDyNAlsypxN5cjPAv85r+BHkO30eKd
FDLcjqNwEdGZMGHAfI+lZwJ0BdLJ9b0BydmSX4oO23bI2L7nrflkiXvY7JcN3GkbkgazPsoZ/Zci
wCcRyBcAnpkcc6v82soDzVpFejJ3ksK6iNSCiEQBPHAiEPBVmRGC6mIJ+sQyBbtUSchtjC4Yr0yc
gDhpLQRlmvx2QClbD8E2au5w+BoZwHg5yZL74kLsvrEJkjQYiGolGMF/toiV7WwASm+HJX56u1O9
AXg56Yar/ZHe77nynxQ4wBM6kS0eOln+n2PmHhH6HVxf3xIhwcpRWeIxwsNmacDEAqljNPJxHpbj
f0CYeQM5p6SpQ1unYJ7GfOOkaf8OoQVUC0laFg8+5CCcCEx5apDMCJT6AfjyD0hxx/AdNahrViRx
JpHeE1pGhNmpfS7bxzrkwA3IlZjw10tFV9Hp4uDKoMJqO6Z6ztlYg6d4VLjOYvxXj2afV3bN3IOL
42pwe4XKkIz6/D7h75rUfZETlE1RlXwsyB6d3naT1qM85h31pJdM0W2W/69nTVsuZYLcNVs+KW+D
c0pMylb/woWyMKBhvlu8xBKYHOZQjHZhIm5j6vhNnOZGpLRRyRTxmmyNO5gpYvL40LWRpdHqJEOy
hfWBKhhPvYTcuf3u7W4tUh+cLyk5s+Mm25gqSaX7iahWhkm9gIs2awiaUF7CZNlQANkTRsxPiMLC
V0wkpdZVaaA7YT+q/al4w3ld4ZPs1V8ruwYUUMVjZCXM5D/qc1lQ7WchYTzxYLPXu7JQDsj21wUX
6TtzKG1tIFt3pfg3DHQwEv/BODCMqFhZQ0KPw4GVOva4jTfN8IOlOUL0O3OlYxXOqRH2L9aLkPB5
U1XEZsarv1noqYtk+3j8DS2Cs5gi1G1YSLsmvV5w4/l8hoQRBJBF6LDYA5idtuvUi/XE+GnN9FBM
DIeFX5/fLxRGQb/C3gFCJmN3KzTS8/DlhjQJzikpHmWLEU3FDh2H8w40PK6JnOb7/1eFbs1LbHju
EkYScCW8bb4Ntz0QINaTYNpAsslYUn4RTRVkqzOp5GA/QVhHmrbrYg+Ka+gE8/ABcPeWZjdWj3Zl
AJf9n+9HwHiB1yxCnBkV2luw9QeLm8dw0tfzAcNguwaVeoAwe8ZHtLKGgJbZ5bNpvey6dLjrBvux
ph720JO48W9OeEm7/pmHyBtcxaA3FF+0qB9q0LCuSSXpnbwWiPtLTflrFGBgUJVkZGF5aGqKyjMK
6Fg0OuvAtbjGBi9BO4U4mb3mm2VfYFam7lokKIE8QN9Bwa/EJ39oSkMjP1aGe6vRrFhChv28zMpr
zGK3SkVPG05NqjQfOJEU2Tpr+9hCdJBF/Gurw5gKi0rbL3B3MDu3kZ1i9X95e41VUZ3i12JuzJ2g
hH02pxU/6iplDYTWGmq4elmwd7clbEbewQpZYpSt1KcHBFxVpja7EgZQlijce3RoPWByLv6YAaX3
Y31RBtBdeE9Ol8Z0GcK04GDPx/E3aCTW1ler7lDsZY8Nh7mv3E6yIuJNkAVqrQwm2/4AcaV/ZEhV
yrL2QOk3MYVhFmWdRVRqZVFR3FPZQKOy6bSxjPBFulinfio9PLJBMgnxREBhpkVyo9Sr485xSdvm
1IlxWB7Z7CxnTVcOSBYBU5/brvgBJHMoBwrYsRhHOIoGhjiGg/JOrrKRjZJpPjMChGPLvxt7ocxD
j35wtET08xSzIxkc5XxaUp0bAKQyTTKONyYKsRU5tKK9zHVHQUDEDRkBn0KO5zSvp5S6a0Ty7EiW
jW5EHV8wuvjpuhmgp8facjKIUNoUfPWb6voOD+lHCcTfIOFam1jtX5+1P0WJ43xkkjMrYPXko2xL
aMPRmxUTLKOsQQenhxu0lkVLVnyVJX76hurIdtgS+OS8jCFdV3PQTl3Nn6E/wvwo9+BZP4p3zaaB
b2iUlh0jotZOGkFfPuGMDKJeNyNKhi3OpdgHvscXxw16oKSxGKdbfsOs0mn2fZf5EvM+admepxa+
lfUajfVGPLRaTGOWXSbaL6ogm29UnETrVdLXWITgaY5wqb4aQtMdjJ05LQoLuoHmVcAfrHvmB6i0
jQgfB2lQp9L5N6dv399ekrno+bcw4wAa7ZxHeUKw+J5rwORf/ZHVvwgbYjQKLmruXm2aXn+hT+v2
JX47pG/6W/vzCUuibrVnPMOg2VRihSchGmsAiMWawrWku0UjCN3zC9jyiXUlErIFfnLQevnlzVRo
wcHdJREqQDNaQ8RbbHu5oI9/6gdzMHSVDzSCD499KwGVjlHbuGSclYKLLqd1tsoFRz2bnEsUQHnn
3QMmhAhyVEQzHe4JEiWc39a8hNcb2VrNgAAuoE04ENhmdTLY6ChZ7a/2+IEALYZ9QyrqydXPRo+F
OGdo7oKFJt+FNVFJ0TVLH4AYZs0ruaiQRrsQlQ5bDQNa7qfsZs3GWMobbARMmp950DBCAc67wsQj
szsCse3DkwVh4auWR/HR34C5KcSkJmMwN1vw8ZQ8xloakinvnUxUmof1lbfYh78wNhGFZgDhXO/Q
kO0NoDFeWmzPQnMZGI9a2TXue02auCzf7eTWqpK3bFGKChFACmGIywk2rUzCsXlgb0au4D9Mb0Vf
GHGyHnS5S99Va23nKQs9mprSLJ2u4hm8+EFThegJ6kM5jT3ZRzfL6KlwE0U/GffljsZG1GmMCLYp
Zk8ajbJDEHOttCjuAam9elLbrce3Cbcs5fQ/3G9cB2RMdzFUL8md+h00xj30FSto3WQ2UTM8TEAY
vzkm/0t531iLls6pSW3IZwLxV6nBEoSuzxDPGNAyHCxuZFExgAsaIuwgoRQOFQjokb7P3doYN6kU
xs2afLTnSIik8oy3YLAj0bB8yq+TJlKZmDVWpM4bvYhPxfud4S6gx9LYeijRzljiK856sFeHKzBZ
MNI2Vv7PrxzSMhJui5Q0EnSeSPTNVr4z6bdI4eUWApMJO57IqsAjVfuPX+dk2pxfUP2aSnaiPnE/
Pc11OP2pKTo5KZbG51UHMg3zXb5ifvIvBlxTmxRC2dDxvQ4Tgbi8joMdG2Nf0bDzJWyduBFpkcNS
dLgRkxITufScNtyvmZbTWBWnOIOP9SgZGYCh1Gx3foSYvfeSWFfS3vaUdiQIGVYUTnk6t9lHxQ08
k7fWSCC3v22n5r5w8pYLSC1cbfM/gIJfNzGiHOoKZoth4CXVgTofdTATtCAWHlw+zPjaV5uXdWen
47V48N5W1uSxCN+ZGTlcpBaBWOHo6cJkE5sRmKUtE2zSvjRhLfoBQ/9HimlXZTYpdVazuQ2RxbVZ
soFVF3L7RD8ldrb8lp6O9aFFZx3ktqDERda+KVJu+DPmxHGRw+t35AQ6TNvt6OyJNQWI7Pu1gQkW
5eiXqZjb/AgySB9RN20W4OHkkhlD/yAr6Ee0kFR9WPFhBF976LwlZNiw/3fjssrVQCYzmifwHgBa
48X340ntroIpsmabhfW41ZMEOXyn/2ulO5CG5M/LBFlYKE874f+2ZrSqYCk4QdHNH3g1rAGeFElh
fbJ9zWRQV5+n/2dOPTtDThLBG8rfA0eI8ue+ptFEllZZwhb1SRmVqAkuJ/3tyoOyLMjUnZ2dOkbM
nNX/NHzYGDmh7u+5/brZ7Y9IBbe1gxkZaavora9PPZv+3/WBgjZirgm9ENtX8n1rW7AACoe33KBb
4NkGSE+wckPt7BUdE1U6B/laac1TbC61f7szjlCs15K+XWuMrkr1fTELwstpRL5RnKagFigNwTMr
eNbPDKTeBuPmHSBpnqxA4Pjhmk23hR7/AUKqZDooL8ODhfHTvQqB+2F5EojU1m7mry+z5MDFgVVt
P2IX35jm33rw24FAn+yZuu7rFtW7WlD40ttsvTA1ezGvab/AwKVQW/DEm1HnwseZYuerpNKhPCNr
3N5NalLpA8l2Vt6Y8Zcp3PNzmyftM/YVrK+dTS/i80J4jkwQGtxW5127atznV/lew9mFmu1A7n8z
KU1TgVfBUojkySyfA7lJXQuHrveXgWN/ag1RkftWfdxLv3GjSzeU2awjqBTwZv1jfeQebu3r+sPm
kM+x4LF6Yy8IgWqFyJLL63AIGKs/VyvoA2wKVy3XGuAU/RloAS0WZCTSI206nAD78/900Divye7U
dubYt5f9MOJA45DXkhjDPbHP3Sj3KYZ+Q/5S8QZZbOJmWy9/wcTaLXCUx3w3Gzr8gInUDqEGSJbt
mmI+BkTsr8w+UCQBQULm9rg7ZiA7EE5Dec/kdlbSfOE22/6ZU6QBNw4zx226FIALjBfuc6JxGeeA
2Affp9kuozUtqzmohqHjVlRq7Hll/skG4fgtHdkbQFOtoBu5IsKC+DjEeeIp4FHUUrXa+xG4E7uZ
6BBv7Infy8kp/rscjsZ/bFBZ+m7YxR3NJPcj4hgbVkhcxBqebo8KF7XxOQgLex9vLbee8DWO5VWJ
80g7cxP0cJjhAfRfZru43FvYDv7cnH02VbaRMVQaO3g2LEMVOx4TJFHwYqnwsniSK9cP3i0ymCQv
Q3v58ylj36J60a5gnFHYZsbgmRX83h26GCP6a8u4Hh5Bxas9D6dCcqSyf17u62Wn2tmuZ5kSvXlO
GocQtQFtp7zQ5gc09OD+wRxg/OLrXKnUYy6CXCulFLBKPGb1Jl4YV9PqVf7Tpg5d0PiUqbiP5+tp
Gkf3p1K8A8HRjlQZTMUEgaaYvYAscgU7bBWqeGiWy/i38ApUZMwaTMsBhu2gC2lkWD2NKpPImgRk
iW53qowhRfjojEn15UNEr6gYYDoCKH+KSNqbGXjRjq6ab4H7AOfdFHCe/LMcdIUoHZkqef+rX6My
woHnL+thFuZkkmwPgpaJQpmYiti0BQWI2n8lQ/vzE4epI32G7oQMQtqfiPGUVy2Y13ZjB+VzZ7nA
K68VSNzeW5rGlAY24MIfyFpH96/3JdRHq2zaCt7x+fG1jMzoDT8ob/X29WP6kdGh/jhnbvPD1ZXS
sBDFYMtOjCr8Qec+joY93kdnlIX2KoiXfXAhUcdX3WMIp5anU2XLIWRli/E8rzjsxkzhrmqk+DFw
D4XgOIuOb/iPbFNjZv5uzL7vdnduEZyzE7vVWBxB4rPZZsCiMXUGreQ7rUpoyn9dsvgxKZPxGzbk
gKogF/BDUYOaxBGJbu+Fo6iR33aFMX9l9DuX/DqAV8KkWumzVlcpB7li+lWvEYcMN5b6loIyLCcU
Q39Uv1m0VPGBxQq7BdPpp7pSB6Bd3nGHoGRlRbp8nEnqg37PEMNj/rWDSR0f3PGZq2RbYq10hGMg
MLfI1SDYWn9QLKEemwe9+0Yud0Ab4qaWW9EZ3NmqqfE6+BITqvZbJn6EhZ6JOQbUhWEp2bUF+7ZY
dL7XInNTVIeVfvehA/yrU/iL78yVpSTwhCn0LuAX6W4R+xs3MXRYwOV9ns+raXVvoEOG/RwDj0SO
o9SKwlXHDBo0mIsnWQOYcvR/1TgCihP1wp2eQxXZlzdRfcheTQxp5UAIIeblFJjoM5CNZFKavGNt
Jhb65GdSSzDVHQn1ZkJk+oxx5pn/j3qzflueRZZ8+xgIv+JHMCBs4NRHjmpd8oKI72lXfJ5NkWW7
Vb9zVui5JiS9I6baf3TxPXuaEqVxMU0SFxS6ubHp8gVO4EjNBsEDoB9zkDefLHQ7qGKDwSBGvqsG
6O2/+FimXNlS52Aunlwx2omhFnB94z4LJfl6IeK833ZhnCqbr0xTPhFchKDoKC6PcoV6SMllr2Zd
tqqOdgMnmi6gipDvbuVaoNbOeIa7Sk2yQnH8C35B+x47D1QJRNxZekOuQJsLp6897utWqoQUzcJ1
uPhMVmdlE2Y32FMrDsaYLCcq0yGoOuqYcEc+aYWWXZRyK5dabs/mkU2DBkZZR5RJUhkGQU4c3FJY
j42wsVDNx+R5WwjGrxZPw2nZ9Zm/Kj9gpPxi/AdK/Emg+w/eqiCrHLBYxQvQn4ddvJ8k6L3Peiou
8OGnWuA+oodyUAk6/lQ2lCQ0DU7Lz2ZOYDr5Inqc2sjPMJT+/EnVhUfTdcv915OQzKpXu8oz6dTH
lp+5NsPiF08aOgx5177kwX+f5881nsZeLxpVbWNB5R5ayVALvywKaDPCKe1fhUd77PtH0GOxpXUa
umMt5uVI7thui9XEjv7Fzer9J3xzRP+Z6gU+PKpPl69VrEHrYuDtR4NhHWja4TK1XtFe8kNatJRY
g5l+xu33LOivA1mHB6Y+HERGTVhhv60o7PhVCaMd8tX+WxWrFAWJtjWxNELUTY0Hk0H22mMp88+5
1i/GRIE/mfNRf7juEVGetNFH95kqIhaFV2Wbm8/s+uID52h+3yFH6gQNbWVjIqhHliNtEUUsyBv+
xIGrR2Tdt207qLd4kZXe52jL334A3tQpyyc+YUKYuZnxi6buHEWFcZJa5nXPeRzbeZHEz8vEMBoP
hbKqkod1xB7tqZQ3UlBv60iuMPbE02yj7jG/wtmm8gJNyX+u7G3x0spnh92JqYAcwj9acvxIGeBo
bkrhx1gA8ENBu5woTsvvLu8J72fHGqYPWzgpIRVRUZitKDO8Xomiw7MV90rWpwRVyClY3xnY1jcS
u30ciZo2zVlQiWeluQqFdgcTPviC7AElM/xhHcYfpw4zpzXw8XTu47Z4ZzFE1IWdC5vnZMxBbHWc
lKDsAgYCoFdOEiouNrrhZ4zV27Pxk9Nnt2b4ZtuGF4EEjuioF4/JlwGci+Z7dhFPiZuYap0Jz9tG
11YYG7Iqs0v3qT9wG6YgZQ9TRNVKpmAK07zcdl7ErQvQWJhLTHM8EHlEIuKk8KhTRXAfWaWoQUrb
6Xecx/G4qlKzGoNLJZhevYjo/tO2ydf+HLtgcLwaC8hIS7AsaiRfFltVurOasCGbPwjaWmx32D2o
wZEwPHqU64HcmcyQchUYAE/+GGTH53JqZOUB5EepoHRxsf1YLSnnZsjsKy95ix0ziz/EYDqy9uFD
ulADEa1OJ6Gs39+6jbospW7cpe2W/wTnHvz3BtbqQXhNpGo7Fp147dehKGYsQsdaXhODyb/GmevP
PNnXvNuJsd6frZm8/u37q73reFQ+eeSCeDt1ULKEc0nHYr8jtKyHsqigWx4rSgbi5c9ivRQzV7fm
Z31shs5Vs/Nn+4TNZX55pmfwXfwZvfuHY2jfOwfpKewes0Q9kGkZPrI+xJnljilsmq47kIQHMVx8
HIlImRwucFm7BpP/X2tHQTZ05L7pm4DvGCKp5b0/zILuDPoQ5CaoN1easJIAy22pbRHWOmVTprGz
6MNJL05C3cSKefaDV+ixx5V8yUM55p/7p15JAlBtjwOaVJQDLjBnFQNzldY4WSKPq7h4w8pZA+4h
cPdPR96lXeksXE9cYPA6wUe9sWTObUWeBFkKIErfwGGW/07xTLLi/0oLq+gU5jLLgabK4CEUl+O1
0x+oW6bMm3ZoFrvzy7qNZOi0CHYQSFobk3OJqcrpUwHuUp9gdGmLTGtmWU9xALSjHAO+BYUP1q9e
uUZXDxMbXx2oe8pAN1f+7WWPjiYoJH32QOybAXJKAR550DYU1hdHj8QYULsluRDWFFMHpflNvUHS
W2f2glUIXHwBfu8FFrOGiNCXwXYquoZ4R/pTUy+7icKUdZ1+dd7I7BvbGIg7B4etMYU+QhytBjcZ
2i6jDz0oOBeS4sQu80wzqc0CEs4ATWuhbZFCrmBYtcTX/4Tq2WASBj6c4EshFpqQM61pn2xbb5ip
slhBZ3pUSTW7M20dRLa4uxgERLqXA81ML5DttOJMRL353WiTCIR7wYWFbH0Al+XiMfg0LvlXQp6o
npuZG7XbRI97xdea8u7hme8HXvUzIkIppoReuvyTBXl0pv2h9P39+GBuVcKAebqggdfsoCvMYAhd
tcO6GYliXSlCuW4l1d8DrlUW/Yo0XeTieWbweadmoNNdLIs/kfaqCDuBsp8fStjvPlqed8SnipS7
+a3TWeGo0I9HKeQi6vGJDM+q1+S+D3pvoh0MgDyy8JGYUVrFe1do7BECxVc+l9Y0H/gLIVAO+Jmm
+ZEMwqp8S5Q0wgyhVA5clDkMjEKBunJVZZIzh2pIGrHCB4eGAItEcyAVq64vCa/csjbJNcAix6Di
u0klWuwEFWbd1PrZ47MAih5cElb7v9vy9y03Vjs+kqQERB4Co1ZithlKD/EtlSsdWVeAmafK4T4W
VR9suZwtNc16Z8FCvPxCxDbWuEAlxDJC+u2FZ53fGvmKrYGvz1SCpIYouamEJsxyOXjAsJ7Ml5ur
oQhjfzbAwlLHOzDOwZLFBSmJLRzSScgowoBLC9yOswUIoFgKHFpr3otdWDACeo+zVXnD7j4Tp2W6
8NCP+8MuySkbAaHRB2F+Vvo9Tutiq7fmfsG8bZGv0jx38LeGLR9DTy103ZIhXQBc1VtR2anz5Gbf
vQHbkxxu+yjSclleSP4NtM1j041bDWR9LNmo4S9zQoOgRANJJ+7upx6OqnVSOlsnsf8WsQrxuSCZ
HANVNuMx8YEuFK6P7Rfjg5SrOBf3pHevaDQW8t2k+xj/6Xn+ekMPDStwxOKIijKWsLrpWWYjKb60
BypgonoSK2GglVNaGfNcyvN1t/6Ct6R2e1Wh22cLKdA5eeqGZQNjWqJlPRGdxR6nHOL43eOWxZM8
o8yTNVOI7TNiklcOBME4ZP5mvKQrogg10mdU5nq2y08gWbh6l5wtvCo2fQkmjoGdzegRGbAnOOWb
Dh/i790PjY6UigOPRmxUwXq8jhk4LoGgzUZ0Fcy6CcmjVZMxIyv/NR7n1js4qcXSLricxTI+9Wub
HdJqe333n2gZQ66Is8gbeYCl31WpWEP1m91ZdyF6hYB5vB2L+iALiwtIXYjtBB8vntvHZx2Z8cWY
YVI1t7GvmESIrUUXcBZkKW6PUHc9F5f/phnaHLG+tgk2153UKDN0vgwRZkEQ+vpJUHMnUmHPgUmI
yxD9LGo6Bd7brtzx/d7MzpfzEDowhfmUzNHvXZSmnJXC4ZyyBs0tXPBDU5FAJgM8NnOPW9ixxFtc
/4tc5pMzycITgqi00+KBbOl8x8tTRexBLsEC1nUUGHXvXATQisJ+h5bhPqu2ZmPVuSMjzJsKdCG9
7/72yqasmFxLDuZqbCfDxUUcrqwdOoV38HMyW8PA0A4I9WX90XvPOHTcitVm9sKdLN1HN2I2iDyO
cajO1+S2IAW/t8fIpciv/AX1kE77QqbbedGjDpN9zoog/+zt7nn1dCdyB01yyYhnq9bZrcYcRiEi
RZcSU4ETqTog4DCX0JMQ4TohCC9Kc2q4hL0VWir0p9zgYBsEG317lZFRqSv8aLaLPaH7VpwiRx2/
GwO+8+lBfRRbgvFuYnKKlTchOoY0MhaSHiSHjHP2KDDTcGs2qiI047IftVrSsStCLts0fcDs5VmZ
sOtOFZ7EzTaTXiOI80Xp++7ktq3qdp4YRO/3xV12lwJ006TptBV+isw8XzSp4dIm8J9ZbUT3+g+Q
S0syQlIg6gZ1+66OjVRhm3wXE+NLolGPrMEnDsKWWuuAWBqZJcc9zHTM6dB2Ctda/VRy7U43/yIk
VFe1lU5bOZmrsxoMn9//OjVGQaSnZNUV0eQjtkWs/Bw+lmKh+aYi0kd9QbGeoWyLkYXQzaw4ibS7
MSRsfz+3duZskQfGrFu9si2YfC9+1pZXVIoIb6mZzXQz7guVIjj/iV9sxiYyEAgB3Yor+vlss5Nl
SRqjPqtMvvVhPRp6v2htbB4lqLxrZqnN9a4H4vn/IXhXmEd6urdWSM5A772sS7JmpEJ2NVZ42mc0
wMdBN+hyXpbwgpFua+wt6A+G7mrIkhAIVdBj6VPgPlkSNGHSTf8Dtq5OJuWk9mSIiwGVrN1dXJXi
UnB+5s9RHxK0ZEDM7DIW5R9YCHG3zeh/l0DxZd0Ep5LtPMgrdFfMWKQxkfZCmSjngUsCYmQzVTBM
+mXzHsyyR0X6k50XanHDeMw5PkWIFlpMudGENr3Vuj4ozmrwW8Ef0Hh03CB5WpIBk96IRmJrdnk1
doFaKsP/vS95KF1mhHzTZnFq+quuaelURab+ThoEqgR0/8fS/mVkwDBSDLQBdweynMiWIIOi7DUe
dzzV2FsLwTrtR2xq8UHV7jE4Qofh1dO2rUjj2WzdeorV0zCyVbgoH/dNAx+/rJK2zbQQckDmW/yX
6nS2KtIaRj4S85YpnhX/ajRBZqFkqJ5ooTPsgn6bpq640p5sao1xAgjLnhrwYv72KXdFF3GVIvSS
lJNGpYh9Dkw9a4NVy91Lu4nWEBwJ9DDNQ4sIPDkKbAHbaql6Kaw5jAnoNmqzHsPeI4A2lWov5Uw5
yfpJdBKqFm5pKJEe8DO6FzdZzJbopn0Qbq7sbJF1l+FqLOqVuoGdnzMA8nEb5GxGXnltyE3tys6B
Xmm3D8qdQn+ZXQanAkcKuUZEjjH6hc+hssfbYQMSGnbJ5eQ4pHaKuiyvpUnH2Sjsrw5+DnTY+/tO
koy15ga2tB5Dp2TJAniH9VaCtRNkspyDonZjdv6Vq2jKM2NlGwJBSy7F7i1nEN3ZJG4cootWu9UV
6pe0HMz/VaCZSUagPIzwyk8E8g3vbkZ4gtuSFC8n/4nmiMeHQ/9n7AXx9Es34zn5GpfDm3wdsdzh
mDWixhN7xjG4k7OD5p/dML9Z1UOtSWfQjmnF46Kh1167nZorEnrann/xphoKSEu8iOw+lqfVRtWf
LEroeAUDN/2/Qwp6aKsISXsj+ZhfYr/sOm9ewcOic/b6R5LA9dbvd7jQ0jrBF+lZbJX1z4dXPqRi
5TT6ZOMG4N7sEgsdhQCaXQRXPnFWIoXyxYp0CZBKWWkIcYiB31FtfSo52UtcGKB2+aYgLT+2XFP8
iCWdLr23QlosT3L6736MWvyyy3K5PAjLjFVZZbR7evVAx3CvhWXqUjqWgJycvRHFr4vTHmLCChwW
3aDKOWzOyhOAoulCwBGB+SCCuHMoigmya2uqtyFOqKIpr8JrdiC3MhEdDLF4EOShm5bbn1UOH6S+
M10gb3XqNrCkuVuyR/aCuy9peQlSJdq17FV3wCIFWoRoiFagHe2khf5esAtlrP559XOJsZ4aQw73
E3UCBdSFEiGS05gpbx1tWPePXg4sdcP+f4dM6MvWosGz4ISbypOMvk6OiKEPMQ/Ctc7HTfpO4Ot0
lBNqdprfyhSeJV7+wlHXEozh1qFKsTTUVr1mgiJUoMgn6eG7CQttyvt/mBT5OVSUHF5Zifbmd0is
1qZbwIlCmxzz+tixoSwR6LH6E5vR5YJzWb8nGJ0xVvzwSsHrk9asnuf6SP1SV9tH9wrcKSF9FBmb
MEpB8F2uK6bbJvNbGSNBao8O5OY5FVjJPQmqvrM8yrSgMjDqjj1G/SUegpv17hfVnyCwpuPg3510
rc5sjL2Lf/+rounoxOZTahTDq5EAD00D6iWorcv1mi7V/QyUN744Nrubv9iKrSEaDmksH8NaiTwd
4k22cxPATxB2OL9ATHpWXi9iOe/8mH+C9SKzCedCTfInXAOB5DBjsGwLtTvjIyr8cNbaxdr9cSWh
GDcSGA+lugsRK0Io7arynHsEAM7rxkczl2sKbS6E6u0kyk8uD6PCd88zzSA8jpMIluxiV380Xvpk
9OWA5Gn4yEp3q7sJlQ8EqWZKedjxEhmYXnSXRxPG8sMDiBt0V2EJSYFSaFc8fHjxG5RqtjRyz82n
xe8TyM/UCXg1AIDtBDzpXqpz7UHuK/d2zHomil1gBPC7JsvYdNvtBdGmFPP8tcojwLnHYG4f8aFb
YtysKe94+1AtA9pNvC330iMAEczu1nlud5JZZTuxtjr8znWcKoz/i+0UByfsfWjqN7ySDAbWmEWQ
Rgt0rFDDCppaUFdkwBbEBIkMAF/SATYrOwO5OC9vucRx/0x6zD3IW95EZnmz9hBv7QFKUAY8Vjqd
NE9wyC0Xk/zAsiYm54BdKUmiWaSmFbo3mEQmFniVkZyIigZPE1SalTKKtUELtrB7oBX27gk3NaE1
Lt1sahzKh2iEed2BMWCEhfSGCSohJubfXOmGIOUT5CGPgCvB9OHpYlgfE2jrW/55KikkADXSFcP2
FXwplpZcMpGSHED99WbgUwDVRwEf3581q3Rp8GvTDhvkeVtFp3ozK2qk2Gt7f/B/zKZ4DdaHCLO0
Cjt35rEPhN7mURfOiDRZHn3colb1BhWtbITMv4IUZQt8+RrGLoOxsw1TWUHuGn5U9GHMTkr+YD3T
WimsTStLI66tCJ1QGF1JKag48ZISfUWFRmiAsOq71oX7MiGidFjmOSjDdoYzEhaD/cAbQCf7zSw3
ZFtV24fowS3qPjGXSGwbdOc3lUAW2TapbeKN00Gf/s0KmDKK0vmBhGmZcrukLogzA7vSzK+F+158
l1cRyrr/K+/ckrcAPHOYLYTqRJcBp+d3YiFX3mqg+h/Cd6kKyDHTbXCDoXU+1tpKBP6DikMFf6VE
N2qqLAnMr8fGQd7ScqenAp8mq/VjQ/NWEW7yi9LuRZKNIaEclRni/uZA24HKL6rgOtV8hXDPWY+u
50VQkzar2p5qC/Igp0drFY3xMxOJXKbMqlEgIPBmI7hxUzhSgD1QWtKecpR9MLVYnBulUaTmnEyb
vDV5jm9MJ4J4/swrYF045i4U7d+OOEo+VvH8qZZmc6+ddjm9WgLbvSbXPkvQv8EygeILr1iDwiwl
b0imuOorfC8cWHkS6BJVv37hfyTBjMnVEO8ILii8BcXRiKFXJbmzc6f7uquTELEB8J7kca+GjK5R
fCTlybXqOFggWOXiU1ewUBuzUn/jQ/CAF1LNyrUbq60OzWieMgfCgvQ0KP0uNTqHGy0gchib/qMt
ko2xrgLxxIPFSCs470/scjk1yWZT2QRDlUfaB/ICedk5KyAHgc9gyDSl57VxtuQHmKrlrCLAvzYo
Jzd28roZodTMMQBCpIsYV/ly4VFQa+zOfUUhAWHExMeYMJt+IiwdIb7/OyDprOMo3/gMlJ0rQfOp
ZnnDP3HHpViab2s41p7AvEKgXOoA0AG9oWwgWK9VlmMBcvwofAfCrAysyeUmGaso3J3pRgFKSQpE
opq63loGMSC+rkmN78e/2VvgMflUkXKQuRXpAW/Hk8T/4gur1VR0SnkF4/PIlF2llXvAr4zRuvmF
a5ryhAQAqLl9/Ucw1T1DvcaxNUNTIqLfITYf7cIDlPn2jutCMtdSBqlVpgDRxeRWat/h+1uyHe/C
56Wzg9Biq/h0+E9Hn/rIYy/5G4dkj6kHX1ufcpyZjeiqW12iUFY08gA3KQ2pWutnfa8Lg3KhVLJp
0U1pKbugLkcHvASoVaCaBUgAEhGgrMywW3T6aKJHr34tDSWsO8VauT4MMoDPSwmuiu9SIBiJMftV
Ry6oh6K3/Wt/aFjLCtqzV9ucxsCF4XjcAsVzoFx0JikkBoi+pzPluWu59znDh37i38CXf5C3Bk8y
VQO/yW6bn35dwCiEBo8iA485Cu5v67lE6BOsUM05wJ8XV3fNbQTCOe/GYRXlNxztzuy89d8wasM0
SQyCGUGA7YNBVEylFYci9DCahOu1yyvVbe0/kiogc1fOJ1TY7Hk2Zb8CPD/IL0GPejYeCkBHRTM+
qLvvPulDZyfBuzDcsIM+HL3x94IalHlWz+FcgrBFGr9YrI5zfCRHTlU9vgHD43uRVN9qwgPbJNU0
B9zEkxWFXrQ5qdcWwjznnSDaDxHqrzjEEytJgF23fBjfSFR+JvAo3HFidbXy5z6St3Zo77C3Y04u
6JWPydCXIaVfxGwkbfsXD9zlHbAirIoLaCsUy0qgpS17yMWvr7dpj8WZM/g4785YSFIZ1tngSt86
s6jgWbSKe0c42MS1KJH8XpxzEyYHABwlzMfGNdrr/i3Np4bYD7N9sSA9l7axq0qsoGFKuirAKsCX
hc/x18zrJ3+VidGeYRMAoLjiNFLVEzv1xNJBaaVPMyss9a/v823P1M6G0Cz3wRM4862WX372GAw0
0h8RnnP58BltqB1SLdqkcGeu04ZFgpQbokp62vIFi2ZMhdcqw6ijpODepnSLHsKM9CBKrq69vS0U
s1xUjXPnAV0ghVIEpPajDOpfWTOev2ix2iZ6397LeAHc8K8M4KOXcw+UyMezkufUoFwsDMKRdgtq
y8KV4jWlYXo0giOigrSnaLeiiPkWziVVkGMJSCmUg2vjsgqDNtsTdVWcc4bezjbNsBK4UqGiRuws
HwWjYQ9ArZmivVz4TLavPyh4xeQ4W902IYMa4ukqSwbbqCIn2kg+mDaLdww0X0zcnEm6/kCssxKg
YKJXz7pBXhD8qdpPsoxbKdqd0Ukqg7V33VSwa0MQQFRLDgL316h94TChILVUJGOG7ifK68mXUXEm
9Z5GrwjHWaoX+Ryc31xU4gfdjwJrkICt9G2ncuuo5FR4APuociVHaNCBMyH15LHrz2WPFfd3PE1o
onmdwjZ5d6+lTvTsx7t0KujvudGfOAWjOASYkQEM5h6/pWSxu1yqigTpaxwVeca4gBEtH4jHvAGw
R9szT/OZJ5QOTgI99ot7zqE9bQ40iNIaDsXlzRZ44IW/oDmhkCVGvQJKTsTr/B9js9R1gF9xrU6L
PA8/baFmz8SxgUv6MriG1W7g3jAjj56giR9yIWmjTjaDd/VJlKvZtI/pb0zrHPpoIfeqRCQLLfQm
Ht0QhpU0JDZUsJTYpdc/yewYC6+MJ+inXXaRSKzLcoTxgxposgzfKn2YqyTX12p9XqUuE3A9ETKP
yRlcIwdMEDGUBrmfmtWbFUhjlE+GBaApIYL08Xl+Pq6BgzqJJxaNa8tGKd+0g9KDlv6cnx4wmm9D
OZSrVw4rQUyOb7/g/rE1vhiF4yxeHY/H6MIL7DJVw0GRFY2Rr8VfxattQ9xjnVuG1LHZplXVuOTt
MxAGOHE+mi3OruVeeIlIaBVrEJCXrhTY6g3lTYHnk5VnUT4O+tVgtFKfmqvimh+jKOqaZ26x3v9Y
3JvNmfS1k+ZxZHbXCMAKV3ujL/vdo4ob8r8hNrtPBcNUL91VmXO3p3s/xLa14MwISjYuVVZgu66l
f2pJWSr0Sw1bfFH2XH7fO+pkiKvdm98He/h107HEzOyXP0dxXHLzqH3sMufXWZsSVciscTSa6g8t
T7liI/u8Q6ZOAYw1aL9JYE06iiFZUVod/1Br3PhXIx3Pac3CKO7o0TfuVFbHyNzcN4a5D8e+A0Gl
uVzvgvXtUJHvYMCOaJ80B9Y/+WvzZCpV+6YDumBU6al19rE4II5bIjyAPMM4jD6OwG1eUZCXoc25
uO1nfuuPX7txrT2Qh57IyptABN4lz1HK9mceVYQK5oHhNavpzpuNUxKxiZqZdh2RZz8+Pz3RCIKV
6ThDtKBF3Y2ZKS2M/rxBQaWRRZojcfLjZDHqyKD1k91KSxzxWkBzyMLdw8W8IU4gZq38+OKUz21I
gpqsMen3vKNNTDfUKCJcGRs0TBWcAUAW7mkkQasgl24wztDDiVnf/KqPNQkH88VJsTgAeEcKlQTv
u0DRWAAkbEoRc5hkLUTDTAhMFfuHxZd3J/uGWOvYfbfkCRQLz/XMZgBgQ6VWg16cWH/vMrVLxMk+
RjFVMzTiU66tErYEpbyewtIrBJ2jbzNOqoB07k40lTyvb95GYicDMItWJTh/YnRkx+OFVyuD2fPM
Fh+dxTvS51pOJKUf4sgFdkK8oC7h1xSplcBf6T4xFdPK918JKP0S3Z7ViSNqVFfzvP205jD4FKJk
7UB7PwyO8LroSYSsWGK5RNWhmgd2ZSS04WRk0msuV/qxzx25o/q331OX7oqki5FtmHxv/vmirxDF
+Tp+ZBocaAhnlQEB5FEF12Ask343HAqBBM6/wI5fcrET5eNMoYnGf0b23ZKTzWMTnX5k6vO8jWKz
evEzBwuDXdgQZD1HMmmz5rk2Ukc9LYJcqI0RKW9ie4yUgWZM0WV+DLP+Hr3aXuBtQYSDPw0mBoWn
0PeaB2kA5PP0/ygTr/E95Vkai3454AEvEP5gM6zlW382N6RDgIs+o5dgU5DiWASOF6z76IykxkGD
xOxl+eQZJrx0Q2GpdcG6ovZcAiRP4ygzG8Vhh7aa4I23iK/b8CuuNR/XezjhgK62LX1W5jY5eZwu
/e64Wn8ix8lzZogoQxqxX56WWXasVkiw7L0zt8c6gaBqHAgB+TE1USp5fW6e8U7g9gYoQtpzRFIX
nTYxY56zcUV+LWiqtrkLsVA3SdCHPPll5dBohXvLoo0+rfL1nUzHkBROS8by4OMN350+7QaYkH6s
fpfr3tw/f/Jz8rk99rnQSu2FMqw8nVEAF/sMqE8jIw8IkS1jA1QG6oIcvkCyhO+ArN8TCPLV+3J8
lrqqsVmdJ00gemX7IxS/7XKwzDQgeMmC7m9WjEr54/lNAAvxNLPhcHitcn5r3fgj9ctRk6lOC7Wy
XpiC7JzLPuXgxegrRDfnkBzQFPKBzmsVqpJTD3Jj/uoH/vTpmOGdO78CcWgMqZAsKyopSrdCLAZu
cTIwfpW2dhh1OPKARRmgI9FfLyTC/4u4iQ6Kk8nkxYzE4K7Y082YvNfFZ5z4/fh/OONxiIVoEjxN
W7CHQLVFdQ3PSyw8/k9kHf/daSefb6+MD+GqB0h2WvEeeO6JiKxY4xZdhY1couJ12BQdqtds1Wam
z9k2pkugdMbrqN/wBrq0DorQFRPVX5nsVxN0ef5Tk1AbfEk1SRLEpIspfYDzR4uOTxmu3G56bjqc
ptATuyeWu1PrlYZgPE6Np1iH2WsNy9N9OuKyIY1kd+bFjAIKJhuZx6et0RFxnpNh1nQpB/EX/igz
CynzFvotB9+af3nUaA1xfMxWLzCJQaB7yevZFLatMTldDxOTNKkBENr3JzB+YhYlHYK8HZXHK/ED
Vots63u9ARdZJf0lxFRtk1QPnTdZRkk0p5ppl1qvy5u6Kjg0/ADvZyYj9nYJMwkGPoWzzpVVngzL
d0jusP+9cICWunTo3THi0TRI4/6//ahl9HlTFVoyReGu/dCde0mpeW4+RVLSLnLskswHYuTnBW9K
XFE9mfJ2pHRB4Fi8bNUBdm2S3rEblxUOl1iyZBSqOrtk1J5O0x+dOj4YRdU31BEe1U4s/vCo+mCq
HxOPHlszw7QTr8uyn2Neze8zXivT/olRxlCheTwcPFp4LrACgSomsRWVjXhWLLYPDow1rSpEpahO
WRTNcXrrpTxxC9q9DqvndMjV1OOymwTJ8gNemRLSGVz18N90Xf51jyudWwgdEHlJEEmlKJmpeMKT
wQa1wJJSjnmNxUEtv05Ys2zcO/3NbvTmzEzYdObp6pggC5yzLI68hFQrDOKiMMf9trq3m/L+kHIL
B+mw/WgWiWbYnx1FIOww0WmPGs4HjlCdUOJaIlRhTZAF/vFhkONYUfGHokj5+GwNZBhB9P/E0ivb
NW7WJYP0JTwg0CUwVjzCjWfwKOMbr4g2n0pB7kyJdLLeeYrydenzUq/sSdNhr9dXLbVYmylytY/m
uUWTYM6+7UB1wN1NU1HDmxBFJh7mhBlwaBfSD5W5e6Y8AiYXQcTmOWrgDZJ0t+6WaVxDdYo84WOg
qQSvrb4ES1zz6LIOI/sV6dX2rjXJRv+4vNbEwPYqXlZBLz6lbNWE0n8PWqiK9HJ/nrAsw+zaU9Rl
cbIK9c5kj7zLD/U2wM0RazWzE/glnO8oLC3MFvMd4jbULPKj6GqG3GuIWFxCO1xSgvcS+82HPBYe
k3bcMqWKXcR8EzEKG9y/z9yg7hSKyC8ARotyZ/b59FXa5ZWiXClxIQq8jmbcys7Z1y+/ukHO7OP2
6cr7OtlLkUA7h+YTg3LIF9ep597Lh5ZweAui851YqBxOxtgU2i6XzW8OdRzeJCEvRkVLm6gt4R7G
mqDWoQonJgUiP0m+s3X9SptF7yZjK03TMDANbSKUMvbrQT2BEHM3VXtfOJWjoy9TkaADOgtTk/zq
bEyb74zxK+41WcFVB1KUZOuaKroYeo7JTpX5pExYBsvRaVtBas/WTJA8ZRG0UIbie0l244w+II3U
vZ5G/fmJeh8Bl/T229Nuu4qr4TY9Mwe239m0u7HerIehPccyIBGIqCDxzTy5MdchigLQej6PJ5Km
fMKfn/LOLl9RRT8N/eTkfvdIqk1nc07KII2i3TEr4/HvdF1/Uri6W0M0h2icz4Yv6nQsVkEMJGa4
JXwq/Ef6ofNujJHz1I6ieRTsctgj5KVeaPBU+swaPrlOPbLTPRVyDL3n7h1tVFQg0CnaHBVbYwec
SUsdvfu/368AhJdx7/U2Z7VQLPUHVgRiDdIhbTXj0M86JVxYeW/pZcBAHvr2d35IwAR7DDLnRusz
hQ/A4vqiIcCrUu6P8qlP+raxuF0ORHuvHhpwzSYAPyNY5d8Ffn2OrhNE2uSSCr5IVtFzX/N3Y12v
hiJZI61yPM057EraGcwkgPdXdRAUpq8lVGPfcU2TbbVYIBTtmf67mWS7NUF9Q5WxC0I556Al3vrC
hHQIsgbE7koo6urDSek3zqrR27E0RweELPjtYrw2WcU7oyvd2VB/lBj8GzjHdGmEnNSXNmW6ilfb
qTg9Mw6y2Ex54b1XxHOX4EMf1z7oxHMwotR86c66Gg+VS9iuLPNgoDC4G+5TuLj8LW/EIJyLXOL7
gsXCuEdVN4WyaGniOMGzok8fpFsfT4FJdd8H0hknfzi7d3YfPzn9+MJutVO9H20ktHn1OSfDP3nE
trslbT5R5plaE+877lmx1qCsuxcoi06mw7bOIAXLCgdvqAxz8g9VEq6ZHEStU17YB9jTDghQwCMt
AVDt3+NRRrocD0+ryeWTGOUQ7jRSvKkz31ZEj6zncNGqYn5UJ7D9dT+qqhzWWIa78ChFhmZYt02M
rOYWUxC7+89h6+MiAFsUSuPHF/5l5enZP3WT37L1q6y/fBqh4t+NAOiq9XkrU/a+lz5f0bDzhHSq
iE8oK+iMQE0rWg03miAATn7CA+dZPMGMqw37SMO/m6vRO3AckOvfIpcCjD+AKZeEcY+sw8qsYzgn
g+8pjcHpbuH/GxgrF9C4buxHsApFttH3BsvaOc0rBoXWkiNtMETzkMk0DMPK7NMtxZ/1nsg6nsMU
nyRHRtWupGq/rHTXabj7nsLn9QdX71v9XGB3h9StOc3+Ty6Sn+HeGmsH9cRJdmxk3RttLhmwTvfv
Fkp7GKiPTcbjGB3H+Kocx5yICRvIdbFjxVwex3qwYYpPzxaCsPyzKhN0Hz28w9HMQ8yS9+o8MCZd
msCySDBbMnWEoEKh3LZ7yOQGwwMjOha7kt5MTCQ3KFLGNPZs14hf3R2WJcaTeeJhK83e3SRt1irK
7lezHo4thMwu7SPAX1O1lcFt8+b/xn3540AgtosAbzFdTaeZBtHRq4iSuHNyVIidqbzibslnkjvL
XryeRIP9o4D3VzuVMn5oK7HsMfIKEsF6pSUEQzxx99TltVkczxVtL5aHK8otua5n5qBQacq05XAt
9C/9aXxtk7wuavfd6vroYtCY2VUbpC5WsBo7mb+OwNqaDUI1fB+OmZbXHaZ9SxzIWcnS5c6/Z5ce
dkF+Cxm3HtJYM6SYF945w+QzFzFF/Xvc8DYxMogv6aO9vuNLTum5X2FZ9rScxikUFNJBzoURnwml
X6kujHl6webZAGjlTq28bLbuK+PRrV0GKuRYHDoIZcxh/0LMM8BD7DIonZ6zKQNwaN9q5lCrZTzS
mQ9xiZ7GxWdKHIF9ng05UUlXn24rlO7aXvVLk62dIRvY4vvjo77+yPQOaFDs8KRtWIOIPQzB1b5b
OSTtEnbXHTGJHTfmoc+m1eOPrEjlcqqfB18K5a2LuFrSBxr9p1nWb2AjNYP+l+axh46f9e1a6Y+Z
PawBWzHjph4vqaipvX3b+sLsFnYpY0MkAXCkUwTyVvo+AXKGObDoVDa4tjO6DqKd4BIIStDmL0F1
mg0q3s07Dpijz0jIHyUmgDUK58SulKJNWerjdLGu4epcfhHK5VIL0tyKc+PEasIgxCWLXq2v1JcI
Y5Q7wP5Gg9pH7rkNJlCqsBNaBQR/ACQ+gWUby4EO7OcmALZZPV0O8Tv8Ey+RiT4C18qDXiVi2JOi
8FuQTtwANSsURSnzaWePd1FPiDrDQTYqnNUxLMDACplUnTp/G6P00Bg3a0MCOp0xjVvOYWuV2btp
wxoS2VDPT7exkhCIv1W8YuOa8Zu1e74TPDgWrlUIEwRXtRZ9jwNmD2XozIV0iJodzcV2BSf6H1qR
c2zHsxhrjXncdG50jpFbUcWNyanEB6pCtQ4IpG+4kBfi8nEv4zbTM/sSnCXYRBABc7rF/TE6RW/g
h/X9SdSUh0+3gk7esSD1Cpcnfhek8JZSTFViFrh+RIkHVPl9oY8FGDz2DEMB0HFNrvQ30pAYqjB5
ztNlgVLW29YwY9kRn3AeC4VG81JvjPGbxxZ/a3UsFhht9+k1SzxEYCyC2D1ykThyTguIpSkiGaRR
iPS76eWeuW2rjmo13RaxzOGaSuYrytUiQ9buTsLz84JL5Z/yA6emEWb2qiS9X41UX0DJ9UWm1Vgr
MKxflVVxGpAvDILj201F0jW2IstgQXdfqmn42iYv7MZnHodthyvN4mmF7QYziZdigcLM39vnCmnz
3i6ZwB3ChATbHgq5EbotqJ/DcA82gpuxP5z6uyfIw1EecU4Edj3+CtBZlTal59ZLP6crC1xbMSwF
glvOpbjsqruevw95f/7ppdlmfyJk94jUadSeQptdS098t8sOHTkEPHAUsDh0BlL2q76JUIEU2PHi
qjd2B+iui1OQVKtJ9uUZONHwnxsspF2Bx7W9hOJuE4rwKjsR/7t+q4uD3r8KMpBky7AlbhXQI4fy
xTYEsZ2xsCe//n53cQvPlR1vUzjzUssVviGnEjFdSa1rCMXb+RB5ISzgpJyplr6VgRiWGuLfGUCn
IoMaZNpFufTOJmfWyDnsVVHNma0Uhi1OJCKluO81KHJz3gZFc+kiF1xOKLXMsuFlWx/rE1VopwYc
f8EiNitXsUbsAumv7XL1fPGZdz8m2manH1AfcmSXK5kAhY/eX7fXAic/AMmWfr8TURY0GMGJWGWW
+MH93J9VoVdvrv149ZxDjS/TXAKkR1c0J0pjNv/bVfpAPdVY4GIHa5gjAnvxIjbUoIg0Apxn/seP
NcUuQFO4LnXgK0yygWC4coZvTbClgGkCin6fI6QIQzB/Nz22Vn1t1qE8QL+NnM0mikt8w27RSQe4
jRWC8dGCADcrO4BKF/gEC+hshP/Vp4+kanWBahn+4yR82DMzPi+LWqqXmtZjq5C/hS+/YsrYu0H/
VwSO20YqYzU8/LWa9GQwT8I3ch1AvDKXYjiYLJy1cwgiucKlTNBtBtmASveQe73lqFdqSuvVfkhU
Bva7Od4GA3rT6fWcHMixitXGIJngVSDXcpQAB5xfgjikKpzeVEunz4EddOHLj0Hq0RmPkVAE/LYq
90MWvsAr0BBLLuAVTtJQFKUHYuOUqQyUlC1/Ghn3F6X+lnjyJYx+jl2t9CJzNiiqIJiCdDX9KjA2
WQXGmA7hzx0Xoru9kTU6A7xhlwglZuhYBoLA4ZtLRoqT4gtaTYHgAUcmieyMlLf+DsI99kdzPspr
xG5dwB0pXCcM8MFKdtmTTowCB2lNQYsTf2HVOijiJsFYwLn+bxdTrrB6TEXgzcHOv5yVPM1abkXK
XFQkRSxQ/FWESDbLdSxG8r1W44uOvzcju9cDHis0VJy77X321YX5cx+nJqAo+SpVR71Fz87ytais
J3kpYqfcVKxURgQvc0ePRAgEI50p3Wu/FhHqgrVsqDVGP73v4h/jDOvLK7JvSfl2CUzPCVvr4PWt
9/+W4hGpKg3N9JX/LwdqIoMKxjHUkXxL1EpW34tJj7rwXn1KRA3O+CGDZ8KlRxBpmQQJsZTslOCs
QYxA3QekQ/2nZ0sAQ+LkxIENnY0j4ZodR3boYSosCUI/8123cBKyU0Zzmjq7Z6oEYk/BH+MFZxWw
pCPjZF1h9r4NiNjjx2/5v1EI/O+0dnmJokFJJaF60GocY/VrlZrovamFweGJs7vwfGKS85SrlLo5
bhZ3vYbT5Qsbvn2X/Y1475hwfBSqUe66p35DgdfdKyJO8OvjM+QF1lMT4bWagtIqMRMjh9DM6q8c
sjprpBK431ppdoFuCAoeaHEVvqneruG4L7ZHH0Xmvgmtxaw7I7qzEx1Z+AZCbLSztnJgGTPkV8NU
dMGT7atQklzLs3cv7GBGdT9pNlXm2omWxRI169AlM6CFsN/IRcdX32p8r/aqCrnCOlNE6Hj/ZFZR
dErTqFXEQ+atmFRfXKxXzT5MPnQ6PfSG9mGTx49ORgUoRbANssvUmm2nqOLj067qaLc0JPAnmrMT
ItU39UOoD5NaFFz+72qH8ddyQBfdQAm4fy76CeVEOspSpr1NbROZ64xp3SXNLCPUS/6LMz74OX/q
lAMYyTGjAyN0AGMJ/5sQIi2rJn8HVMpIxWMAAULJaa4LcbqxQDt4h694glUnTyA9qv6XYcjZi+Cp
uT9FjN1AQ9aszWHT3KoKzQ8+Khd8H+JsV0O6yavIh49+KkqWYagYBU3LcLB8OPpmww/K7GPZ0BD2
xqOWkrCm/tol1so7y0DFZLVceQUrUr0UxGIh0H3nmspYMG0Xs8AZ055Rvqz/aWRvnFPzrvMe9/tJ
hDDjYy6AINaC4OFjo6XKYUnZvbhJo3Jopgzn2oZUChFdCW8vYLB37PeAnsDPvwoN6ZEFzyZMD3MK
fZv/jSOSDW3FOtdhtWqzFUWiti9e2AOkIpdCYWYlb2PN3hk2GJw1KbLJaodRCEDjKOZ7SGkCQ5zc
yWt33He0Kh6cjigaRdzvr93RyVaIUTfh11PrU82aAHoLIeZSY2tlU8xCNB/0/nxjD+7tTmXNZtNR
uiGcqpBWGstr3LMcwUSyfmkor025l4qnwWQz8B/2h0Wj/fLQ8OxEb8l5qgY9S8PMPKaXelCVAxWL
yk3T/6NnFjkpQhro+2pGcASdGyDoEQ8tbXykWiTm0OdTZNUm8XirzujCieqGjKOyg4lZfOT0+bB5
yPZ7X7QSBNaILL7XHxoTShBw3/PexalAkpQquLz0kTmHsfNkOO5j/w6VhoXCDpGgwxuiBKXJJWP9
ZnieAGV3Laiyt+1D8N96PPkG2S0FAnSRLN238G6r0s8qLt4ky3K3xGaRx2P0Pco7TTZmY3g9Q7nb
9e/OpchTAMyctspImvKgcCjDd6JPUjiiLDm9KfOWbXt9qOLKJlr088mqhIRU15y6D3AEn/M04Uzq
g1g12NHgp5q581QnqGWPjaiCr7CZ3lU8bn30ghM+SsJ3nkccb2DJLEG2V6fasV26GAJ4gYri1One
F0hTjyTN+U2jyO3iMsyGl7l8q4QE53/PQ+ddL5C/DdylgmJ9+xaIUxMOJ9xCnZHtZ+38QPhQPM29
QUB9xzlQlFXnw7/0MdhBxU85Jls6PAUFnkpkF76YeXAl0qsnpCWVFZT3zTOYY0OH92QGP2tl9ZwB
0+AWVlvPrHceWwGI4IaPRTjRHq1yWD/ABtaBI+8R99Wwr0X8mNNRyaM0lhH3crf07rYSsWOi64LL
PktLhlxHbopZ6iIfcpfIETOSPwjY7+g26KyAjMMQha5Dit86SI3x7Msy2D6gFAm2Skp52QGP8c2A
Ba4EyM1WTFiOSLWXVk9jbzoJZ95lHr4ggGIchcVnQYZvaj3je8LjcO2LoWJIou0u/xG2CgrrjTDQ
lWH9MBCJ+/zlqHoXieDElo4HsI7t2aPYJx2aoTCyHBz8jo8ySRRwy4Exu5zn0rS0g+Uhf9nUDLOX
7vHX398l+dNB4d9raPtWzAp9L9XGEXaRMFZohbUvmI8ulj+JVzFYfnD0bi9AyIsvr8Tfr0RxoCia
RMquXIlOXNOf5EOBTKvRsROkZB6NGyw1lmxaAq+5FjbP2gN7T18NAIBX7vmm9bLqn3hE+RzljxfV
2zQZyE0dSopTKveIO+tKq8AdMLYBj8lhhuwfhtPlJN737DmA5tZMst7mUYMgT2RhBdB8Zw61IuoD
TYR+qBAgd2vWr3wHzaH73TY9rtJJz52o2ZdUvZ5q5TilRY8ocBmZE1Vqrr+lj6CQPtGNae/iUWaH
UULxN9LK97AtOExE01Ku7rIiKKi+shgYL4sbMr0BR2/bd3qQl+eZB7NIj5rRM2yvXuQVfiMFWVjK
5tP+lEPPmvq0xJykypEyYyYCq+z+zrDaKgZmZg1Dwh+XijEuORAeW4cdzWmLu2fir5eMSg0XU1QW
tDlhCSRTmwkowHGqPiv8klTRjjTKrRVgXCWhaD3Tb0upauQCY0VRMXknC8Q6MR/wZmZzRpu3/iPp
3eiy0ZrulF091FjH/p7rYJ6ccGxhvOgYpObdXtRwnpSTCUMVxKTKP7ewz4HXPMhae1h2DKieXdQ7
STT/wsphFBJYvoo+XzoowIZxQg4LBUbO5Ys2ODjrKNAGVgHA+iay+4OvBKrhKb/L1uqDTbTF4Ccs
rYQ1rk62VD9NgkG4vp91CJ5drVB4LNEkVWVy7aULtOCURhfPxBcO+lps4ih3kXF3FV2eCu/fU21D
Q0Mn67KDBa+JeYaELEMDOpqrSI0HOlSDfghABGtruTjfUpFz8M0iIL9UUJdht4470sMsKZ4YSlfE
7vX8JG5wQDX4fjU2hIZFdJOw46BWxDagJZkfUAyIesXBG8cfjyLEJH9pkwFTvk7fggtM+t+ixkRs
EOtuEhNyDAEg7ZXOCkgN/UN3jcm4UwfiviW7Qc8MYOLqOYBFXWUkNHFLfYFNZJVg71Ad6VIgQCHF
1P+QGSrlDNJ4L3ZKCMUReg8y5ek9Nzks9FURRb6y27wla5cAvRMSw+jZe5M1ZUdW8n5RP6TmAJYc
PtaoNQiS3Vuys3J1rB9Ttgy6NFijQ0I1+5Fi0an6/htRVWr0CbuuEgO1+uMLDgxWCB5v1kWvt+Mf
oWO4SPP7DpL/94Or5lt/9jH1NSB8OmSTLAjbIeyjBdDdcUBq3nM6bHoOtcDSgoj4BMBKpDbEnPt9
TrQyJikQ7FWIrgB8PlB+YfToeB7cCBjwXi53GptBJCFdb3Xhc2ZET63fS7qgtvUVlj7hx0aJayQ7
FDvqFu11TH+o5UyG9JGFsVV6y0d8eHvphLR7HytS32bYuN9OMo2mOT25gCiF8sek0M/MknIlTScH
jwo8HTKmG0hwJR2G3Pa5iJ7pPGI5bRpoj3GAKC1oP9RfIRB5GqlA9U4Q2vHV6/je/0WDVuVRZ6/x
WwXr9wj34ebU5yLsJyPcg5ZhYfuWfNfg7EHsdMDIQTIs5bdaqPeXzZnRxcPzwWbN2PXnERmAjjlL
rK+2bdstwCecx/M9DKNqpjvRe4OsQibnaPB5D6j24IKSyykYE2VLNmdNR9t968Yhz3Y1RDPhLwvg
/a2d2cJhJrVLZDBYqBAcJQqHWFB1pQmfi38A9UTkidxYw9gguuaLucKfR0uZZEVsmmEXhNuM9HkX
OHqJAJ92GRvcaU7zU9slJ7kiJz1Lh8adicC0cSHWCf/H+e3/3oDn5NZ/cuTKSKHgTd4DpVNC8Y8w
dReu5co6JFdYYfCipBzLWksPKyXFCLHMfPSVw50RfE+EUpEPAfWS8EocmYaiT2lGbTGtueQD62rY
OevvUcGrTVyCBX8bY9a0MhZteveHaDwXRN+Y+7G5KnhBBPVNFuLPqLDmf7Esn1qTSbA7UhO3MUls
+OUvB8pWhVXaZq0iqY48wdRuGv5m6lsoLwv/3Uq718Amho3dUVcIgJSFLG6uPsATODRRW69Csvsb
L+VdvTdG/LuuZKThuVmLj7wcbOu8zWIhm7mASsy2T8S63AFS4YR2KoyIvx0OvA/qsvFypXupnNBq
topbUV+Nc+ys3uBpI77X/M4sJ2Ryq4f4w9SRGCJqnvC1idTs2cc/W/JkLFiB+APgR4smwnVOWh7h
6qG4qUCsvTuQkR7cQndC7d6UUta3Qbw2Tdc2Ui0U21k179JU6N2ZS0UeLwVuT/GmQi+cco1DaWUz
hYTq2BQLeLZvRDeanvFhkQsUMia8HxBNtzSA6o0GSJhRmALBXxQqsuEGoyYLIzJoQ/EMgIqz22xP
0imq+sgCYO3Erza8ZJ2iDOrkOJS6IWub2+uEeyGFol21zKWqljGh8w0kYz/aCrksORKFyq4GdknP
ce53+u8KI48brd8MYdsM9kgypJ9vg+NRZUgC6zVqEDIAKqtCk216+SfEaXowmwPmpbzWYS4nfVDW
mNmSYokAD5pb9f9LWZpR4vfvuRvymYlu0Aqky58+lblAlrMHrKnhxE1pJHZmxEE2Aqfr45Zxpf2H
962JrWcr0aop/XDI+MkhGlcRG65kgv6nxoIP6kUvBAVdbjzKHvQsTBH8Xyv2Pi9WLW8UpJ6btT3I
xifbRFpgfauD/fPzvetcjD8lSaDG5JjY9BaqDiv9yXgl/TpLSbCCSkfB3/ll6MsmAusa+oHpbV/L
Sb9SFTzpX9cD4/3JeyJRxlOgPWJDebZEFOtlTFuYAkEKOpebmI37+uBDDylj6ZY6GVQ5hOUGMYAY
wwZbIDDe0Iou2WTJRRIpfRMgvMOTwipYRPeolHfR++n2BJDCuybhLzsOMkrckcu/XRW4K0+x1kk9
zZATULAyJyFy4N60+O7dUFZr4BICMEvJJ43ZxGGOBToYDykdCqTq7XrGmRHVjZgZBlh3G7Q2ExT2
vhb2qazebmP3OetDeoa4nHnEl21cIqIP8jrUMd3dz2BQkTqFW7ckUCmVTLhEsnZ5EsfJAjDT4KQZ
T1xhKGgiH9BN6Zogguw0jD99RWmpF2Va7+drp+U+1k+Qz+VlwikPzNRdGD1s8wBAxHRnFjiSnn5f
AkIlsGUD4vnrB2xQyO7KUIbDM8lUEl55q+zMSWS0s5wFdV+Qke0A1renexCDDUqPCux2Ae1vNngK
bzLIK0n+5F2sMNZNFOI7fH8sRFTkHG+e9XrmrOPtSBndxqxvyswbMPQDPcIqOkSwWGxsFOuLI4ng
+Xhjd2pN7ddKWLm0fTtbMQ8RoWzbyAf1Kak8G3r5+P2Vb4E36BJ3o4vuIdqteiewZTw1HQhAgMvk
X4VY2YhLvwmM5HjJHyPsPqrlHQC92xqKO8nUOZRewlSLLU13uIsozYszyzrrT5QA7YBKj13Vp6cr
1mmZtvUGsWEJjGlMu01zvTMdM9/HNV4vp+d5Uyjnuqtzuyht/dB7U8OlmwsCfC2sBZF+AM5q8Z6M
GolBX7YbMgrCTriZOh0DJaPQ7r4fCluZWZpIZcjEjqF4le5avJ60dXLszzdLsnK9G3NmkuK4OiRM
iph3IoIRYX99RdgCFy3MdDWDOAT6Vg+EjEL2S5Id5ZAzgNwb9AxMCGKSukl+ywxLrVif7xznTS0Y
CKIZFQPaYTnqLQR0O5TzyA+9FX/9CKaooXxTa4m9J7tDZeOFYbGq8zZ5p6xs2piRsi/2R+eTtJB+
gdeRDqo0NSSPozRh2f2R+J0ov9DtFOgz+TduVZ3EPm4kio1PpEoCcvFH8guSub+3rXZTnksu4sud
pNGd4uj5hRQdiWrZz9xHsYyv+ntEiE1lNXtPNlDb+omZVrmzVF3mz846SCTSImQR8zZET8uaQRfB
EWDitWn+7jLDNHtzXxT2aiJrVU0xwuXRLokWJlEFzCk+o/O2raoYW+2YuSenCCsNWg2ybkN7ksSW
wQLwGea8ge8r1z3usp+L7uwgKCI4wjeFxXIqGxsM2tAbMGcYlYOkm4/I3KFvVH9UCOtvY950gs0w
YNLuRurqsUEvY6Smad8Z6MJiVAo49IfacQHyaq1xPFx31aadGcnXwq+DfN07QjiDrlNfVhWmK/Fm
ZCWvvEtTidjbPzu1CIgke/lYg8NScjM/kyuu57DNXAogZ1hYTLeUu8GgvYujhtksDruk2kFrA/Oh
Wz1CU6BRuiQGCvQiJpi92FapdCq6uBcVnXiWI8jHvaKRQBFqFjvpQCSS/ItA92VgvcQbYmI9tzsm
nJv1eT1HEJTeHfS06VLjkDgPslKfCOGKIXCXzcW/UAa8eAEuzQg0OSKMVVV6GGGCUXHSjEDIu1Qn
xJ30V/ExpMrP5iqXhfE+IOQ44JTrxnUl77ZqF/cjUyQ4cW0N9lqGCFS4S2S4dkyxcLjnIuZuJtTR
W5bYc54VLlyJJQCvAd4volefRGlxQKGl3IP6HwJyOZOSmaJoA8NelWnjMnVDDTnAQJEKKa/sB0pP
vEbT8wL20hKs+11g9KgmdHoFwVPUPGGD5Csh8K39YQ7+SwtqRYPnOskXW/Jd6DNS2y7RxwhelveY
XzkEtOJs+XDcrF7vNi7TgH9Zvv6m3OyBPRr4D7op1V9zyv34ns+PG6q6aBEa6NgaaXYsORmYaq9U
CFaIgmUmIgRwv6pZrIJlfEQ62yDft0vfmwbwp7q92npYObuFscLgznqhYCgj3+zpOuJpO/l4oCF2
sNUfwm+6aa087AIXmFEXibuMqQDmzqBGj/LF/ZHfA3FmSoD7EdC2eop6MNraNAaVHbvN/WmVPCqC
nq1Q5dkkW+RZYCEMdTl2JC26YNsCe2uIObtUxl8wPaByXR8GlMXaYfoI8rf94cj1mi4146QaIsvN
LtS0Xophc/UL24B0dHsvgmqROUpQiE7ILQFFzxS2s9ZHkB/wnd02vZas8LAIaCo2QtaUsO7DoTct
7CwI7pUq7ID2A9z1jEOtqrWHxqe2w1gZPoc6kUKLBsKGoaagvDlrY0iCPbak9nB2C4zOQ4/EEdEC
1Q30q5e31Tpty20as0Ao0sWHPH58qKZ+XeqmvI7ih95p/SeLszZfY/1vm7w/Ghy1CjiGawj4RDy0
/YJDwgknuhDVZ3Di/K1DVxudzu1jJ1O+TxBio+vn22fLHbFniuBDEpEpk3qyKCTjVg2ImgJJcMxY
0OGKm99zvMSy2fuT+khVRht5InLRHMmcozH9p60j/W+w6bHT2rq1W7bGfd85lX2vXDurF7DXtJ70
qhuGO+oeT/QrttcA293Q7GwNpEpZqrVbwxUdw3wv2USKwVI0t9ewYx53KDkLactHTLzibmxB8JHg
XuG3Nr2jy7GA8CktuAYE8QiyCMkb2e61ARHNGegfjEnKbkaIbexn+1qbI/R884O/p64u396BlxjP
k+5PZprEx1SHLcYhrs7KpbYmnk1YXsoijcIfjMeX9HhjM7/zgR3clVvcbkHqywfqxrElU554IMuN
dZkYHeJ03ZOoIvBXs87VTBPIQsEtmX1sP0Egs6vZyEe4GMnL6F7lVXTO3rQkbOam1KiSwQvQ+Dww
ON0abTici6j+fA9xleVsfSFwK960AVuehtbuRrnDmQSorSCQx4sfQqZXWq5aYc4LD8XIDPsmehws
hiIYoJJaMyTQlb4I5GSgeMZKR1/xIYdzZaKmuhPYp84PGep4+s3zQp18M01Y/+F6fY8kgma5WBxO
vzYIA043WafEMShXtA0aWc0jz200xPFyGf90k3+aZGIMDSthESPtANUQnVgcUEXXYHoMz2ADAZbG
UhNTceZxuPeYGuWTX7d/sS59Hdq2dLedCGyCY4pu1LXiSxxBnrdlA9leOt2gREWxHdB+VsjhiYRu
FfPPxmUVSaSTDE5F4oDIbs0kb/PFjVtIz+Na3aA7LvmOaNUJsw0Dv/VDoaXVJuK1cj8cMXDqgy9k
NPVOv+sqR+6fmk9UrA7sutN60fncflRTFY/EewMjq4nOz0yNBYv8YqL2ne2XdmbgXWajENSYzzgh
nvOecP5+30eRo667cQQDgj7m4+r5oZ6ZyvbDNuSMJiV+MDAD5E8KwkN9YwxOfQxZQ+lXOKe0lItI
h+sMfdWPfgnzXSRdHU2OIEVetcbFah7m80tpH7GixdUej3mTtWH9fc9hPtMXbyjQQeTurBI3oy88
t6bEVOq5QhhuIcsxzXvxkmI83lr+DqV196NX+mUgaamNhmS80P9Yug8siuzy6WnS0TQT/UxUJ/pK
lpZcqKHGj1B7/nhkmP8I5akusc0o+wQelSUp2v8dNOfTJ83jxoj7WLJ2JYRHaWiS86I7Suu6Xg4D
/z/gJB7blF+l1F71zPhA+2jJ3f/gkSgKnrOHQ/tIEanjqKXsUMpxMEOSJ/nBJlrVC7yALGLMNkuN
ndJLmH9BO19SqlYrHYcCH1l6jErzaK2vU9HIvRI/f4GkTFEEd74qqfixI6GLyAI/DiZ8m3kzvEB5
5jkpbZVvj9rWS18wX78cuWu72I/kTMq/L4yrTO5YGOtcFEtGkgcDznCdY0ky107zlIIPeF2QrN1A
77X50j7M5Oc1ZgG36UFKrKZYBbWp9sxdsb8H6DYETzwb4q0Wbe1COeeP6Sb5rP4Oc/VshCMH8y9J
/bSTwFNvXx1rAJJMX5Cx21Zcjxzz/mqlB9PmIWJAmWnflyYu6hNRpzDUyvdVrrite5vPSLdrYlsp
N+bbAskLTy3ArC4Opam16SWy5VTmPZD7FOIRGC7Y1ruvlClaeAoCRnao55DkiiPvOcX5+JkJyLiU
VlN/TBcctyy8DTR3zvzfXBWlo937+q7D74rZ5i53ax+MKo/Ved7Joj8EmDbVwjr/i/4+bOkN2p/U
19ZS/VmVLAmVeHNuV400rcpMGN7/uron7czjfO3L10r+oAaLh9Ktz3V6Y/GhNN1XBsGAP+6rurLa
hJZ12uIjBA8aeWWdLY5xxowUNwtpHzd1mnzo6O7H1H4mJBd4AXfJmSXz5OWN1+LTsq7FNKhu0Fus
OOQ9oay9IPabKWzKB046HFs/QngKg9oszjxa9NOh/48PA3Dfq0tjyEa1VxTnk7fCr+HNMrYBsCgs
ke9gIsZ4VpeM0D87BMgt3myhq7trhhtJLwZJu5VXD1rImjoS6ZwttPm2m91g3Se6N46IIYwuUTgd
nvsYHscEEwqPLY46B8lqeqV3bxVE9afugE6ezHwfxO80cNRqnDjHxUBNqbflQGkkhZwSVhBWnlH9
X+X3A/WmgW0MN307qRerqNLflDR67/pUkdBBq52bw3rNYs6EhOXb+rYUQj2k/vJy8UlT2kO0e6SO
/m2EAggYGOirpMtVPw+5FfILTOy5F5mkSps4dqhh4Ax/0jPODiSDQGfdcFMmUZp9dESEVxcY5Et6
iI0xlaWQck6dMkbo/P5zrQu/3ko9lUaBC/rihm5GY0oMKcijc6xXjpsv3geyLkRMvPbJR05IJtzx
e1864IWqZZSETQX9EoUtLedDAqu92uqjo5rRmPLrA20jXDcimnAylIyGlxyw1sMEoBYIzm/G7b5E
Ekwh4xATA1ZP0qwhjabuAjIcttYJmVsZ2w2JryAgsDIRAJRIUfeOFCTRj/ba+AWrfSi6Q0JyXphy
uZDyO0S93MPU8PPiAC8YcID9hOoySkjUcVEIQcsaUrMzp4EJNeIrQSfaiVEQO6NP4PE4OCzAwDj9
Znd+kFgRChF2GG2fFJwq8IPFJknlFsEjfL5GNfPR5x9T1wwKLAbA8AxaMbrV9huNkZEuqAZph11O
Pw2hvPjvEYAu9Ijb2H4EI1Tq84T/pbuI7gQjx4iMcSiguuEsxPRZCFf6+NA/JrSrZNqFLkCpQuiP
NuQEayPgfbMwCM1eH0vw//D3hFqomSvI79XO245NWIfZU3mbxJnoLFntNMQzKYmMt2NvHnf/4FX7
fEkrLtACUQsrxTeVeMT3pnOaMF/i/cqtwi/IEQjXxTyIbzPw6CGQpT7zbFO01WLuDghQ1gy/RG4x
+GM84dBvxSFAfGMfXQtPlh1COgowiM9+yyrY2zCORopIxI+l+Lq0Y2L9gTxliDR9xBAQl8zs+WQF
mNtUkV2sI+nI5c0I5E8FrcttoAXTQnh36JRj/+t/z6trIGWPCgZStA9SrgVjOyypgVlpGtzHhp6E
soO9/6A5Dq/bxVRJ9ul9eeSAPPoepFduLJB3OaG574PYCP7Hk9Wwvt9DMoyuVJJ/ZJK9OzYPGvW4
0O5RkzSFT6g+kX9LuAm5UPJxMfhh0BpJxrNJ8tIJWIf99Zq9FGct3pS0JQP5TOVMSXFJQrUFLySS
l8ifXY9bAAGvdOJdrobqxxtSxX8j+PuWrGXtUsqu0XMaSNeDXLX3FRhSPvC3TM02co3qXTz8DGWh
5cKt+dWdOaibDcWD7Nbj03vZcRsmZv6Q9gmrZ86ZJxrUjDAu16oHhlR+AUj1YGFyruVbqOSqj+BR
9wKHDWY2DvsDemoJaHqFAXoLBEH7om2bu0/sortcQlM5/5khVzUqYT5CinkudiraZhReNQxwDYfM
744489JpbHd9fc+AmFZgbXeTJRzxw4Lvn1QCjcbtckL3VhT746GcUfOAGVQMDu5eoHrlXpF665BR
ZqJJqsLMu52onxbE2K23QDnP1oSzKpozkmaCLHYV+CyYoBtBVYc18ItAzuzHz5HM487ti9BBWw2s
rgOGgVicFPUjM9R/UIrD4sDxSXUIc9uD8U2u5ROFyqu7myddmrbTeaIz1sRTUIxf/TncFCK5oe0T
5nDGQBRWZgfXWrEAN+t7vUnRtiMztpIFTsIeOz0E4gtN5vIcypKYjjEVlfe6o1XVqtkQ11GLCaZf
SegWBmXgwgajHB6ypUOPRJlEf4jic9518N3Ojomp0hDzaihD1NKP3uncJVrgOUNymK0kur1H9t4u
F2TMtti16j/c+pTGWU/g9rqXHX0ZQYCbDRS7qijQa8YrFc7QVjHXwb1f+XbW6yYPcEdPj3ywQnpo
7dh3mFIDNOo2Bi+X97bAJ+eTVnb1xXuxQOnGVfEftvm88D61qzbMXTIJVRDcLMvHRKvFQlzt7PMz
NUif1mkIDcU+0fZSZEywL1IwB/nIPz/myCDAP7fpillfcdAXJJsVW1t5KkS2VGnf9LtsYUdXBjI4
5/r+1FUPAsJ8jAb5dKT7WWn/bT8cjGMCG+sdRwYGcSQpOvCBkY9UnC5HiCuXl1CJIYt50NF+imWj
5LUufDw+Nz3+A7ntOE0aW7a6DbQnaxsLegQDSHUN4pXt4bMHq6gr5/WGPfpatmWZCTVTTczq6Wh8
O/ZFs1rcN/GxZmKT0L1hkUtwfINbIO4ji8ODCHAP8sDEUxa9ulUC6DZ4MSXt9MypEAH12KvHPVR7
0btOppQlPcxg9SlufnOUE1M7gcaTakmld1PHSHgvr0fI0VyUVsm/iSXUma2BTYXCuOxC+yR7eAyR
6ZQQDYACkBpHQ/hAq0Tr/db0jYxlPOxVuHQezE/tKbP5b1DcmZLeVQoV1v0TWdBLhbjZZChhNpzp
O0LtXkEjIed23/ooOTBObbEquyGWW8/O7VvI5uP8CEbGvRwarBQMgw/OQXYtl6jLYh7QS5Jja9PN
OvekguoZQi/1RAFSyArHs4bXmH1QqcFX0zz77tSOyHk6JRNYOD3xgHvsRe6PhmPUIeDQ49u62ReE
4KjyI03k9c+2Ma5GDjzKl2t5mGR3A5/aF0J4chWfiIWkNA9HnP4sxg4hQottGwJ9L83LSkYyhJTd
fqkkAdddjLukPF2001h2lTqRDWrD3/pqpVH49SFJcDiGZT/B2YJzxVftUaQM2Y9QWGwMKtoshm4O
eqqCK4cjzya3Pp/n66Jae5sBbHVYGNXCK0t9Fn5LxJCCl9iwxFsuhLzsMHmoDEF0Q/tg0DBxzrWF
PIB5ntyt8wgGtePVotOgTw7DHoU3iRLLKoB5g+UiyhyAad5wDJl3a8w+9eTnn5hugpiShZg8LtFy
b8volKw6bHDUEq9YrytTTreyVkGGARt04EDlaNoyPLDpZ5Nijbi1l5TVdzgWxg+tnZDN+uUZfg7G
4ycHN1iINejVQs3RLf7YCh0o08D1ekSTZWBrBEhdCd6tw/1cseZHgdQt7lgZIgSqFREjZOJpoF6q
hqWPqlk/vlIrfee9+I+TT9gdB/wvCMyBPy68mq8t2SA9Exv4D34UZYERyo1WRhJjFyroyaPukiSh
3vwC7RZOYGOH4px0gpnb/OGe82QuymKQ6TGQeVMe515vlSwMlUHXH2KLbpBxil1lSB38WeuMU+AD
g3Fc8OmldRQRf+fRuTi/YqvWoWfu3tXrOWtkoTQYZZlngugtjaqA2mf4WZ0J+3iKdlHW5lrIN1xm
+xCqpilq7Xbuudfl+5Zs1nW52FB17ntq1korLKrV2fi/TqNE5S5FO11cpkGTRDSpHMjM053aOQ8E
YcyLsT6am/Qcy0N9C4CMcB/40XJRo8bJDKJOSvd176Fh5q25TANtumyDtN4zsc+uWhqqZBEueX1V
Jn4l6cuH65kG+D80tKpP1ht1MfujRq0AMSfoyAfZrDLidP+Nd4FjG7rqqsfX0gE9r1wutNk+pybX
FPGkeNq1aTPT7cpbaJdt3u2CVkxZc5xTV4qNn/XJODTis4XCVpiBKkB381BvQddfv9VAxz1zoiCe
CkqzeV5LtPkBrV81nt7ADqeFbbAmbK7FjUQyH6QYaisEvnF1CZ3EnUViDhT+FjEMUEB6iFyj0qUv
OrGTHIZRayEZIc2dTTmevYo2FvTKLjywMYDt7pb3sGY5Rm0WiE+GZZ3+g2h32Vvbp+ILiC/BWI1j
GIxX6sNfcy2I+m+L5155+7zRHGKYAgt8XlskQKEwkYps1hBTWdaf4JeNGl4bRtuzju1GAdzk65v1
kyTLzybaUBR7zG0h/iiFWd/GBcKJHTCW862eG9qgSwZ+q8GgJOhIUJZG8VAoWWt7DFKfFYY79VCB
RqIqivxjzrZrDdaFx51DpWQ2xxIw86dYL3zOTw0g1A2XCa4n0xLFYRBqhnuFN4ZX/aDXSn32LA/G
smFjA1AoxRgeuEASNS9Wk0tB0nV01YyrwHg5zPmVuHXLvmbVOlzyr7OvO6yBRxReQaTNVzp1cyTh
vlkUaLPVurtB/pns4MV0YXfJGbjG6ZokfWK6dwr5XoRTdChtSsm/GCZr2MSgkpNyEEc2vsGSYIBy
y0PQ3u49AqLtFmBPxXO6gPHpsol3YoRCsneALQQl2HgZpKU2raw66JLjO6IpAA96GGcAdQ2OD5hR
QqQYHfXkdm/BRY29gYyOwBzk1fzDp23Cgp+PwETdcUCmAugU8Zjfr7TuY0Vh6b5MPbgPVVVNfMbt
FAMYKm5GDgLnlnzHZb8aIea8nT1bNdHflf3UHERRjwYIGL6V+lbhev0uR8c+wVPrAMpFEteLR/gd
PTL7obTTNxSXGQQqjSzlRwR5loRpfQx/h1WIr9+uMU2wArpAhf9HU6mbEz/CcyTCUncqAlScE8Tx
w6s0Ol3XCMbuEIY0fyMArCq0bI7wWs7vRzsB5dzpGBNTCtJmR7BzlwXkuvzlg4zaXVu9vqPGoBE3
E1uLCrO5HciwaDP1LlcDzK1Ibu5muHd3YsJlXgYGX9wIvxv4/aQL419Ra0BHdQHv6AkUDBV4/LF9
Aj3oBm2PxHxzgwswluVy0ndc7RLqGqUutPiYKf9WSEkEGWDptutw25eT5IkTnhNgELWJHtx+TvKh
33IESMwggPgPh5P/S1F3Qmd7Zhxe6fLvw+GDCChB9RoznKsDzUgFliT8xUR81GnVDaCCnz6EWAwT
cFHpE89pwcpSLiVQ/FBREJBKC4wC+duf1vGU4EW7W+cNMAh++S/fTBvTrPpSy4TCoDzp0OS7IB7R
9f+PU9F5pXWtoPJpcW2kCZGwYJck4aNSaFWtarjpmiQL+rZyCnG+trmM5oCBgLvt1PeIU6OYu9cd
y114EgYwuWI2lG6onRgEWfKbeF9etn3xFxcubQoLfO+fXwzFFRMBo+bBES4PD4bwFGoSBlzIowIh
WZxweLnd1xlcOccNDoYgcu5hXsGeQWmFoN5tEigw1khG8JdQTh3W/NqD4ew2/nst+t2MTrgjt0uj
sR4Bf8elLArKERy9PSz3tbGgYDWgXp7bRN3CiVTthwPWBpWxyr5KyErkcIH6akxTVj5BMU8B5GKs
E/UZeoviAkRmtN29Zeki/JNrl1843h1OUAzhuK1yCjXbDzSuE8MdDut0TFvGshp6F1Nv2dKopOKh
uXINRlChnbSOxc0Sja1N1jOFkjnaemkaA+I1mph5eEi7CW1FM4l5v07nJaralFnxQwhsbAarEn6t
psR0I48RfRacFChmQNCnmj+N11Q7kqi/0gbUCkNx2Xk/NPGabBcDYWdqk5ex5LBr+mHrlKS4HZni
3wchYdJnq+c/HoUf/6Jg+djBkHG1rv4HEyqhNz2F6cSMYaFhKDkW3T0qXWz5dvZ1VKbaTSvkEPNy
kkIGjcUmaJsAaFydpjlgeYxeXcZZwmRtqdzAIk6bgNoJMYULIZtW9WnVZMadsQudiR/lh8XyudiG
zffGsFF1NpSqWXFd4kFgfD1GXsOR6NqpjgsbAtPfkbUXMC25V2BPR//hM/A8b0L08c5+BP/b/25U
U0oZ823H73C+KqInKXgQEA1KGpLG5csfbzpDKC0UurIgNFsFeA6O/oKFBgovDFXq9+dg/tGe8uqV
0XNwx34IWPh4CyGP1LSFjc5xa2/OaFNrnZkkFKgUSgkRMXj/eIJ0XYT23iTVIzg2HW+g/nCt9iEx
2Qt4AyDMSY4Lan72hCdaDGpvZTjqTj2m3d0Yn0ZoLvPTCRhO/IVS1Efmijqk4tbiE1dNuTsAZarB
Q/8TNq+BzKl3k7jCoA60sA7QnUoNDVN1h4RWg+7zTvOjPDTJuicAAT3eob3XmlkwcmZWZDpXL3ZD
wM655u+ZeqnMZahkNYlGE2gKT8BLsSavxUQUCFiQuICveJBGANCh4Fh6t1Z+dPr5x/XqgJ8jlM0V
0nL5oQ6k+UFJ14UL+KnaKHE8kZNGsqnRD3JdxuUBEp6m2vM64TDgNQbu0CUOpxa2VFpLZoJlURLW
u6SinfQOr07h1WOEUC6+y9pxdBzYbMDmf1GxlSDU4taAicrcX3cDzy89Qx8QhZnYocJit3Ja38ft
GfkeGs7QzFz1skErzwSGnTP64xtybSgGqqtQOUkAHMXRo23MWSm/Co0omzb9T2iBfHus0qFXaXVw
YIy3pDyAwNyyQY4GseXIjijno8EviGEz5MBBbrAR/YhZFpiHuVJlrnvKaOW4e1yFY5tmK8NaZJ9Y
DY5Ofp7Dl9bUN/LOKapzUDvZl2qwpTGkMjHYrdRS+aWHTenl1Ys5x8s4gXEx027UrCJtTi8AcjwF
cUUJR+N4R6U6hVjZMOlXBQJvNO9g0QqIjxYod6kzNG4G4KKiG+N+6WhVeWD3PXb9MZLKxXq72OMq
XsNG+ehk39lh77+axx4b4ljwkuYurtsLocR8kh5U9FtpgCuby1pPXd/duy0wEQf61W6O/L9UGSul
kDX9/Goxz2FzPDQ14BQICbvujyluAD738tSfX/b6NrVa2iTT0MW6Qi/61td/h+2OyjDOkJPHEECK
SsMJYbqlNG2OJcjBC3aNeXWZ3iClpKkPyktShJhUKl3PYytaG/U5+o50IteiYGdd8/UeJfHZoYQR
tIDh2wTOnqwlgld/jJeCSxHJ6MIpJfBCCiW+tj/z997EYjh5R/o9aIoFVoOE1eDhEOePI+Dj40YP
5MMfNB20YAMvTOWBLYZ0Uj59ZYiCWPwCsWY92EVc7DR0jAhzNJQYyDvC2yn+V71AlDHGTEeD0p7/
AcR2HceV+6iKhX7Gz1nWptHWvzTeqvgqLpeDN1Wbv8TSjLSgnVCYqguF1M1re0LgnHyXY8sCtffL
lDbhURNhKu9E/pz4sx7p6Qz5UkoLFH1qApdnxL8l3fTCcDhZHxy3TQ9og46wRskhtaOLxFTDvs5W
8JSSigPdpVGkkXe15psSk9bSkf7lr/5GKZBrcNYJJH1UzWm06jLp+/IrhklI5SR9M3Kv4wAhwE+H
V5n5ZWiZqbPmsTfDstQpa3Mr0ZPlQsjfnk/bMUUoHlj2W8SCXk5OA1Cn4/AXyAdB9s5Ju2S+SRls
Ncxb2F0yorJYhiC07u4ZXS7C4KtuW+Bks1pSEPTNPGF+M2gv+YQ4gsaPQqMTDl7ZiNywn6bihbQp
ZQ1CNATxvKwcdAuaKr2mb6mYQNLs6y/XOgK2Mwpvzz1npSZfOtlDj/NmNm3gEY1F2jQ6dNoekg8p
R2+h0xl5RDG7PVnynLF4c36w6J5p6uLYt8afRBs/L/oRiY8OkMCSWm4E7l6N7ihlxIk1VOauegF0
UcwARk68GZgudTearhZtc8skDWIudhxvsWZ3VTKaBo/Qa3UO0gUQKf78mKF1WKhAnVOfdnYK+fG9
444VgAtWXSvkXi4SfhMtTxyBi1wdGZmT/hYThNpFXO7lPtCD/L+HNdt8tPol5gKzBUyR4Q00Xd26
CXzaIyDohpknf7cTk0b4YagwoAx+mS/82bi0mQEr0IhTN1vgyQcGC22wJsW9zO+6IXk/vMbM4Uf6
a28FwJkNgeMaPNbr36T5iiTIshujLyp76dBDNIiZ/5O6RwUDGnZf1As69Jf8FteELh5QkykUaOz+
uT7wSwmWAZcwMGgmhjgK1WaeWQ+n1y4bGmj5aILtpX7Ez12S7SgmCERtMxVbwAJh00YmdBhG+Sdz
zEGknq/PbflejCXTrxnEWwX1Ch4kjlvZyDyMl4m05LEAaib64H5w1VntJeOEzMO/jUYqZNPtTB7S
6+cpVZfN1rAC1d2JCqpEENni6mLPpddJLT9/It0J9cF5eswI0462e+Pjw094jtn6Wrc9d3JRsQ+h
ZiiR6nuBM5a1DQ1TsrgfG9TQtz7sF05m8NJtbyozzCqzexTBWIIXwuCqlEi+r6HwQP7XfCw/Oxod
Mx1Xucywdxro5UbRqb+9sio/FNdfsjGdycsYwlGUqu7e2O2BpiKfZYBiTdSIiwIJ2+3fQXCogTsU
YWzvQQX1zgH+POCpU1syYe28//2/3WolSY1kGEnV/D5CbSNesaPHCY4Abq3b77D0nFrxdzdm3AhF
D8rhx8qKLvbiRJsXxklPm+M7HjpnsmcxcM04n7AXbrTrjKIk/mTsG9/228TbsIYtDal7WETw5jTM
TBbd6xKS5d4G+txlL3VAibZ7MmaIDHYlv9d5kSfYeUxq3zJo7BU3qL/at7PJwQLVqBC9os5CAXsj
sQ6WF1nCALs9udnHaLdTrv76PzcHgZsGkgDxmthk0n3vBjlb30lo7EmXp7Ivmr8ukLJWgGuNW4UK
qwu15+O+lV4HNaByDfAxnPyc2OdIo8z/JpXLyLu9NVYURJIYY7L0xz8xSjbxMAR99xEYBDWWKwpe
Mfy+kN8WbgWAY8QNbu7uBESRF7gzbntvhp05omumim0XU7ygqx2qmDq7Xw1Nws7UG+L/QrpqCVVt
aSj+JWzZDKK8HKKKbMyJ9FxEVB9N8DiOx7+whS6FUVAww79z+pKQ3e03HVAOcFMq44MO7zHwKG+K
PPxKxp0cqacRhNuHi4pp8qlIsFRMQ+5T6aE+CqJ1XrUhmn8UCo1aFJBXRua8INWGTid8gEgsOBWB
bStoB5Rm1Hbybe6ei5bXFNBY20lJ+CRtQc+FaDk7znwzwDcE3zLqA3UqmlDIbP3SqwpvpetCkA/C
kn8U4fw5PXfXHkuPab6G4H6zASNZXR5qYz50WMR8HZxlg2+AHQwUcaWL2DJ0qbhcgAmnryb2BDVY
kM92op7rxqICG0AHR5YUbG9sIH21cD3i7oo5JWQmJJIWplsY+Qbgh3pn3dWXUfVjKj//I+kRbvKv
EAk8zd3CFgyQhSRHbEP7xktUcLnWdHK4Whvw8LsDfTaFIsQhS/jZRcG5muhMXwfRudhGhMfsMkUd
ngVCdQzPc4ZZ9n42lEOIWH1OxjzJksqlA6D1ap2qIX41qGWQgeqASG63j5Wpwe+s7qUkgpJNeUvH
OZ+B94KsuJYyvz+qU8qgpP398mNT1kIWikCDbUUa+5Qkx5fA7HOy15W57MTGpD5MnooSv8eYBTpj
gVF7gzgjBOa0eUfB2v3aGI1qm/wT0BmPTMAI2HEhdArA7vIxOdJbNhF5L6CPfju3iA5ceXizRjqC
K8gFVccHXaxoQn/efbClJYP3Lj2yRNiet8L/slPinIf8GUBP9eiGJx0Y/E5XkQJojZ2Cmtopkh2C
ZcD1MFKOld0wajvNfvSRD/kwbongxO14vVlpks/Im5jqzmcQG+Jp9250UykURrWb5R5kwAUio3h4
cIq9UOlG75msz2bxeeGRLiRxftY3zBnsLfrCbJ5vAt5zO/bSCkhlUT0LOOrHCBf5tud75Op/MlHb
onQ/gxSQn5vsPrpvgSKIN53UxK+PS726L/cKxEtLr9sGpclhRko9VihDcy9RKkIu1KNAtjWCjFpz
Q7v67M2uOvcxMRmZZbifOtH3XPZ2F33IYV8pod4xc86zT69r4cmAe64m+ANpetjLZOoJ3UVuoIpD
gz3BnKnmSEDlDZlRfjMbYDSJSy0F+6eJJnJ5CZbTw9KY9q+NYhdOTxgVZ/tztxCOKBoKw0s/ITxL
yLwijiN4P0Gf2YOtOMSd4ZaJa/nf7nuKHs5AvSqgbNkSi2JuczHghg2h4XdOwJ36Ep69DmwVjR01
hJcHenpxjuIUxRqysP/zmVoLwH9VycLGNiMP3J5cMhS/bOWTwXS8/oZjMt2hKgWvfBt6MUop9VfS
XJhUHBDH7rJklJatlBFduigBRS5rG71rR72PJOdYdbYN2Rhln5+jt69eezGlINQAlCSXHv++tCch
oWw3yUhvZSjHdpvQ53Je1SHp+zTlhmlj8Yj5YX9C2kt97m7G6Y/QbYl3uWesTzX/Jp0CaX7HH62X
RT8OwUCFQ87/1b9DxmNdJGe/uUVcKd8Gg5xzoTeMsTRCptG+waOM+Mv9nQwr3KFC7NSf38oPaTz7
C/tjh4OEbryAGO0k3aSg0tprDcTkXFNXJ9qDmJ18MmGnIZbgMcLQEsrxCf04lSSSbxjQCccNCXWx
BeZ1c3psW3Iyb/eVlQiIMqhmPUTOVc0gZzKIgIlv8dlYJ6xH9NuJEb3GjZfmRR0WmZ0QReC6qhMO
YuUVJOAu2cG+YUuaykl89zqTCb5VFVejHVWH9v39aY9O8h4lm6Ihn2VByq2CkHUbYQBqzmcmTQQG
Ol+k0xdIy3Lim+eNsamFcEGxb4N78iaGEilhpLwPg5RI47AmbLD8exkc6sGXVEmKFF46G2JsEQ4E
jrMBgMRSmtYYg2EpFVhw5w9VgQej3qslejhnNdfgupfNxOK34al9bjTeaKZbS8BRZ1yTpuZyOWBE
XwF1XuFydjcEsjDzgbPEsiXcK/VOcqe4/Ew1N2lWWJS1grv6lqplcZEm1yPfBD+A+xMh1nibxLqT
BKGexLPM5beYhcBTd1fVfR3AdciY9/4Au5N09w9g8vCBm63Q/D0MjGfeBaWOp3O/xDMfP60ZFLdm
fjUIWrXChcu/GVhFJDPvCCQIkwQgMxVoFE9AM25e/+7TcZ8PDdJDBRj8KKOoWACUE5CZC4QYEPn/
JoUXs8tEvhnWePKJyWYsnsklz07JCKaIcYVtQ1V1bH/VTNn4cKaxd4+BqJpPvgmbVnW9PLQhrolP
PsJOQBvzultULUzoXLW/VNdEbSxRO5EfSUKpWfVoIwLKnkBOm7QFeAY2BZGa7wGa25CYPWiOReFw
SFuRFJNHgRjVrvxzwnJ6/aIjUSdUiaDERe3LtxhjGzy+OKIpF2dTi06R12fb0u73HS2z8MCVYoU9
WpMfHjsIgq4xQtiyjEK8989j4UtuKudNuVY9Mo6AFJ8Z7c7WUZtAiU+zHFECZ+F+n34XRPfYxCe7
oH/mCmgKYZJRAGtRAbQp0xaShFp5KmVUD8AYkeTyOpthaC1nYf0G+cGtB+qSUJCnthFO5gxXdxfE
qHYoQxDEUdghco1y9IULv5Okjwk/earHrT10FpxdWzzcxA6im+C+Vz5BjlZh756aIOXAngQ6OwSf
a7YWYbZ/mL0VPoClykWJjr/g7OPwA1jH10GEHw3CxFTyLBzavJwBfl7jrTgYIkGDydghF2Bzwi5G
KEeQVZAA9PhBChwa/LDxxWNGA9nz2BG12Su1mz6FhAkEv1T6ypH9Diwislpndx44iuCmkAXwwyEH
ExW8vCUaknr0Tq9T9lLOG8AOWjOO1deqZIv0HeGS2jUqY4dxooIcJOgi9cCT9HbqmdL2oxbmuJOU
ruuPdNlRt37pITJGXsrO13P/Ym/tmDKPXkJUPp/fvQI1HbJmE11ojWNbbkrmndBRlr9KELWybKD8
O5Crb6Yi3qEWyL+4GjJKGtp2wEMuJMnBmrsBfnbauf9PLW1nhEeg7kkMX6suQxkrnYyxDRfKJm1N
BgHcH62aSdOzaP1eR5hLSp70G5Nezhp2+t14XoSXnD9NeYaodEC9d5dYclqsL5ZviwVWbWoErAqt
fuA9bGMWzn+z4Dy4wXraGVXYMt6KjYSHkjQwcSnN68Csyy4zJ5iPM0guwMFVSGd2aUMgcTQ4N99k
DbTsMg7J+0VemnGX2amftULR6EwsjB8KO/7tU3XCHM17SIWbCZx6CpUwPuwbT0JpfltbaBmi9K5p
OsTqUcVUwdUI7GPZslGw12KipNOX09WVwMU++dkCxLzYoRrF7ArcyG82KNvVjZD551wrSX+PuJlC
I9vgezyiss5BwXmxUiY53JEx7wV6TdXZ6vKsFA9SFP9zIps463JtLnbzk5UUmuPYQ/xKaAi6ERcH
WLa5q0ASSjx4GCPiyUVyIUH2ZBOCM3HCC1IZVXMDURLqY70AchXAfWyj207n3ir9BhdFI5apaON3
3Q8CPgrDvPw1rich7lpR+rnjswZSC5c7jPZYwyBn7HBrfdfqqGvlw5EgDABDGaRHd+EzeOKWygFw
5qCjjUk8QFOg9/3xO3PT723tIBdKyVeEuNElH4M67L/ahYhzoFX68PE40AJoZNL7LuvC5HnIEkH1
BUMILRm7DkvXDVk6k6hCMagWeyjCVc3f0+foWafU6tzT9WsSxR1SLL62l4C1hFafejKkTjOR9Fyt
S9jzfPJ/fwL3bpT6znj7SGIyxlS/qx138D2x1JKaeVwK5usCl3gEg6I2DMgBCkBNHw41HQH7Pj3P
w6t7EqrBsbfDmDDkox+wfcWoUHN0Pc4S8dgZC5EnCvrlr+Bv21rt4XIbzBv/nUy+DRDlDJfRPIoU
Hz6i4bCzLMUgh1+EqzySye/bacp0ETpqzRbBbN3Yn/BQhX1v7h2Gk4ajBUsadkrhPCRCBAXAR7KK
nc3hz0/Bt98P+1fVABojg5lk9xf6dG0rAIhhlfQPuHGayD3o0VdiTqJExFN7PYn4e41I7UNQ5xnm
hh2nKiEJfepWLGUfTRGpEMvoamTQr6YfR9Gxg/DshLi31EAH2dCElowTkykt/nsYp1UpwA5kNyFj
xsaI9UUzdDU1UwJTY3BfZU+/JeH8WTvJhLBnzAn0DBLXq5Z8YgQxB9Ln1fmqZrEE7Lkxhip6Uycp
b3j+5XmZKU6OerJxFUyC2BAZIF90c9txYYXfuZEocGK0JrTDBzhEesBe7p5SMaXx6h2S5YvOpCCu
Mk9sAYZjfjlWT5cxGDdnxGN9heRHfChl0hHoqifoZkgrjdSibjnS8SEv4pZos5gMjwknGuS3PjY8
06l41mQylIqaHgLjAKpfX6j2dVh8c2WcuvYNKGXaqpNdj1hmurM+bGOP9Ip1Ye1Sss+EK340Aual
PFQmu46Z5eYXaTLefkoN4Mm+qnqm5HD+BM7ZzVH5QGkeLn5yBuxp5ZLnCfK/1HM6AG7K3H1VHodV
lAX5Fvk42pwkzTxeVJRFdh4P51O28sq2VBPHwmSrAH46KRjVdruH0IGsfXOWsJPBeIG7Xst/p21w
79J0QNkHAl7LsdGFhjTMUExTSk8GCWWwajPqD40d44Yqs9Pzdr9OqIfQVZsazWu6/iij3B+GXYpF
+hG01zXtGhfj2NtsNxSv/xZxeVBIwHaHuCJg8FMq6Z43MU0chZUg4gLAvIIXdUEOcCJmT9ymwXoi
JtO7/o29UQ/MN33xpUB6mYa+tcQb2hewxq45I+n9wx8IKiSibh2ldfVffzGOHHnnSdqjgJhwP3eV
J1nhFhR/Q2qAiL3o9r41B5GL1nNeckartof1CRV5ppQu/irNutnthJPdmUudB1KV1K21PXuQOW8a
7eosFLfAFOURjQUfqRF5MMloo929NLzOBQtFlm4oZD8qBQMGOPrZFLR0EVnOC45gmj/iaNd3yWIE
kvWwAXgL7kzE+9DP2B2TkT+cfNYUNJmR7e0T6Y0WsnkzVxjaqhdBvMPUTgRUweWt/seNBqOU6cOL
cbJDrTij3WN2gQPCWXBDW6Tq9E49JLi0dUNrFGCxUAOUuRQ3dvkEX1/0uywrWwvXUJMJDzwNXzgx
gewWGB8WqkFeKpklD6jOOfQ4/grlwDk+yc6o/p+uiiYD9F/95HdrDgP4o97uw4K+tR2o9LB8b2Fc
Xmehdy8Qfudcw6cgvAYlfWdGIQyV7bChFx1FIOYwleAim92+mLhP2EXw1FdkhQXRWtluUixJ9Pwg
hrtkkq9mdKtYCxCalRE4RRhknqa5fRht+tKsBm2YPlEmsa44EE1al0GV1q76BUdQAovb1FWI6lah
oIiIioajOoUdDfppBr3oyW6lNzu6tmEv2+w3QeZ/VDjOrHVdfo1I1dYcAIkc0XdWr9r5jw1vgWJz
W8NscZOLb0rEGsA/pECdkdsjpMJPeK5/6BZQLtg91wrvfX2YRLAz/T6xxEaL0e592ypBAGyve3+g
B+Iy0XKiYn/cJMqw0MAMZXMLkbHGnWf8gP/Lu4gMPbmO6OkYQCKwCYFit6Z8HTaU8MzA4fQWAFGd
tbl+dQELxSv94E4aMHOyPdKH43rOnGrisWrS8oKGc5l+69Cr6v2Qby6/DbiGMYb4HqV6bKaMVRfD
lZJvu9xBn/deyKRWXk4jnfXeMDHUPy6zDpeVaBirYTRNh7WKhps4ztWDPAXjkeGj0HaP8/Va3u5+
wy/MyCipXQmZbW24E2d8NZk9uOaWi/d//LBw6E5cZPpuO4xq2PY8kfGobqzLpLOwDB1SI61qx+Er
nWGTRemIHpVTuBN7a+155OfeLG1ZaXzDGUDXCp5pkp65H17ROf2eKlB58fprvVPtSBGjuRq0pyqO
NPhJtYtp2tky4qK+Soc4DGJeacO6G5bRaJ21fY2Qfm42O1nIKM4G4RASv6573MAb0qXOrV5zQeMe
59Id3CiboxYJeVFA9tL+kcxZieX75HPqBrC/Dh7TiI1Fyrrdwn0dtlZ1Boo6R3XOB6tBcqKi17mu
H1COkm5CIK7F7fxDoSGgLhb7KWhm6jd4r7Tjny+y+ORh9P8RK15iJT7v4tJmxm1Ob/C8Jy0Yadxm
PxYPbceaHB+0D+vo8MLSkG4o9pvbVZz5Ls1JOa0Woqc55YDRR1a2ZyxoafqIs14YrMEzIQt6nYFH
bL4ijHjm4gVqVA8gwOXGFxsmcASKBEjo9cA2B4ZaRxRpPcHoqTSXAYEzr4bEWR7IqiJMw7Qif57w
MjSnr10mJhaA2ZhpPzoq5zbfSnjQay7HkDpvjd2s7say9dupNA82b0nrXeqqIyC1f9F1FcCv3oiq
9Oaut07EXSrEuC6tJU+RPgTJrU0wgaVJGqcwDGn2ig1IBfy+jWcraXps3Iys/Rq0wHrt4cExYG1D
bqwjVY2PU7rMZUp/kGXzFJQFjZkAjKsm5OKkKF/l/K7NKD5R15ZOLVWx8ovwIyjYrUMIpQt+Y2f8
dkt4mDnkBDmFihp0ULWNBlLfUZUjCkugm46L1orQLNfUEemEj4NJDnRxN1KwlW4Bo/CHrPTDOttt
ez6QJhEvEdT+uws10ZzOjLJ5Njr6rgkUuB56DdhTNN8BZ+3PR35jVsYF4gvxyVpAAHU6aPS0K1RR
DtsAXNy2ti1wha9ICG4otreRxdNBHjafQ45SKrToxpCakxTFNtkT6P2FtnI3UY+CUfkE7iqgA3Tp
hGc9+l1nNwelQDUQQOrvyTrkyYFb6ZoL5QLyZ74EIwLy/zJ7QYn9C8IDcHkDpvAJnQokwLVFLuRy
9MOXH0oU5hTr0RTDQWI/u5MeH7ndLQ4rPhR2ZDnp5F7s0/pP7D9MURFKu2jTOAdSvLEu0QkNHOo5
FHEdHJEm93hZBRfEzPKUtxe1Xz4VHmSu5MCN+K2darpI13id3sxkeyHmMYRAm3DoPtdS9/HlVWPc
clv4N38IFn/n0DyCaL0w+DFWCckVTzz8CysiN7MmjFiyFMyEyj/jSo9hOmKgmX39DvEzhEYhqEyb
E/vV7r6yTw4utBUs+1ToFnczk9uUumCP9DImtQxjNK5td/UFh1PZvvbDW4m7B0/9Q65H9vo13NG5
6FBLr/XrsaJVaPqa+42hqYH4dLG+5vjfCATGVm5KuBA/vlGGdP5QW+8xWQtwERia5dntt+FIbAP6
T0w/mixGg0y7sojPX1aciWDkKzgPhsdxgTxKbOuvLkkVNMIqM4fnNUPEfYERPpxZx6u4txnigu8A
YIq/+X3cPibK5ClaU5u+0yuScY3daTeApHyE698giTQn5bB5XA0LTB31AVhnCQ/FL4cr8BAlf014
LAmD8dE3B2dzDWuRJf0ZqyxlaXoVfX5qT4d79OkOCw1DDUMxRIPxKrSuoaA0vM+K1r20I1hkJ8gj
Gl4lEX1Qw24+G69A9x+7AzsxP/jtCLjp7vQiNyaHh1fd8w0stUrRFf8CiORTCgYSQSWR2WjFmtXb
zVg9ky/YM6G/8EGdTXL7LXLWYCBJlgANCBCX2aXRVcckTOamkbHBzrbR/PU4c8pThk45RV1b5Qfd
EYTzKLdhvqcC7QKPb3vlBPSOjTTnt/JiCM4J5nP9KdY158YNpqv1vgbzy3qCvkwNNBWSGrfyK/hh
RAuMevx/L2UxSl+aMcbNWPvmhFcthEA7h7iEkAsb8hhpOyYYOrOsmfbKgzkkuVsat4Cgm1JLodQM
JpFSqJwclNtgbLahVx1eIwrId/OVyclOf9z1Zc0CRSmu86etHCrd5Z6P8I5BFUi/YgSlk/ibCnVB
1HSGW0G7GaRT083RbP2UMJfd1BMg9xVppmelTznJe81lLcUAkp1MRvMviRYWZHG94geq78H4vwe+
dfp1ObFszSjB67caEcd+WduODjLoDY6PF753FfhIB18QuRRWvA0oJ4vlTNCsZo5zIiCkEdzfnZ8L
ETni8LVUHQkNhJI+7h4kCKijC0xakpbj4alBUn1chaJ0keh/DzK4700p8sSfvL3HtWJdWKJV4+JK
bKjAk7sEi0jOFXmfNwwAWiKCMPuN4htelXg78R8sqmVcLaAG46oD5o4U251PlJuxUlEYjA+8VS2S
JOdlTVMgzgyrlWAt0OO20pzw8CoT/A5RElaU/OYGKw47DJX8Drf5mq6Qt87VeHoRzo6EKC/Q9yWN
ZGEwHf8WoWGT4vsuJE/tzN4Iz0QGD+T7jgS+7mRo2LtJ3kh2D37+AmnlhXvrlWuf+qJHI3V7zqp9
4uNHuMVk6FwjUL9O4AG8e08W6mmV41UPnY/Yp231OC2HqBOz/2lQzKgHrV1RYpTj83YHwCSwjlpv
DTzH/9eSv60DjacSSsqNXSoByVsjbwV07ngHKxKaMGkwDvc5SR0aHu9ye4P6SFtDeJ32wfFiKNaO
oJne1ucwUqd9UECTZ43yNE4bxesPZJEcol5OISn8GyqmUUfzV/XRsI12OvmU099WAZTuHiFXARyb
PFkE1g8MyrzeHNY5XQ0muiwoteEPrSdLrCJ+CLBsXxEjpGg36lBsW9TwGqk4iBBulJYegFQpqjDV
qz45HDRox3cy3wAgoKbzIQDOmYWqjvHtRTyBU5N51vRoDFfZM6NSIy/OKygOa6SmpKrAcdmmhnB9
jg64WNwcW9GUTIC6J9ee1/QYEHXLZz2aN4vNoguTAN0wtBMQ1EeHsugrG3SC83MTjkwLidpgiwBb
l2KCZTu71aeVCRsTL9oPuQS4M49WmGVq1tXX7nZuvMllg9orGoTWe9/RWsfYK7sL7TzJMr1cKI9B
6/fx1jJ6i/BfZmVxyuxf7ZQcU6mzyhxD4DXMpvWTBBCLVSGSO6T6G7Y10ncE3x2ZPWpyv//q6Rrq
01puu7Z3tp1zkoaHXP6q7sLrUpJf3b4Kbqyi5EiN0XGMtisIHXNsX+CkqqZHo1EcDMls2il8tAWn
l9zV+/Ock8BBri72Xsx/QB6RgRRc0MqMJyv28yCm+KA00CKmQ1Mb8g2CvXl44cLMu2hCGYSF5IXq
ZypfF0ekXvccmilF8Uf4dqBLhhzM0TyLkEDr4NvqDSqwOG154Z0057JruiZLI3hM2pFYNirXO63M
wO+XhHiiNhy2jz3vJN21dawRMDEtj5vELFQzZJs7WIJ8cMXG8voGJs7WDV/jw7XeAsxWCf+06P71
xNl8Q2sVl9nmfWh/46JH16YaybdqM0DFRTpCAtQ22OgEzSQxSg2eujwTfg39pC2NSt7EkfZcNowL
J5A+wznrpjTtRNuAu6Flr1dUiVQvEhAjbDTTgqN5WogxubGDz+UHvfZL+49T6ojeTCbLEOZqBxK1
e2bVT5WLwMTTk/m9zVWfR6FeCIajTxQO0AOc8wroTutjKX63mR5pF4UBSd1yX6hwmrsIuAV6m3p5
HcDImgvTPa2qm/VMWlmJTiu5Vi/JKB6guygaT/WdDhsVoM7lfQsbAPGuD3vVj0qS1d8uE+/YhbjX
KvmD2VQUDF76OGK4mbKv7YNtlqBFen4UAi8graMQXuwacteZnJvkCnXX01HWZBQ+ZY+jPANgpVjL
tNcyY7q2Bu2MPrF0etz4Gl4r8VnAmi4YMu/lddRGDwxTL2vLTn25cZzjZqw8MeX9pb1ZwI/OFyzm
iOFqvCvlLlD4+Aoirfa0L686upax83tsoBOcMoXN/rnSQKmQ26u5MXT3AicHurwcAFEHTbAqHeeh
vVy1OsUpvY0PerW9ZTP4AgJqzfmpnQ1Lx91zvT6o0WkfO1p9O7dF0OPiSxNzu3aj0k2KRv55bCXw
TqNzsn+N34Ecd45LxofpoRZ0b5IJh2ULKn/oDC8V9hHE3P8rtl0gyBJeLNUzY7qI76bhh76sbXH3
bWZSZ3xjWS7U7exE+nQher3w5ho+pE5yhxoRyxCGvNgDnp6/6siZijd49w+oct9L/xwfaS6K3TiT
c7S/nmwdGntgCD/uYoIbGjRSp4ibqFzU5T8p5SHE3meRLsLsy3F8xcSFW7IFUUpxa2A+Q33OSgRz
mWdXwIsgXJw3RteaUc/pDbAVj1pCieuMjLCJNBJaGJqAaWwCCcHAoiJQAVWXX22rXS+6//+fudKT
NImAV+8obW7IdnufkTmVtjfT90khv0DEEj0MUqh9APH6sJNqsTlrOLz1wy4hR1WoSJEcF03Eq6mi
oFitVp2gKbrQyeAL9vROGy41mIF0PpSkN6eShT4vGaWXsy9EdAicGyxERsEER8xlTUAIIMpGHPMZ
/7EWGwX8bLmCt4GsGtgTporrmrCtnXxzRd2Av3Ir1yi+wBcsRrFBmKpG+rnggZII3ObZ1wzVcoZP
XpTL0AITcEtJxqldobpLKbh4/e/EgeHdHYmxtpx9UmZleMlpKw2uo4Xg/A1kENpswXAm+zWyunU1
ESi6dm77TVXdijueSLEenffYrOib+kNMobBgwkxUSTVGMxOd8www6Ziejyf4EYTRZw/bM9SzO/25
m3g2NQaKhy7BMfpcECb2w+58UeiuQJLYvFPBkQBZHLFr2t7nLpYxAZTyGqATA/9yuvDk6vOy3MUt
zMqbJ7SmaY6D6h1EKuez7O5tHIifUtT1GKn02+dkKHnwVTWFn9VJIaxOUCz0RjlVEwkt4zGPegPu
M+8enz4LXMB0c3e8xsMe0rv19f1ZDeHBUo1I3D3dJfKJHEm1b/77CTltM/t1PT5hGRF3oB1Bm/gk
wskR0s1vZKBRZ0u3ybhAgZ/ah+Hb/htM1CragLZ0lBvpi6BJ3g26Ae3jv/5fgRQ50J1Le+hxpUcf
uL4n3GzbXdAnixC6ECo7rZTS9a2VCM8Hs8zAtofRS3EQhqldiotKMm4eDG/Q8c9TqCDmh6ZlUM5k
safALx3vnEi7g4fKhe+B2EwstA1gWrCAMIHVyf51cArQyfKcaonh20VUlhDKD4Y5u4YHDGgRhFR0
EcQrdlCdqsiAUvGXvK6FfPlWYDjD6r/Bscir+qErE9kHFvKXbtqKRqBwY4wZizwhNtUhwHo0jalK
aPHcZ4lpvxN/yYmpy41s7fG3N+b6k6uwlTxMgDl8Hd0TDLO6unbeXxP4cDGpJK2rvh3jIGP5tEyF
XhfMfdwr/dlvEtz8SGrO+NH3L2Tzoil3nj4ZVra+2+SBgYteaDMTF7G3zbIzHMdzdvwbjlrvu9EE
Jl/oJ+p7dbmpo/gUvdKgh5oQv+BQeZmVwlEX+AmLIH7rJPtVssJmV+iLbhhlJheX07Y2TyccnTJe
rSkRnqDgFtMaO1UWD7y1C+bs/10/V1DYbYNEFEnbzr64UHCmxBqKQ02Va/neEDTYantOhf6qB625
DwpMk5FRJakhZe7hvqFiql7N+FHLl/GAmfqoV1jtATBXzCNQ+j/AleQDmHlMqygjGU98EBLYgRwr
8/mcjzSZAlhnR+LxdtDsVCjxWRbzsfszELEEYYlQO/rz9hZE8iU6sBtcl6RlKeaqKONd0Wfba2Ak
RjvGBXfs+HdKF8MGXS1vw7O8cium565DeSAsGk9cG8EPKFdh4k7LfJ+AL/hHAOfukKCQ6KJYDmFS
y5AMPPJaVvKhS7c3AhJrAMEq1TL0EZSX3/DQx7FoHBYKi0kVZ2fEqWdMEsqvWpyhBxBfmAl4i6B7
jA4fqyJjz3S/lL9j9+wkNMYpejoPw/pq+/jrpXqUn1ZVuQDfjS3icRLMXnSrF2ewEG67QHf+k1b9
tUk8UISBgZP6YyxSOc/BX/H5pngIXT20cmkPJRQfMbvhqmFRitWZ7hpUVAFO8WCTEMreBNTLu4kk
c0V8WejsiPs4nXGc9dfmqe72c/b2VSKIuXLrYsRBVp0VQSVUllxEGf211CfGghgpaao1KU+mZAGJ
s1q7fAzkTLpJuAutZrC80obNEbjl3pw3OsajxoIF1D+1Z85jJ0CokTkrgm7SmDxYVVOPNqDiR/rT
Ff1gWEQ11CdJVRgMugAQUbWqXzkW6eXueBQTvZ98c5Nw9ci4dHV0jpW2yWznWNhIPZmubCzNHy7x
l2couxjVo8xkjK1s9uwQq3Y65cfVfaxyDwCJH2KU+2iFsH3lHkUbyBd1448qmWLGxlQQU0lWdWZS
3eGsOpz2sM8Mzh76ZScJTdJC2foXM/yvVq5JCl9EuY2XCBL3WkxwVHzeNqNz6EuFy07LFqFki/zJ
gwS+FrQqbzsUHOnro/zJxjtTP1pRfB43F1kPASmXT6nG2Esb80ybcvdZtvqaR+nkO9w6QLmpDu87
5XhI2ScWrV/C4361GYHWDpo7867uGbNfHfJOHsDYjkjY55UJhJNUV9e9rGiglXyFFegQEwxt/EnG
9MvYJJWoEJxc1XtWLyuPSqAfpJhqfmoubnmeDlQ8GpvSoqIfioispHyCwdDe5wDBP9rdzEKW+IoE
wbS5Gy5tuDTR+qjKphFCxT0EAGbfouaoQ+y+rwSjYAAu4dGauokCCgprIl81Y45hI6ENVM3xbPmS
Tp8YjpuBFoItu/yex3g7hd06CND+wS3yvlhe/SedHUbgFlhR9QM6wNO80CTPtUg9FrB3PDrodRzd
0mOWWhQU+5SlkWh9N+IBwMD4AQHwUa83Qmb/9vnqm1nw9W8XAl6N+JRPnqpDOKQlLolvNZz+sU4d
5uTR2VmzFXo7/pB+eztqBR/JMiq/NcKReWIpQowb8r4vVV9Hpt51hP0AHqrpz65NMv9SuaoSZoRp
XN3Gy9EP0QjoRD6hYomXtLMevTV4Zv+gkkVe+NzCPOLucTtbOp2bAtVfmZb3hsoVHsLd5t7UOVdX
2BBiKJu3nJAdajty95brUFR75l9FUTpdPN7yrVxsOiTjJkHQgv6wPBwyErc38IimyPthpKTFgH8n
9YN5ikHwDwmJr7R39fJTb7+xwvBZLaay4YJ6cC6TD7OzX2ngYXd/8R7/es+fclgd/r4av2Bh3wtp
PmQfyBIDKKhgoVreMBXC1i0BK1Npe9MdneLti8Sfk9WSP3S3cP/2SKq7XhF+pBSRgwSGagGm+O+9
+IYC8ERMsa8EXajMPLScowVTqtkx+M0zR2SXryS/LGY2JbD6WFOf2Rp42rDeRdP4ROCGESZEpl8q
A0iJeC/NH9UouykVWJd7emPCkgbsmdA66wIfoGu9y7FSv5CJ/L1QmuiGuMYLrGIW/5J+ElIznGDO
59edVAvw2i+/rEvqq0Z4QHzOojvR+9gBJT8O3Nrt32O59jtHRk6quOSdO5Nr/CaOGdcAUNDM3TNO
Tyf0jpeLAXsWPsrdT25q/9qoZylwo7nBkOZ/FWPupwKl79Xr1rxYq41tQ2F2raCfTtvqGESLQZVn
gqvlGLqR7E6SCG1QDK9sWmTiXmaiaxYKtdEPtg0/QZnhoWulZkMAt/jIpKU+c8HmgRb3kHelNb/v
YTKcTcMRJgMWVLCYV8WQq2NNVcFM3M523H11xpUi2765zgDUk45WEoxjFsmfcR/oZu9pKMd5TbTD
EcKzK9zTsNyVjkNVkqgOqSLU+csRDXQM3Qf2EdfWVC6D1VW8sAzhzPUYQ2HxYr8l31BMwdW9NH57
3SZ6EsziSuRom2EGHgtNiedFYuWAWw3dC3vYZ/NtSx7SjgJazgH/Gbwk4y59kRTO06iYFzpv84fk
Yjc0mpVsrVVVnJcaeHgLN5rg5520OVZKEsFcM7f5polOv7naDj4gQ0ATM3KRp3tJmNAEjsZz0wgw
Kpdo78lUGxDSSqSA4FYi0DDEsCmdifjRiqwtQrJvDuABPOiKMvgPobNw8uPsbBh0uwFtaXFqPGfg
tyRQ2QIBSC5vyEQFEbQOVzZ7+QKmuynNc/5ek0AWDN4nxX9aIR9b4nP1aOLM3PYoi5WbQcDVEwUs
xxYbhCQgxHDV1vjEeyNtsv1LZIFrova0Z+iL7ygYGxxCzFm4USnFiuoKe+n66/Rur6JEW6ty76M9
55VMtmIoXZkYoe1VUqNG1EFTNCjah/QvBP1OnPdosFR8ezcpiAMhEdIpnpjabqeQl544bW73wwRe
0MzxLuhtP1MZ1x54KxEubngEliW4e+sdV6T3NxpGW9QtC2Pqv7CgT6KKJqK5YCT51rsObA0eaX3E
ZRHNzOQZextAtaK3FHp2uZlwKXEwKYKcgJecNlZDsIpkmVIF8n6KpFV1ijawCfwRMdIpzwvjuZNG
nudX5QQfjV5hjs578y4Ltnab52FSQfB9jg+iR4IipSIKMBR5o+FJNbGRdKAQk3IhiMV/iMyEB2Sp
u9zxsvIrKdlDrnzLqeqwBrYbCqvKOPYPP7+aWST3vLQ0KyxH7jtgLVzFluFo7ynA6g1hlq59u08/
60kFk6zWh5M5CDWU3mmUJe6yXwYXsGiZI8ZU9yGKJozw8PtoxamJS/oNvWy1UnBNfEz+/CJnCoUU
Ri0YclgiJcGBXWohLHfXXNJza5v0Fy8PsW7W5cXAGuEu5SJanE7v01Ojr62R6/fhtZOHL+er9s3U
7+xdBS54INQUgLf0Aj++sCZHovRZBg73RRz0HCLfZM4mA/TNsmiSDbwhQYKsan6uG/9vmHhjA5uH
nPejc7YJhu20RhAElVQ6MiAbGWHxhu5Jzwo821qsYq3ybBr2e3nPOsjQsPrRPF/lSXAk+NMZiW/Z
SGTqlQLuZmRA6ERrhypOkQNmWXmsO4N+bis3ziOkGQKZA0211t1VRl/qg5FEpb7ga7Q5PlOSSNeX
K6tsGioJ0bLvx4zssVkAlG8VdvLphS1UzL63BOw7Y/l7WzcvTbL/tQnev96+iVlrx4sBWIQa5nmV
sMA/n9kAYBjRhYqww02jzMbGiIOIXrjjsjsggRFbgK2C5eQ+j+EXabW6/QFwahVGa9ubopZfYzZQ
Qu/u12CY6Cc/0gNzP599t5gMJmeY4CCYsxsBqn7jNxSwlMj4CL9wUep+RmYd0/Bok3Q8gNgyq5uc
7y1ju8DUCaMr8JV+Q1T3dclnyAnqQdiTA5IvLlTQzWDeaMD6MCu9Ov5SSISFl+5zvWAWVGu1vZEn
VmFfn4YUE/JPAaH0Rquj/4h0WBLwY+6P7NjeBrGacldkeagA3X+LaQlz6iBeZNskZp62+cRqzIvu
SeUW7yztgf9ByMjUe0PV/H84326NpZRZvknYFSu+E8WYUzERgGGB8dbrzT6nY7HLdPXoIeLjj4Do
PFSu6qq183JmxdDRoKSYMIY0T5FjruOgZId4+VOZA1gJ/zFn2WfjXRTjp/4IBLKZRY0iWjT+j8K2
6GspTsbSUtcYg7roPkZW67LYK7ki2L3MqjEt1mZ/s4E8iZfUa2bohJTA10lbmlDsRMeWHi0vBUMN
Ync1/rnvDj+VF1NCvDr7cYZ/KS/9jO59YxFEB1uJc6misqu+RihPklLo5dsLZ3fHCsHBxjfG0rM+
UczJ2ePP4r0PKGQbOA6WleSc+TeKkTp5ALLce7OgErTbBkPkIX7ym1kOgF1eo22jKc1ZvZn+sVCt
VsOg4wbq7AA6W6RNEtJctX0ouAiCAG35lHNRJmMF+FKEdVgZ2/egT/CFKrVoxYxFb5UDgWwEJB01
PYVe3+vXcsrHAjW4No7AzMjfS++YDTeq+kN0hoqUo4yaG3Z1W7nKG9obZx3hzaT39/0i/uQ9NmGp
mgXTRxeieAIYQHn4cutMvBcLV/Fcp7XbXhJ1his3SPfdgBi+gfO/EocRt55UYnpVkIHupACpWW0z
WUJAYhuvh1pffqVBWHHFrwKqe7h0zPsUTbmt9P/bBpEUhGQRoJbSyN7evyJFGbcnp1dOzuE+KphZ
lQ41C2boxYAaxPH7z3oubXAo3GgfQlbgsMIxAnIpenuRb1Oy2TwyXIlKM1lD+SAUVrDtO8d5Axl5
UReLpjfcfSyZgDVSOGqc/s3DJUT1DIwrx9LZipLrHP8sZjfo1OBc2zbYA/pnQrRl73TdgqiZgidL
mNbcXcBkNR+DCYZOvJRunmB1CezTpZj6LFFzwArmgCOL9Hr0LiZBTu46KT2BgvvDJ/QrFl/ew8ui
dFjw9Bq36efmTlNFmlfltWu2Ng9qXWUukXA3aBWHNsB/4mAT4lRgUmIe42jLVm2XDOaQ2BrFN3gB
MZ1XWNK4jSJwZSTifwTXev2XwoEZSTse6AWE2d3ZP5hTRK9O6qUL7INDw6QHqWx0aH+9Ttal3wg6
G2qfS7X1j81nvft7SIuASM4j9WY1cPocLsL0/aNhf2tUViAKmNXlLOBwXAecC9R+VNzL849DE5f9
qykfsZ/Z31jhXJH5RkvmfDpByfbS1ZoBAXEuJ2CFB0pNAg/nOLPCu25ojXmPZ2vF+iprzBWmktn6
CJ4kDm6VITrS6Wa7GtOBGNixgx5Vlv8s6qGswieUyKzegWXHSMWrXjX6cpoRM8XNYFUJ95NvLPQO
KBbNP4yukk5HDfaGyrcz2oVj5cl3P9kOR+o3guW1S+h2bLumEW3OIEELPjT8V7rZFBk6xvu7m08Z
RdeOrZdA/noAslXpMvaYCS3SsQISB9B3dIqfAclk0DA393f/kYwREgV8a2Jp3VVv28eceYmvUL0s
xRnF6L+kKWrh0BMJ9ESg+U8YfMpy2V4mb8CvZLQIUcjKKgDGNEIbeoug8oLEyKHTyIPKqcL0UFcx
cRBTmwzFaMSIS7L2BxtoZCUXRvS+v4/VCH4/Xt7YEoZv9Ws9x4ENkqxrP6Yp49ebuzo2iXzbwka9
VEhX0hODazffVzvRR+OESAco7SYxkOruAm8vdzfBOgVi1YopaPdXBVnabyELUTPlRJOCS75Fqguh
nZ4046uNnniIPRI9ZmjU/P3BtGbtP2MB0yICg2IDCCOPH42/Fa+wlRabdFcNbLiIhSA5KDWE9pNq
jc+Zi06qKbBeTm5KfUL+wHGiIs1R2+q7/mrUehTmMx8wQK/bcq5nA+uIEiAPlk76EI5UlaPgsl0L
ZG6S1F2Krb8Xho7tju+YtWRUqUsTaCxDjQTMc3uWyrEuk44p4PK/1Xqpgk/MV/qjXAtiFHZsHC8B
H2/1vPiWyIUX8AGse0y6Yj6WwEW2qw0SbEv87SEsw4mqwOeHK6FJoLg20bKQq3EbUTkBedTsTsMR
4qTlTO0X1vRTSspCW3Ukg5ipymFzj1A5WeNJpsSqU++qBgehrM6gTP//myqeamWnTtHByAA3EUWv
ZQXAbHe+LCKqOQ8TgWJRVGNSV0imcbO9MQvKKe1odKVdccExOCFzoP9/bgnPhbYUmgjrZyLkSIYu
KPRScv0eIqXqf4t9hubpFeeDnSiNLQ2P5ceilYEOY8KkP9y4b5ilJVMYDyRfcr8Yk0jYQqEZR0ZQ
q3em3zjPtdnhyRwQ+QDm1TT0wqw9PmyL4DlJQcs19D3Hx1Wn9UECE//IWngmRO9wml0IJ8nBVST4
1LDNSyB5Ww6eZ7jmPeOq4lU1soaoeP0/bttdc9pIBRKrBOZTyzhWOvSI7pNF39FpDtvcItB6CdIj
S3F60SgUf4PJ/6q//ZrgG9h/YXI7LPbFlIzBWH4VmLN0Q4nUbjV3sJrYp7m1Jf61BoJukdaPSZ2/
S4u6YI5+rgvkF79cSNfRSZ6hNOEzOVtCUaKA/cYgGwT97+PpSFLIH2STTW6UyQX3cqXRKtYgUMce
STRFxb78MToD3vAUKaJoheuZxxPm3EJnHj9RymtYT9BVRjHxoljAEIs3yXWbhz6Qc9jD9R9rGjvI
OmNZiT19+ZfqKBL4IbDGbeJ6H2Oa5UQeE+taQgzk8Ed6zG3x1Pq1wpbpRthLelssb4bLFyXDsTSz
f6ATfqVQX1U+jhtP+7Svpdtm2r6V84NN7eFfpCKeolfcSe7FTzwUoTvUJs3r07svLdgQ5RVRxS4b
dde203Rr5OPy1xLzz2hTtgOOFWnhHdXViQsxbJOIwy3YSjDBwCfW9MSEh/43OWHIV9sAMkI5qP7l
Jb66/aI2y8OB7aRTWUt+8pEAQM0POkuS4xjv3/1M3CD3udA3NPL7rN3i99/wsCYKBVHUYAlEYwfx
SH55U0CHeFJbG8VTwsAYqa/F714JtbnRe50DNYPGamFwCHHqmnCkNQSmVsRc9qk2u5OwPqItfwK8
4HwUOq69W+YvYsn+O1VlowAanhsf+aGWRfylWH4DxdXW8LFxG6OqCFLQTtoZfcjLq/gXQlyktNZf
OBE5PzfaH7KXD4A9v4JNdgolFQaN8DpxJ0l/RumSyLwy8tS+gbv5R13iD+de+OogUnx5VHWiAq9a
UCVIw9kHX9NEZdawLJON3U2SNUd68aMm0/0WtzYsgnh3uJ3wXYJWc0he3jc704IHo2J3TEVLJ5uj
Z1Cf9xqywjE10lYdRPPvL8S95bipFbCEq+WaCbVaQ0BTCNs74aotRJNCXyQITVvkYAwwyLD6mJ1N
1bty6p4S7/BLbceEXYFBNqt5PALiBuhq234+L10Gh0h46ZdlJYWWcCAoolbeQUvprbs0b7RffBMf
H842BSRRD2NqLcj8M4yiVwHZoHscZZb0W1M/gbP6+XQspabXVhJ6nbeVEmcfagxoeoyV1EpkifbS
o+Q/NJhSRMeOqXhpr3v0OAGQBxQaC3Z3cZJPQ+pyTu75GOMTlBiZa8VQY4GxBRdg/zS+m2U1urBp
fOOwQ5i9RQgbnKZHFmzpM4uJetuahm0PyX5H7VaTVQZ8yE0SYY4Bu4lYppzWMTBLDFeGv8RhavGJ
PCYqZ9132kpWcxaLJHwUKyXpEmMowDtohUmKbM3b3Mfx5kXG2KjdDY2SWx1kOiNG3Sl4Mg2YS2fu
+rHrQyAM6S3JVDp1IzHaOMAuOBYHxyLzQuh9L+tCVaISG4Ye8lzBHKrd1/wNNqjAnl3SFbw08p2p
9W5Zkj7prVh77vQ/iSgJLIhIh6mmIFb4CrGk92ZDNsLV+qBdRbfsdLeWp8z+mLGCJ3gw8q0+74Dm
D2KmCFK0sB0KkbRITgmmDtNJws79qo4s2D8o+LaExwWbzHhwg7OYnXEZijk8U5TcvCz32zZHVFdA
TD+2pk4JSiKiep9Jx3XcuMgJ/fPOR4TduITRcbJKnT0KPDRIjUYR6hIVIABt35g0yHy558mKIs6+
LYt2iyXiT5wPCCzaQot9Z+1bJIywDxqMX6tK9ILFX259n0+rsHOv19YfBmHgr5rPkXL+AghuFtGp
97CAqJNRaxIN9kqhsy9Ky1bDdoOZLtxOWgOfPEhjsp57mWAdT3LxOaPCt2p/Qxp4MAlfwYW8eE8F
juF6xvhJTe+oklKzJlUyixI0/Anf36GsymPdll/6rQ87cJIJXhXmstdL8ZCNN5TqDyume9xMhYXE
RbBP+k9ZDSz3R2skC7i737IALI2/djnstvOn1qkOnd46sCYYMEX4kMmrjb/Pb5hpqK/zf/FeVzcs
bdkwebeHNtQqXU5hKlirEAKDMiTWPHdAYIr93aW78GxKWolDDSiC2p1YOXIXirlBSuSuhrlyTvIB
JGak+RiIu42yW+mmCwN+DYQdGoL8PNzdWT1hKymavfAWc/JNA93RaZn2O5Yu58zdOwV/vUkb5hHD
NFtRU5YIn2+VMdua5dKvsDxV3XSDuaizWb3zF+vNjrcjNyyWb4V37OQprUXiJIAr4qaMqE7l/8YA
TCxXQ0S0Ammk1U5otQYOW8S72Tj0M4d3Z62DFQ6cjLsUs0+3Q0B+uCcO4O1j9LeCfSNsv3XcFKEJ
DmtrLCYl76G9xgdwy47Q9r4Q2hCJzbDJqAohJBek28XJHMjElZ5V6T0cgyB0QVc2XVKV6RkcScn8
8FwiolvaTKK1zeU5HFZL0Afn7wGE5EkUZMrG8zkzaJYOduPVaz/Ua9kQhbmVtUjN1nN4M8tVteeO
QTUT9XtgNtZNepjjaG+ZbsRZKB3DqRuFZ5bFz6IBxoZlOKRN5I7FFQ4eAn0oznbjbwiohbmRv6wn
sUAYnNswJSLTsFBRiCmuU/XdoKThnqHviJy3Mth6Fv9Oz8u7caRQsQj6ZEZr+DDfmSiUJxfg6Teh
oLxLfwhSBzCdvvel2WH9mgjkmOWIyJJ2OO/gxOcbpe5dlpj4VOV7Xym1grARyfAD8Z+cfAqZ16JZ
fKpeLpaxgTQonFfElkmUHoDp7kZQApR2ZPqN1xH1/I2b6i0i0CSl2L+kVdvcz9Y9UtpFRjjxWv9/
VEv/qyE6cxpkBZCc7IA/brqznAu62Swe2q7S74VMIpCi7w6fvPFugjGHKKmx2QkeLOYEr5JOYS0U
prIVJl7nmerBOnWI5mYN4r4DTt5fd56ENK7P9+dn0jvvqdNYEQ0bfFGpVHtsTuGlvYZUh50hDWYX
56QnMzl2r2G4SBAjqsI3wUPhESPmL3vzo5fjtq4B3GRBtz7FWY8JDbk+3Q/wwzTzwTagAZ56DoSC
yQwk7aJlTbxwXoOQ/H+Rt654xE64wQK5+r5P3/aZbzgJsxwtLbJ28BrHi0DoFgmEVthQiKhHZv17
meVJvFZW4sHdKxnO80tbRdHfc3Kdih/qYC8jIG2mImVPbPoWjvgSt3foWPQSYPEXtHRI3JRjK+Dq
V5/+UxbXjP8rRZfFJ7ELjviPRsc2c5njZ2mwk8Uo4dcq5A8vuzz0CxoHvc0P0QZ8Zf3xXDIbH+0w
77VplTbbZoLP93zRj8h13nqWjxeGR0Xl7CNeJUKIoynzpHMGI1EaAY+qf9o5u+9FHqtB7Bu89rWb
1OQFHEOBU2DgiHe6oWSYxdm+Z3zyyDmO9Aoa0otrfJFFwoKny6cPV7VPoFzOSDV1mgf2wMdSgCYX
UR38tW2sAySJYKEj+3YomecOiRRyuWCwS2kw+NqTAIXGNBRy7f7GrW3OyjZuyEZRwqf1vyj3RNvD
ACemRhUWyvSW09uKj1HQ2JKYFbA7R1OP1OVqqmZN72Xb/Fnlp+8aBgVWoJoSp0pMiA7UC9kmPDIo
HJaWd7DcRxB6SFtCOAp+ZH58dEwcsk06rHdvnL5tJUnSDU72U6FPSdYDyMDKpUgPp8DF2T4hEAFl
PrkFPLRHvy8INb6RLioCrxwiqd0thXCDJYBfv3AY++yplLfagfDaOd/q1SEp2Oue66VcpqJCJPrf
moSOZCnlNQbIuVl1u/NpSxGQIrLT8/NPjPcbHoEMP+l0ibNf+OICnUzGNejzb5RY1BK0tdwArACs
S5du3rvgkD1WXg97QuQOATMP/yO4nxxKrdv3ddc03lzvJ6UPU7v4wG/X92fvbD3L/2dt0EWn2VA9
JPY8/2nu3EPTKGHYC7h2j1OIS7ZfnYP7uYIiONtvSiYF2feoGXPTmUv+c7l6fzpmGKWylrgrgokC
rN96m6kQdiG+fNQDET/r22/bxH7lOQewigfMYM4sTkDkbUIaP5MNtvZjdErZCgI+bz3OxRNxT/U1
3sqG6zQjfJXOksMdqf72m9x1LMHaxYaOk7mjtwU3tQtmrrkIHqH144CNedM2qobDOTELI+VWixzj
VqRcNzSHBDRFSGk1vEKVT1pKAI3UUX04muxKINRHUpYVQ1eW+Oa/GqWJHGlPy/fKl0rQ2XAEB//n
eDFjVRezXeWo2cF9WTcfhI+m5IBTU8OfTMPJ0434IBFlayeJ4rLZGEpd/cQplpHo+S2irPhRQMS2
6tGmBbzFsrajUH/zKSh5XYZiL0DFHv+D6o8F5PvL6dpLBOD+/tmgMU42JX0zeKSRk49eFWOP+DPf
bkYOXimSebHbclLtw4Jz1rF71OX77olkJmdPzvopWrnaXakmFSb7DTETBcBJhIEeh/INnv3nJ38T
VnWrNdoOtZWwehiN4TNZkcLYSGBApogB3DYf6toOI0kdAyb+BChkGW+d8SfDEjZB32j3UGoa3dvv
IZbVCk7zppk4fx0OoQSuVFE/L/n6HDf+pMhE3FyEQV97b+iuGtj7jsFJqTd4EiPGgHwjxRnZjEUQ
Yvvm06IaDwafPjqCKxmV0IEWOatrcTvAxY1IEBJA7uyHgR8SSveOmU52lPUH09rhHrZB7gJirpmj
Yrsic2SIT6oVzypYXLumFiV5mKm14K0izwddgfTgLooOgRMdfduiphMky/EleUH+/1KhEjCIOXMp
CHjgcIU+TpS6fPX7rJMPs0goMy2aXihDOUIsIBSqu42PH4PKveuIzrMdw+kSRRQZ7oNieHfuH5i9
NxR1DnWJ+CziraK9mtCQc71lx9ZSyM9A0IT6tYCntk7Ac44dxH4BGehPx/PklutF0F7V8pW+UipS
onvjxVxz1Hkqtag64wF2EJ75S+OiigKUFC+rHB7hkeBiBAAiO2FiaAlRuBjI6LgD/tKfsHIzGJNu
AcWWPdn+r26TI165TtHGRgfwvO30ODKctXSyFggXUTZIqt3PvDwBhdA1U1uyXkwtgZHsHLlRnrOS
5okNfig8Mu6TI7Mc6BlSVXR2rX41rDjoTfYjDKHn2avd8F89wQS8yxFjfDBacQ9swSlQhdiHjUiQ
1zBh2qxIJ20Hnt4hXwoOuAKFgivMZ+Jrpi/kJQSFP3tSYpMYl4l9naD2t8E+3/7kGzjiYG+We3Am
nNqR8lX3lhfHS7Wzqi0PYyBVdNnABXC5bhAPQlOSbPrn4xcnVPi8dvtWZuV5Kzs03UITcocHJmUg
KRVqhf/iToDvlgLbvbn/NzieoJxCVvS6SElUvYuGtJ8esm1aIEeBUM54ytsgm9Aseco6lnMF2Mw4
tyxohXMmP+ozJrKDO67IS5WcdvehzdUQblosKNrSZ61nnk96aLTJa/J/6tsk7Ou+yVYIEIKKipNZ
Fp/CcRSNPvFgo/RMh+oTurs5Aa8Eam5uY+gMQxRxUk5NMdwZmHoRdp4RDHAE0jAA/+7m3rxB4ak3
gKFxLLE1ZZv4RH1Uj2U5hzfXQkkoPeR1G1zab+niEMur+M+TwQS3bovDd765ytLg4JQCJ8SbCtOU
w4aQnw+xF1Vb+MJ/YNGIzslGcemAbcvIlZoTtR7EQi7/7G39ExyokZ00uvI1Vhfuf9DD6RSFSfYc
/ilAwABYou4QNbp2I/PmUaPZYAzk5wOAP/Zs/ut/21ymtzRbB06PIJdSNWFP4sQ8iobMl+b3xJGd
aEJawBlmMT+s9Nz2iKZlzwaluxNYNS2kkfHje2zMDIpxuhfahSR4mSCabgbvdlK30bjxWnWN5LJz
5aXXokOS6/LfV0IjchX+ExDM2O5LyhRKm/mioUyl7mYfKRVe/Wd2Apa5PeFe3AY/cy4yZODM1E7m
V51rQ6Rd8F/u1eRbAyoj3jm3JKAT9o+NqxHSlHAG3mDZAIAtRvnVLXFBcnto328yXtd5h2doC9SV
L06DI/9t3I3SO4A8Er8/891Htu6WghJOai1Fcc33LbXxjfTIAeqwV8wSMdCFVgTwHC3wW+GKGliw
n7luS6DrKO1EVJNFHSwhQx1IU812UdUGYlEKya3zJLuzTunJ5V0zEFJHX/TPhqPBmGW9IoVu5csk
f4dQicSrXY6R9C7bENM6PJlYkO4/UsucJa8yALDdzeyR2tpvoSi4Dvx50X3eE1pVBbOqIiP9gewi
1pN738ezMU+nalg+FSfhsar9f7aFYm2VG1JDmlWNa86/80aPr+MNOP7wGurSOYcUlFfTmA1QTulC
LAS73TBgJ6iZTQqIli/fHmPe1YXaih0ZyqY4xbggJqmlzBouDadJH0tLLeMD8N1KxvOmYT8EphrO
TJRx++9p803M5fyzX3QxjkhWeOam24dIMfB6uL2EHtDA2it6ZCc7YX/WoS+OMq7t8hBtiRv9TxIe
hoe/hTijoysWPucEZ8uVojoqLGxNCimpWJREPhsLenwXTWCA3pXgkS7Sy8ElyXKtRzOfaWp55rt8
fcTNe0RBLMGSVQL2dWPwD8o+kAShQuvQKPecEqoM5KttOdyayjQgm9A//vqq/SxFW8sRsGf6qGR0
PrR5dvhru1oXFGzo/vpf0Jq9NezU/mhUPdYnKrWxQwuVzFou4qrnf/3VYSnMjIVt4wRxnp4oCi8u
jhaDyqBehuxNbdPFuMDo2RFtFnpPr8OTkKOmMLBIAYRkxuUv9fVNQNeAQoqhATutWg3GeaspSt52
oKLxMuDsVB19VxVnCedpSJI/zlFSAoP2EVsBFGogNz/Lj0BYilVm9TVuSyF0g1w6gdXrChkad91r
/rYnQ/OTRkhSnHq9C7Otb71dn/tdtTA3D/gkl0pvBOK0o6WtfxOIQmL+aePUkIzOhrSO8TbrymXK
q7YxVwjvZYfWnXjeaFVEbzntoAcQI7330wMfn6rmiNRweSl4s7h3JrBE+imBkD9WaBVnQha80qoE
+YAGvQMO1cqOR5m4dfURqZKPxtvKV1AnCNI/ZN+LKiqZcYFF2BOKu8+3B96HWbcEfdUsOVPEHrkd
rhssT3/TrgzIf84qqEn4Jljcyb4gFQRFxSMAeudCsFKkfvHz6WM5AcsIo+PCBNTQ1qW3jFwLwG1B
8FSRU3vgz2PVT+Vda5NQDjkOcChfrtWFgzwltGFp5neunz0QFdmzE3MRlWmTwiuDuyaB+I8ab7ok
f5UuJKM/3QHaA7EyTf42zMJ29wYkr93ZTi2OrBPSwxFuRFRA0xoYs1GJviFGWgaYyIR5SqGnYTru
NIBOh/ZZikDqw1bHt9rni1afSh20Njw0orG1f6iaL0ZdAyOiq3/n346WxfX5IzS4kLAEH5TGHbdT
2A1wNbQMxgkCwUmJi2KdoNMNusPvEbR/FUK4buUROD5IC+waE2/id3ZqKyUUOXdS7XZo2stN4uNo
raflSrqYnGgxBU+MlfRfrxeek/E3DTMpLyFnE/GlVfOa+JdqWdQjcrxIoE2T4Q4C2o41KvqVjM71
MwhcV/ct7TsiMMdGfbzbtA1hJwNT0XFEmTMwxiD4f0n4DfYoQSw8miaqzzvJGRbW/UTYFUq4oWVr
AdS+qVi+PiwtnxRoqCAJUEJwm6XMsAqCl3yO959yAp1YSuF2B9m54UoGoN6Fh2dufSELdbHhADqq
A1z+J7dEwO+1CAUgQe7bHKU8ws3aAb0l7XRwb+vKvMVG4TFVV1tChQTnlS6pfmHa/W99wHGkGlnA
FzOjPWqjsxLQvrDzMfiPAoq/Oj2FLvewxfkzCVHC18ufsXFUfnrLSQaus3hvxc0gBS2aIPE0mSwF
hOOjF+5XRbMJruZH70e2ey84zV2XfZpVBcYR6pHajuJGB6vhQIBxhWn9hV7WuDM0IuFHfVV6Xjww
ZLth7+I9RFoiiVox5Kx7KtY/8q70e+hg6yzM7Kt0zDKRpRodsoVZUnUUAMrYp1LfmxgaZhL1CR27
WZD0R14q3tv7lAh0KE7m5oBJdMmPYClsOUNui1zBpCYnWYadzu82mxrP9/U7/eo5J/XORyNUUUaG
4v5o3uj3Kuxia3ZZfsdwJDMgssumb+/wFsTw2fF6wPiysfF26IRQ9+E79/rOJTxlymxYe30yd6Tf
TEJa0RXfrKSJYP+91kiYBzoUTUgJvm9VW2aew/HI9MJIyHJwC9VOiG/fQ0+voLK3RTL5t47506LD
uhEYakFajTmf537Tb7z5589wxUWM8Qcpy9N83CAe2MVNJFzTG7jGi9bJ6gBlkMsZeq35d8yvL14W
DBwXCmZmA5yLcVHbs6fKmGL48SesuMyq+eCczF90+A7OhFSaOxz4g9HEQX9fQUCvwOtnhMHM9Z14
bKxlAwK77+4znOBdcCP2OZHQxj79xfANYwu7b0q+xCED/1Acs3WD7Rmuy9odIJn2rCTr+2hiso4d
3r/IzpsQnuzqVRetae8T8D1jRgdPdm89EUgxoRTeKytSDD+635vw9ChloZfo+s9zKuRn/0wMvIlo
BGXNTBwNnpQ5/95eOY+l+mh1nJS9iXPgKFN70SNPADxML7KgNU4bgqPPWA4SwQvMIRqymGj16sz1
mLSrpokBkpQGNrcRvCGbwjfWPgiDtubVbDBG/Bsyxwi3B7c9VGpWGf4m++paKtV6outmnkdA8+KZ
DQN3gD4gDk9ks7PN4Pi2h4e/EVxay9qXgrOysqC+NDNlY9u1zk6cFZEJ4t5wxk+P7mHkf4AeimWB
+nmF2XP/VgYp6Ov6O0iAEw6IbRotbiXo203vx7BXAJxIJm7DkbVXvACZro9RLEU2KBmheCyUhXtp
9ow2DjzzLWE81aBF/sIEHhs605QkqQ6ijmIradbL8nOIbE6hjt8M2BFPl7b0ShcFQ2enKSC0PR4d
XYq1vtZOwhmpVPPAwzVHc7ZfwdU8BDzwbkTMMsjSUhfhEtAXj+E5n3Ws2cpZ0fc/3M2LDyha5G/5
dnIDtgRkzmX7v0e5xVd7Ds+UtEk7mix9T8n3Sh9WRmKnuPmTQ5ko47NZ0huhoittTDTyaE+T+HPm
gxbmAmV20LaRPWEde6PcDl3wMzd32WFmduh4lUQIcE/hXZQKy2QUPRuMjM6jK94s10HIUXdoqeT7
srPYRZzj1FWvjPCaqmabwgTUJummYRL0CoftI6lvkEs5T0YyCI2wwZm8X6TKDk70wrQJ0JwWQMqo
68ouqFzPXbYJh9fwHtFbvfqvb0q/U6dytkik5GRaRvSOe4slCr4sYqRx2HFSQpPLxIObhxymRbed
rNgVUxqwK5PTZK3jly2mOxk5o3jYz6zalUuEoe71TBW50UPtn9YrYPoi7bGWqAf3Iewsg/aKT3OJ
e6Z7pjzWp/NjdXHjRpXJBWZb2cbaFprh02jGYUB+GSzaQm0KCVursW33AgCD/cVVueWn3F8kL/3a
MOoiv2oKoLkVglW1UFpBBQ6x2elfZHPHT6jlny7J6bt8a1yixHaC+uCVz5sUzRTKGH95tZFhrW+B
MxBO35l0vqklzp5w9P5azHZvUPM3p6oG1IXNkZfh/TdqpOkoCBGcm28j1fGgtBO9k+ZQM4DsnyLX
r3HSRc/nUIjmQ1A56vxYBqLox0deqj5ULOXDKRejgXVYZnUzJYSxDVr8OJB2CJs28vtczjPCubTC
PQ8bkyc47RP+T932IGMn0lxWlfKZKGc0LAXaz1r0A3uHouBeMVawKivIylVB4dY8awgG4Pb4WuDG
itSRPzMMq5H0INFfYI8q2aKkhRTH2V7UScaqXiyUOZg14uefPkVab1SoHnWKEvxBC5goOfNjrsLt
DgmUbNyq/1ZxCJL0Ep7TASMIRybIMzAZ7LIPDpt8XtQ7FPB6hCmKbigActATS2Uy6iXkjuLyehzd
XJ1YA9hiGgQx5ZJsL2YB2ekF3TJxBuIo9lZP6xt7mgKBS6kLm+RSqOhPHZhQRZUqMb/3rSOXVxx+
DNPHxPXDI+Z+h8aKQ30IriitVUADK5txMiWf6Qi3l8CCt/vs87FMQNxvCxw9CPVNz3pHQ+5aL5C2
wCr3iiF8zZlin/iWebkbxBdusVBo4zGRV/3Cv4CZRkXzrhh++WTlqCTlg5ZWht0bSKKCRxROHDc1
3cDzf2f41Y5FoXo8mXQsThPCEytNsssr1xKY4U9FIaAZj9MFnP5aR1wBogxHBmeNLeFErr1Pw//K
Ce4pQQUGDxeNxndALgqPBTJ0ENAA4ILdQBDtkgMnLr0QbsYquDZBYpla75ghnuOXSPx/UpUKJgsl
DIOeJp4j05q/rtAucYyCWH11H5K4E3CnjJKr07pAve50+BZCEpfeFH5262Sv0gwBcaq10svLtyGO
JEXa/PRt+17Zj6DLJl/0vYeqg7jrBZKywxZja0C1ZrRPxly5GVhZxW7t19ZQR5qmk9myhRcaeNLR
jI04uEPqq0lH/LySuPbgc+0JIrHrKfSJghfJK+AhMFFjdBh1ESMKIo/t0wa7ox7+k2bHV+XjOYSz
JyEvPe4vJm0UoR6E+nzRpSJ+jGj4zPnHBQJrKyvTW8jYIGIjO5tsZT0kY/Ab9JjZHpO64XjMNgdT
zohX1e5fJwY2heC3JcymXFRStp0wcGkuFEAXA5kb5wahYd6mE7BfgQCj0DBPj/Y0I0zj0n8A4GfG
mxFsemE8nth3AWnW7UrOtlBAbc1/0wfCcD8zML9P54JMSRA8jZyNh0Y9eRF+ZXShLfd1RbDw3Ahe
9CnmG5GBcFDd/CwOYgsvN6jk3LV6MuIMuJf44APCGSGP1cbMWQi+dVklAjSXkFqQ5V22mfbEj2Ym
TR56Ms0jPNdsODrOQV8YBX3PFqwvLroIwRB+OvbnHezVEju7MAcZlugn17DQUKz3aq52mHaVGKeY
/x0ENGzwqCgbTJkV0ZC+5Ad95dtGdtDsnjNBxgRH78IAiSu18pH8q2cx0lEvLZgiwOuOepkAa95D
kFsAP20tl3TBjyCEVpt3aEI3UmRfF/7vxt8AESRDLOm0i1yCTFDbh0fVaKnjDC2z/VKUd7TbWQgW
e+nebIyVUe/0mCjhhkWhP1Wjewi2FoCJIhnaAuBKkaFdB1ojjNKux6hCYR/zXAM+DMLE1i7DA3P8
exu4nQI8glIhO7yRxcR4N914P+Em2Jh0kbUWcWmGRD4i+uGl+U8hdWR49q+/YJo5rI005r3UaMOb
TFBRkwCSSoGcg5XqpoUfgtmO8qyBfPErpTcc957mnEmNRY1SXJ7C5gTZL+6Vy8X27zLXg6jZLOnS
/Lrc1d7FAtq0/M+M7b3iZOH7J3e4vyBWOBxab3GPhwyKclZ0PLKDOV3VXXrZq/AtqiSmeXOHlIv8
vHkCgXa/xeXPBTZi8jXAEiQ6+8/5FISeP6p8crDsbAsQiKTLCeprKe4iQrs+wsbDtqiuvQY55pRl
iryKBGJsi5AqM7czXysSUp1S6yr101uMhYAQkLrg3Hv+JW7KQRMdm3TDt/nbuzp8H1J1SG/atpEp
NIY8BGFSNCiMCNe0SLwXrOHN6ksqzGoLCoKK8t2xmYs6BKJtBxFPwChtaPC0lMzGReaoPRAjQI5i
n2uWap9rb7whugI0ga8IkxgkJpsoQPpHTv/GS2o0o7LFZaC3BvGtfVWzTouZUZRs3TG4rPtHzbrA
qoahduqMGjIGYByhh3xr2+scRLbK3MBcWhD62GZVJ90fkRghUj4cECyHNBt+O9TG6ggwYM2nqxff
c/lWYp5/m3XXNWuH8zyO4y+bKJU1/fcaV6z5/vc0aPPwcVrahVFN5+0egxlpdevx6GTKG6iGPDPa
pjauqc9N2KzeSyfR5WQbjOQfL4TjryO3y6l7TP76Ie8OCqTR4lPRFBHGRc2V12d0JR651W21BhpY
50rjjkG1yhmfcVYgMqByST2dzebePmSh9YiJhETf0ZOtgTAXHboF39hiQ7r7pnQ/9K9aTAlatmlN
RYiLzYqMcqS9ugr2L1Y7OCHR4IrJEefBjEU4aL4uroDUwggt+wR8XUDtalcut0TKt4DF4KXk9xt0
eWyAjp27A3BiFCtM0yyWSe6L75qgDYr7nZ0UpZZeYvdinYarKoVYtMKRQfzLZ/ajvVgEpLpn1lwJ
NQELESvaAPsGZzIveI6ySCDlGNLr6g5wqTq9rfM6czkBowsBJCQXKPJrqid91RFWLWGQ3QncbFZ2
USkv8ndDEcxZ9yoiB535gwr/Joq+K5PoULnmrCnSteVbvzLMQXjqi8zU4APGSdLlJrFBREL4SGr5
flkFd6Ldtcm6Cg8okAOPLEghFQHhF7DAEPJQu5xBBjFSExfkP3vYeBTrJV+NC7WkhEoiFgSe4ps4
b2IjUDA1sjsFvDWEYRJmxRP9Ns6dBWB+l84wDCs8ZlgOmXUFodqIC+i7cSTACdcXQ4O/TjIr5N9W
mzBjkmyKGUpXEm56vDVH1RvxF24Y2hpEQTMcWMCIKLziprLoWIvZ1TE9D/9Hs2YkMqYso7q04FmD
/z80c4YMYEQssGUFUN/pdS+QR/e0bvCnmr4UdPSaKAb2e1rGMPaAY/72sEeGVS5jNCzf67ATN6AR
PtqxcUhxQdxYhV8FH25hZ20dj8lPMNsJtF25voZWsv2Vaq9TWT4MyfNRCUsgmJ2dsmLM9EU+KBsY
TrFJLwCrMbeo/AG3Q9GUfPpdhOdbi5zQ1JnQlnpIytpc7kpmxzjMdiyhwlIaHlBd53n+Tnrm96ba
krOqDbmQlp8R+oLjjv5LoEu8iXjNYgXWiw/quarV5uvw3WS27UPXqJUVO4ko2Ix27DI0A8ShKUaO
nsF+rVG0yV1aRJOhEA/RiCMzEfTryXmuKv/IihnhKytC/6uKxdhShvL4leOoLhN0BBJ6Szhpp8DP
KlhXB0AuSOeqDo6GayLt0arvv53uW9CAAtIlg+NPR1djF112vXHgooNTchmtMKFHYV9q1gCIs9rV
WeP+EV3NWDlFKk1bRcuoslj5+4cq6HsysMy0+Pff0FhKNL39eSDSHS4W3esGhG8+K2BKwezgKMgC
m90LCSMrM9jnnZ4etqiqz0cp+nncsD0+KLb9gumMKChJTrMxAi9zEsnV0jisPOyrcQ5COfP4OM1f
Ls48LgDGQFnU4CJsaEuthRT1jpB0Vaf3mzU0jOKghC2s1a7rrmjN+EpdgJtQldt5E6IIDdDY2Btk
r5kY38I/Bo59NhbwdHoNx+SjnpyDw04vGy0GFf3grcW8ZK2EHAXXHLamNhKmoaKyurV7Kwhr3Am9
ui3c+dOEJgnt7Eb1qevXeG+yjEy5hCZmmIGRfvZQJQZ/yZqIBRODT7gzEqquc0FeI6Mqe2/HH/0n
KybV5+dswRU6sVFd3gYPiYmmDJ/w5u444F2iiGEeqZPnC2C59/85z0DJLYw+JliiS8yCKsnSFEVM
IjNHOmvT+ez7UG4o2CiqcDgdxk+omzJDXSTNWFzsYsIxY4l/p/vsxtPt67R3xfllaLu+i9+166xd
x/U9zlNibxxKcb/GZG4yrieZEeh5IHGMrvWMzqSktQST/GJ1PQ9rU462oq7eAivzQLb3jbeSuCHL
fcfmr/CXF3BUenXk/Vt2s9ohEXnyD+cw2p7hOWW63p2xitzOi9+rVKLpubDF9xPLisEqnAkBoWwA
2HakVtErlPN3dcMi/1UyEA/4ntFQbCZtR9P8J2sOsDnAE4DM66/g8W1OTK9UdywP9UPTiBeDgdpN
I2n3RC4ygC3AWHrJ9+vM/FNo10mPynxIsYxmQ195laIgGPvmQJx73FgTguBj6nCr64bcaDe0TnSd
xSGWEnfJPCy2Q1NBqH82rYEvoq2wOsclws/myYLHf9sRLTS8LnWU5DSqVB+Yce6hSJDgCBvju0kw
ndlknKieSrErPuyRnZyr6GWhBa3SIEv45mTp5ynsfCbPklQGAm3v90ueftO2vAewHTuR3IHnaNT8
gxsjyuEVM+M6dGBZiojeQG5gx5txS7cC05X5mR5YBFhrim2B5kB8hofPgYNMaU+GAu7WxdlRUEQ6
NFtudxwZNOonXDY/3flJgCKF+kMSEAXeIWgnvd8b7qIO6HOm/koJ2Y6DMZQOKhzxfX3gm3PjJimo
WBOSblYs4Pmdsnzdhz2texypaXakupFMAUkLZPkRTqALzeS725fqcIJ0PaHDCOSewQrbiGqwcVGU
v/7DIjbT8FdksDvg7jagy7XXmaat65JxhkSz4GcL2OUKTiFlvN4cNemseLYoZaMuZYg7tj71m5Eo
ZE5cNWFPGhbPnu81vOlswGsgxIOdGaFw42tqIHkyNkpln0Ttgc4DnBG+UX5SXq8L6mXLbuxKMDkA
zPXsFQ9dJFXjrN66dcMuRdomX66rEcu+Oj/AnDytrIBQ8kbLr3P09CoEXMDPukxYNMcXfeJjj7sN
RXdVnCRPpPfjIfCmgxlJgKcEKPr61IFhDtnxPquoth6Wcfe5zgPZ7iIkH2XciJBxM6Ag39QauDEw
l1mKP2oXcW6wAGaKUzKitXccQirsVkRhne9KEXPyKfiZxugWiZZwaYWukpXVyy6qyQf/JHVyhUpO
lAeWiGl3M1Y1tpPiiFH2gosa2rkoysYpA1cLoysci7yRwJorZKilCax+Oc/LAEQC6/eZLokH2f6z
E9HwvlsHXA5HPiyYQHvNLvW0EERysehvAj+C/tglU71k5KP288FYtF2fqLUnkhS9TsiQxRyRZMKx
zlyzmbeRnfd1st3+zQesPYDroPwPzzAZR0BEUd+lx4s5xvxpNZ4z1rrFIpTt2/3ceT/AfF9LcU5T
p90jYju+kguMMgrr4U/fINieG9aJsiuL5CWVYaUVe2p5DUkHJ06p1QmVzoyNEM2XHb2tru9QtNgj
ldmBrIrt4b99Ly/3oeiWFbhtR10woRK2zcChPYrhIuC5C5oORA7oBaIsl45MJ5nQMYxR4YSs6s3N
tTVyFphQCDOwiniFhF6DrR+7nz8I8Q26qFzu9PuMzDOywTLZjP/a+wTYXay1QXpXm/ifE8oosavi
hq4TroyixkCMbxCqcUa7kcX9sDUNu/92BpI+eqxNHe+btNOmuyh+mnRFfE+Nq2p3A5cUctm33tjA
0TAovSvHF3I5ydL9SzeP8cNstVtb8qzkgMZP8rICCYnIVL68iFAnlYdrOrMQESxp5J9xDoM9PP17
BzjsM+z9hg4Ivfw2sGMF5kg4ckRE4HDPGCT+QAum4iwxHm1vuvX79FagkcHHuiqW4w7JJaeoZ1sj
7f1XZrGWdwxiBNxvuOgNFLHyRhi1OU1/XlIDKcHeCC74JojYDnvk3o4dSt27X8NgZG5bES1cF4XP
5+uGaexqnRsBPJrpBtHJxJUaaYW/1UYJ+xn0G0207fSXX6lhDv755uLrhRZqOzuKS8BAZtoQ75PH
V7PmdACzbGuGHgtZJP++viUcvmlb+Pb9HfR6ockVnkkwdRPTqbmT2w76sR6tN2qUPC4M6IUwSJ77
enXrW8qZqVD1NdID3GPnIDbtdCeWIS+RPqHWeT56y+40//8s9skbbL4OzEYueVyyWVPXXKReH8xc
BPAG8Z2QlVejrlq+UT8M4z7iiyquEmvFx69TbbXtb79KIYtl7wFBcB1psSL9pXQr07p5k2LrvYFw
Yk+dObI2eYytSzlZ4Gy2nKkOYqjNSp4By5lGfIP1Uj8dTIliwrbDUJB+6ogP1vnSdpCUe30uAxcS
/DiCQPECISTFTF9HNQLqUhBzTn9LjxKqr0gY9kOjlgfD9DqUo0VK2q0P4gB8TRTxJ67tmnIqhRg8
JXubTOboM+P8rLPCIzBncVySdfbfq9sDkg+s1jO0Bj7JQdNqMdYPZzvDk1BYSrxF/nbm8kf4XNSh
D+kUIcEtjfHKCwIBBsbHOB5v3c1NNPqGycAvHYXgIxesIODFd9OYzrs6YEiqoWwzwJAKM0Yr2+yl
1zMfy3JT3LP1j4pDzqHlnsX4wYctDUUi+GFbNunYVyCueMZ62OSJKSc/tgKULY0Fvg4xMZcNsR74
4/0S1PcczyH/7g7mZFmMUMVfetQuslZo3NDwQwUNXmAOp2JprrLIWPlvcLYuAhG+82KRFq5VbULH
iCvBl2z24l3tBlkJs9OUJW4lixNaXFx28FEXSB70wh1zw9Dt5RoQ+Oj949FCwn71CUpFxiDWsPO7
1WVfEZM4WxFbZdYoBsUz5OAjXmL3JaE8QsjXOx1fW1yy5T+3QKrW36pFwp7UycgyI96P83F1KL8V
eccGR7pmaie3NVRbYIdwlkycMrL+wWvS/YJ7yzpeLx8x+fbnw7KtrFoTRaTR6xObbEC25QWjhUnQ
+qDCL+QXrma769+U1M6TXZvwNY78BxbtcCwHYIGGvXQXnLhBJvL2CHp7TDIau1us2Wnny54VKJkn
U/2sIN7Se4ARyhnVwHLnFUZdCF8t2Cz6wPF0hP5YE2P1B54YUCKuBeaAso8vSt1d4ZJ2xjNirSPQ
+DJEIaBy2VDeeVqJKJVs1LKHkNTJP/Ejdm4eOgNZCyS9HZxQ7OyctWfUY0SvTLpF7bUhKVOtfWz4
ZNQAE1Gvhd97/KpcES2mS17s2LNPGfQiqT/+9tMqv40UpHVJNGK1KhYwr41B8RC3j0npqJlmhl4t
4jKFQDWm26IJL/I70Xi3B+GFXH9Pg63Kfs8DCs1IjBjoDji1RS7raelkFBtqRLfZcVcLvtcSHP5B
4TiQhTd83x3aMwBhzvHPqiPQvwSyRSEvlv+n3/u43CkNlZEXY3T+yrxhjkigogqv5l4Yp89sZ/Qf
GkgiLcPMsF4El5dx7/pCsXRKwx4b902R5Vi5pQdVLgpLlGPV6hNFu96FnazokEgs5ekYS62MgNjl
wi2A4+U4lwb6rqvsVTWMnW5d31ifxI96QhoxGR7ald62mJ6X5kH/RxkChfKCIkLODSfkjLzB4vXY
DkxDAJDat/K7GcCxI2BOR6etP4O/Qq9/YAbP4GyuUbrFEJkil34RizOmAtGfLA+SSe46+DjQEEXN
a89FwC8t2Ng5m0FrALuRJZsG3iXaeTqOFYi5q+kDxx6UCcnYC/1bUb9bTo7DNb3tgENyXdkczF6n
coV+Zzcms2JCccZ8yIQz4SSWCwU3y6pPGfdCGKaDSnhgM/cVDBebnLa0zD/tdhI2JDi0UA9j3C7l
HugD3GG7ANHj0WRq95Mzbz9m42r6tr6LJb42r4We++TbPAkqEwExo5JoGj54Gt/KBCWymBXTfMgA
aI4VwQPLSv8DP2+1at3miuFoffCs47jH4oPBV1BMyO1HpYEJNCysm7ByWGIjky2Pjdc5Iq/A9st6
3M0Gi93GIYXRR658Sriya8/D2vU8UDeHAr1aZnQAJeE/WpikaVUFBuMzD+pa/uVcWpkXj9/dYavn
goCtdIZAgfTR7npsZZ/zwwzg3xVMhpFqxaE/1J2yq9upqFc4rEYQgQ0QyYIyhgTP/lrWVqnPIxcW
aSNWBjdgYQc8DQzwC4C7Ws9mZa9Ks/JOxvmRKDhbXjHnom4eirtVpTaL7WocPa+oDe6etzII0/4O
HQENzqpuTol9a4t3LIc7CEx75JUA0jYqvf32rAHH0cdLXb8FG2eyWFGI/8SMJI5uyASLhtajWSiQ
wF6TV28N4iPV0uowllR7YxH2o5Ak8XtJvD3uuQOELOFj38XQlnSmjlP3M7jtUpuIvH3miAQoXOA8
hhXyBdb8GzZba5GxByDGn9AXwH7VKx1lYryrp75z1YWLsBdLY2p3gDfvbkbELFTKFzazpQ9aqC2t
jNHc9IFUlz87+37/HTYRIeH9bS0qwIknmO+ByGMSsAY6WBs23xec4e96/BSuotOBVdUsoVkDWLem
1CJnx2zk6MijX+P27hwgyFXXro2E3E9TvbF3i+L435tHqg8ujfIXPPvt3HEwqu2tP8c9V/49x1d9
k/8qoIC3BYsrft/QqrMQdcHi0/5JNU9W/GGFlS/781M54tHIARVCu/Zk18Pj1ldTWSpiAc6JUBMu
UgoByHYsl/xu20BSbKUi1kJz/BASb2jUg+zKkcPRPqlp6g/RTvTI0mr4+HfEUpH6gh3lr2hVMF07
wwJkavxN+ecYzVNNcJXX8w7StCWN2mIj/5kh3X5utpyaqivQHB8+157cwnWwHJ/4DiUYaY0j05xR
GVVdqb6Gl6Z9zpgWXjh9hPyfgMj/oyqKBrSE+GaWbXdYlTlxQmaq/XizoWUA9sKbR0RGMWjq72LP
N2aQYzlP1K8+64V/8aIZwkRdvYAybxdv+ubuH8ZtPHh8pXMjVB8bfkT8MlH0v+En0sBp+Dd0sJd+
6Ul/eYGoGiggKY4V3Q+wnF8KJl3TlXRc1kLaMwwjuxLm3QXZxnVhPZbigvV+sO1Lqw/ibmuFPA3U
HlVAt16cg1AZypRH/VKbO/vG8IgL+eq0wUirjDt+j8HKUTT4CpwDu0dGNkPTBspDyc+ZHcJ2OWgo
LG4Xr2KnnKbv7/2V66VQWF4z6BreqHa5yeGAle/1XZFUnrH2sFHumAVszBJ0cro3aafcrpspAhCY
lVI3hsK+1+Q/n3ChM5x1pLuIKYanehujNAZ8m0vwGiXaOv25vcdBZoJH3z3z0SUPv6aW8uOXBe4i
KFLsQ+SCAP1dv1aIsM6HpP5IQ7xA0BFIRivOh2oS8J5RkfRU/AzzJyCskhI+nTIawgN94qG+8lKW
LqkSm9mUSZKM4eFb3HuyDnxMxyn03c4kzp0X8QjUz1Yye/7t3bB8gHL8LY+fZyIEanGY6LaEl/VI
dqPv5OILs5GXSzAb76O6kyPyYyvnEdROyxiixNUz8rZYEQOVSjpPXj+HIpyoDa+XDPOmXHbQVUPp
KF1aUmREGUAQdFwjgilns4PHiQ4Yd3Zf3Di70yX9vcHrIymGVp1ecdavxBuWUU4sjxv5qQrbJySz
EieHw/JBVu+YI15gpmoL1tw8qcd8oxQ8Be9b7IXXqmnBjQDYQqRIpgIZeNGCse6l3dRGsmOLBuvG
vM1xn/9etnXa/WGcFEFIWxYZvwaZYE7sfSZT3ZgTxDkWtrHqxErOlAw0Tn4dbw2fml9Hq6xLJk6O
wMFeQwWAKXJf5JyhdKHEJOj0xBRk2fDi/RBGy0gB+rt9Stl7GVpOWf5H46FOZjrH1bB70qNwLha5
bsDSurVIL7ncKsuXHHtxuJrSfortrKXjfXMwGXY0B8dQNOAdhRAeTxnynXvp84RRHGGG1q/cq3ef
9KZSlYHLeWCfjN6zPEAOUCbKSk5OopHHduAQjhjKktKIJd+Tc72frWwI3gn7/myoCdHqRmP+4Ybl
s1c4FTq+XI4ra4499mc018w7OA0OcbzJdat6sCA1bleJ83aJckvnxeE7HKqq+mO588GnLqmzMpm6
xDht1ocKgGJu9XdDtcolVOWRVJU42pem1HbxgP1y+sF0aahGaCNzMvEwlpG+urDMwxzPvmCuza2R
slAMwYwFmn6EW2otS0F9E609mLlfIH2nuxcGWK0ThfbboIHeuMvLskLyJW9IuwggI0nVgIWWfSoc
BLrxbkcCaXJhOQ0GzhFaYyBn4irIlTV0q8ltBJT7Obfq9mRoRSIEHFnzmlKHdASRxDB12iaW1zs9
eMOoct1zJPJtqUql85ELWQNWl6T1CP++i9u6fCDYon49MtCr4Uv6y93WDWSVv93GK8WvBabTxqaB
omJBPPXD5PW4ebKVHapoYjzRXkrfZpNz4hltQQGZlef2T8F+g1UnkTJhkpiAy0EB3hgGClQ1ZNNE
DiiHwJo/KVe0EFJgZDSNY+TcfFTTejKP4kNQR2AO/ZBnWqOO+uYbfpamXLy5nsi9zqqjzlJGRv76
agP8NjiMwvxXivjHYdkeBU9xLzo5rpkGWtfxT5NDRIUuDePgceVqrfkBGRwirTrhLqeN5SKhhQAJ
JkUgyh8EWhBkQsaVLpuW0ngy4xiYhOMcN16F+vNzXOi9qMeUg2uA08mdl1OGuS5o9lXQc2vuSvGT
WamPSv/3B359jtAdXr++28883aZbkfO9q99vHDo6cOlyV35qDdm4hgd1Zf7j5SCJAgAQoLA2njxA
gH7F0R2SC4Yi6NWHT+PWtiXkCahe2XJdPM9UYqWvi8A8/eYSSno1eWCWUgJFQ6nHakS4xzJjd5VG
9hyDXAMlUBOuNhtRBImX9bCGBksbDWmWlrW7lTmsiPmrcnxOtUqOqR9ls/wy7n5IN1iu19VyZTXH
88m18fRVsyga+fYVqDuCah3MCSLsNyt0yebEo5/bTyDdlXPMH/2o8eRO+UIMPRDIFqJ1ivNxao0E
1jm/99FI6+P5KUn/0mndfZR4bfwtCE/7tgJO06k23ynTGNDCqoEXxd2U7HuzfIWwIaCVITrETRcp
OGz1FV/ftMYNsY1MIDUs2IZUnH2Gpbmr00h+cljKnGaDteTpflBTfqXnmQWUumLzucdamfCahiF9
UbOOJGM80ehGCmCsuSw1FNJ4EvmtNDsf5Ds/OhRHCrGSrSgS19SI3eoLDgKdYUB9ibKSBKtd9Dxa
yGHuDL1N2wKuNop1FxVvG9CH23RWj1cHbYHA8gJ21PbekVWiHWKH+1H9fs5HNG8HqwAtOiEI8i/Z
wlXNi5iaT8tUggrUkkSFBRgssAFkVTFK702LVNmMOGMEeABT/zSoJFGGU1eBGFg6BBKQ4aLXjLlV
TOfQlGxM4A5Dj10OUKSv8Y4yH7+metNGG71dQ7EUD1XOALyK7IufGq4MUi/q2wZe0yN6AzuRbc1x
kz2zNycsRHZtHJTTdPLXx9wYBpmTy3bajBl26lwD6Cl777PzyfBFeoh24Tq08t9y0nGPMqL2O9O2
q+kPkbTOFogvW6tLj+CGXI2HgCcvCk+icXhJq9hzSR6B73IDZdBd4ZZhNW293oNYusnEmBspnzsn
7z8PkX+aJPpXN4qbFF4KXCcSE3pE1VXAjWYH8zhHjqE7KwjpqWUs3IALBkGh3TA9WmJ41szhA9vv
DuoD+YVdUN+WGrYC8d4mY8uLXu5EloPogkuqL2PkyjIhHOyf0Z/KhbnUbAJwthhkLYwtJCvNNgZh
QUmXDPT2xHZLWytSMMR6Aa/DYoWATwMpWuAbodQTzdIbOLsDV3GsqQCxXVz7AijIFMAbD1H/5iSd
kiEs9+DEVukzua50T3ruwU9g0dap8jt3Nc/qxjTiPDheXFn/SDPkCqSinfXFHcYJmlpuQ1qcBmHV
kA9heWTFALPQ4WyNNCeggytWhr9y/XWn8kgZ2HuMaHGYAsprU1XUvUNJxn5381/G4B33O8SH0ccP
nyuRK5DVtfbHLQgtDQPMvV/Ou2IOSAhR7UYS04vaBUPhcGQL3Rlts+VN3XAmpiU+uy2DTqYP1nPa
cN8VcXl1zzk2oL9PybkWL5dFTCC8OuW31RovOzvf51ibAIPI18nxXwe6uji+pcAMFxild6249ur3
r0P+rAmPNKVc0/YWSt0qpfheoQTYVMr0+vT61z3+nU0vcg1t3zaKU2U+YjtuMznhLyJlnFYMRsxu
Y1t9+cBX7vPU9p7iUEPEyQurKUf7rVJN1A7NYNtQha2VAPUHrWzFesORVl+Bpi75NCsqe09/nm+E
BstCENAr6JX3smYdCKGz888/K5ORDkuZDUQopJNMyoeOBKyFV8GxdPOKKTt+8ZXEkQZGmynfq+Ph
tcfyAACzrf4DCQYGpQjChNHUcY07SDyOtUihPd4iN1zdPqvzg/bgwfKiZV8a1bNw4xFP/gHWIhS7
4cmRCUvSTccLKF4O48z6StUIEJTFWMZ0SkK8dC5ml4YeID9X6v+dK5kbo0cpuA4FBAwwNm2eEcE8
5rar8GqGmuuFKWxLGEaN7HI11mGw2CQMaFKgnF3Ybw9M547WHibjLi+G4r+tYb943yRwRlibJy21
Sj85XD/hNl0ucCMCTjC7HVjvXjP2OsX5qILM+1xQkeaIwefqwigV+uyuYK7s8Lt9TsDnumkiqC+/
YzFIJpF+8GbWSeqr2oQKFHI2697MVU8mFlSEwFf8y+nK6sJWlpwqNFUfkGeTYSJEvXJfwr5Tc4gd
bhhc54s/AGudsQ3MfT8HoeLxTrAZYLHicKlcVkhznXIXt+iGNMtMg+vbKN7fYmHVvIfzCPNC6MnG
/e106wn82CDz84NIaIo3ZTcfkfI/EbeeqdpKThqXFu4wUzoT0jSnuz+Ksh94KFXCWX90NV9nnpEW
xNEbAAF+gEi9xWCM0x7hj50ZnuwBstg+70Me0OLbP47ddDWWvxSB+ffD4DIXpW5ArWOEmIiXCJAD
zL/vWFxCzR1Vx9GQALIizbf5E4l7QMgVZUZEAmyolSYc+2dX99CxzLMHyn+VFpCAIvTJjYECUgX3
1ntJsSvG+r5Vi/eZcFTVuSzcEIlmWhcEgBZ3eSJt+o7ifmWSTCleYMNkBqwS9szoqj+Qy8pKChvu
KK+xs+uPP3xDYc8EudD/FHvI2VNLm4r6pb83O9TIwRAHkrbdsVp3FU7TkSAaaO63SXttWQmH1lfk
jYDz9Cg/52MqyIodcv75BJJWOr13lY2iR2RMVSbey+2LlmgyHD/UwTZZJr7h2B1g8MZO3THOhdLv
kOgULDkA+4rAIwWEh+KYZRCl8JFvVKswmRo3pn8cFAEnl5lTSuu3vG4gGCwHyC/Q1qwxZMM6ONli
wFMEivGdGveDlC5ltHR3/3Coii2rN1FM1B8iisIvB4V3+plqewqQ1vy1DntFLbv8Cyno+ZHfCBoh
hGkp6rCeqYR4eHTtydPIA8EIyaxpvjEcWg9iVpRo/+UG8lDlONwssayzquexVjley9kWkDvRFBAF
2afrjuSQj4kRiDXqJC+tL5ToG91AEdPqkA9sD+0bvRP/nCFYpOu671ujPaf8hp4Xc5K8HmfSxYeW
/brbBLYCIdcn1NNThAtIxEi/icgU83Jy2N6EQ5QYc4pMEyHp8LTMwk3BDJaeHcbKQOdoUvHhxgTg
LK3bTwvj2ssycd6Bl0fPPIZHldon2pdxiE228czU20V7yIjjFEHGTQJh9NLp1+W8U3Y5oo/Kp3kD
mrRnjCBLrhvQsj2dQ78KjeA5zaX3MI4IDf0oRybuxlEILC3Du4t7vuSyk5wdsAPYvb8DkstrbQpt
h1f6laVq0dPwUTMvbBguCHcOSqtrJoOWs6jAt4cqrtKAmdUlrPWYllrQkjVUYzjT0jdAJlsSBddS
z7//xizaSOmV4DH5a9z3o7KNZEJPCjo9NniLXCpy7AtjjuvS4Onytxag0Ff9KGf3DJD2xlqSNcVb
UVDdk0UKsv6x27KiI39iEmJzwjLNeowwkQm0w98nbDUGIbabcYjQIZyakcZil+7QeBp/h95GSsfk
XHhJHKyZCX7FwwNGr9Im87pMZZ5iYoe/9fBwl+jOsBHonaCm75L8Zbzokh9+O6C8agMhtSDlBSW7
t7WYCGUkdhWp2vZFfl2HBlRvaIJvsIitDn0cKKjakrDJIIRPGy0xQdDUVkrRyYk5VY55nHNODWcb
B94fRSSm28TC+KfYOeB1CMZcneCFUuHQxsLRMqBDJ8+zc9EQla3uTA+2RwZ/wQbFSaPR/w9SHS8q
Ws9pxap/jeuRTsGHNBmF6Moua/D7UQPo2lRETbA8A9bh7LS+7gNrLJQMaQVgqA87KRntNz6jLcra
uZd0qGdfgL7O07nc9/GJlbJiYvwh1pWpRwix+wX6SKfWrqK3mPGVaEZK5SGs9y12JgdmYt2luu2k
b7MWSDykKbIhX0xh6ZJsZBQTXJHicODu5FhjAgpuobRPS024BXCNrskT7+EpmOPQ1xQg1D0grRf6
E6UeGsDArQPkVwLsddDTQxF9GzCXVcKLrmR0zDljgy7fyNZwMKjRLuiHBICjTp5Y3xcICg1U9Vdg
aqvKUGv93BWg6Jf95oFnvoC2pU5WXWDBT7OS2tcG/q0jfCN1deqUWdaUObiAcnStLtkUk3kcHIy5
8l/Orntqo7FxmuKJpn7+bYQcicfEAI4TY1nvBzqQKYsMFOUpM5ks9snPgGuKognXbkLZJxY8m+N2
I3MaayZAccs4B22hDfJJMaoeUK1IDu/357Res2inyD16ATn7RlDFbC8sHseRgZ91jwhWp5qMgfTL
qRav/0D9nY/1la41yyo0Aa+aIMIsVTxXeUKkM+cH/e6geJlavzRrS8BKqdDF+158t/bhFx4Iqy3k
/8wZMhfeHTPRQLkjnDNeJqJtqgexfPu3mP4L0xxhyELkZMcYT2d7FcEne0n/bSZIXqXbo2LQsaSa
HToRYCEFYVzpyXkl7YDPLvsVOvvUdjx55OGklWOQjmpsWx1IT1qNuWBlnviDzcdDWYCBw1GSk3xg
nGFVI7aIWxjcczBPeEyvNfIW/VF6nsQH+sBNpV/BLtnD9cNIm8UBa6OIs2mm+FTM39lOVjZ4SQKM
j6sMWflFBGUYupXVuzWXbpvxCoqYcoj3vuD0LALWVP15cVu4zi7HNTmWeuFuEYss/GOQwoabE0s4
lEpxrjr+6rqHGtHLI7GossWKifuZ723CyJXpoHUAwD7LZ7I+wQWyN/TR2XUnj2M84YSTfoEPtKeZ
rtyAyECsXWG7dMuyOUMOwiJ5x8Cz8dr3IwkROHpT/Tk0+PqN7YUi6ZcE/rT/BqPI2A///oUR5N9P
C+bVRzeMk4WiGKRDqF2SYAsX7nkAJ12dfhJnRaTAMm6T/EM9/4MIxXWfs6MhDDrOHf2mxL+U1dHH
pOtZ5/l5WSMD+7LWWlxVbNqugXhXLpYoF8fbYR8mVjhsTdI2TN0xkr19m+jM/f+xt/9wEFAfr8Xq
0EgNPMJreQgqg7y/0oQXHnIqg5KopDkm5uCSfgnJF+LJlBhrrQbX0At/wnKTeN5w09YlkOqhbH4x
NwyrHtG3NJ1LMvPTVz3B4gLF5IiKI3OvHnxm/RJaUlnyhSdNP/HmERBam5cHoSnX1WoN57j692DC
t9CKycJyrKEwKRf/yG0sgJN/zM4hxBxBdETrBwefznPdK/RRwNKwO4/tn/VzvUPeJM9MmqT05cId
QsgdEoiTT8IzXOhnLAVC2nOMwOsp0qWQw+TviQ3byBzn+BdgPB8etciisV7S22gvPOar39syK51Z
7rQmdMy4zvHfy+1hdt7NUAUIKu75GfEsnEXaZJmV8gsqyR+rQgM1pHp0uca20n/foK4f73V05Q37
KYfI2T+u5UuG/x9ZBqcM1QxYY/vkwf0EfraMbyDFu4gcE9+8wv8zXvt//C7haT1719T4IE0zTfJW
rklzeh+o1kUyaVnE2pqU2Tz9OIudBjte/PXdEkvnXyzXCR+QRXqKu8jlHcsPaEyLZ0YIM8bx6gkF
1HOMV9+nI7iYOXAHbYYYnkak1UOkXhXUQbzogTPnT10vWj5maQUG59Z4m5nnnPUzpqIFwHMkd7kx
J3oNYBYKIHTuo/IdeFQiwTX+I21dAUtZvyiFBQrWmionm5FL6F/sImtxyAubXwdMfWb8EY7609tF
NfNvcQeKca1oC77PePTCZUsdg6PZsPcTIcjy83HL8pjGtkvnadnEXt9sGEtSV/QaKAIwusDJF8Om
mslUhAB2Jymm2cj+gWbnaVO3iwzyvP8wyMmK+yWRWNuDfurSQBQgmWoVDjHK+5dIB1JaY7n2JYwX
76KIBplFyB1R6WWkkS5HzgyvN8824XMgKMnTlQQ7NKoEEpwlyPpOpgsJrDHwtuwjrF226RHIo7l+
pnkSY6G8zjEjBozV6/ZmNCBLgQ2TFBzzmUR1kQXymnF7nQSSFG4MB6jLUG4KXmOqXn5QEXzIfW9K
lm0Lk/f/UU1hKx5B8pSYGHhFZQbp4q7GZ+9H51++zgJgsHAJe3XMlZcpIlRON3kxgjoPCuOWrU6H
aKhU27QKd+MBDAsCUs6yk88DD/Ah9y8XLVQEsrMWPyETRLYoGPhlO0dbRzlhdm5WDDwIvDB7wTB5
YFTp/ivOUpYrAF0LFTEcLZ6PGZq/0UJ1KTTJt2fvfnA9m9HHT2dUUgCKMIe2QnX7A9vi9/2UhZgu
i6GocyWrc29HmtOnGfpurgCS/IkyGeA2X1sArzB12uuu+Q1ig89JQCY6xk+dL83lgjaSnXtxjjWe
bOVrV9mbgtAiuM/uouCGDP9t+2MyscaxAR6rTksdWBahsMC/ysqgA6qxEdqG6bg57JuSOaIWtXCm
fqWQ58/t35TkTnl4sx2wOhptcOd6dtHT7cHCIiuy1ev7TbPymlOFBL/2X6sxslTCiSRHTBcX2NOv
dUljIPp0SUzJXDMOqSMj/wyn7vFBeLgMIJOZjXMNIkHAkKxXl0livTSdvwfK/IttRgfdpgVOnHqH
w/J5Lidvem8uUkf/dsdciocGufP90V3F6Wr1eLd+6XM0DeHRd1cwOkRN5geOA3wzwSGBYaUJV2OZ
a2zKDcBh4IvfMNZb3qjFgouoXXA03iSlPq7aRQH+YImQhsoQm5Y7K0YsPbo9NdwbfCvbYyQM6uWq
aAZHVRdkONN+OLC0Vd3aywSEQ5AQJ6qWPx2E3F3NzokyK9h/RpGRxtXj45FHkK1UowYMfH69br1K
zxCAAQU/xUzFIw3/9LY74DRd1hU6SrCG6d2y2MMRqtfLJLk2942RezZkPooqWeNVc8lD3kzfK8IP
NB3Zb1FPWgXtk2COvaOOLX9fsgrkKod2kaRvXfP66QIk33Lnnt0n5zW9gEh8tg4Wv0l2iNtWKfKd
FmFjl0uGP6/U+TJHIWpAch000ExYTQF2D+sVmDaQ5HuSrJ7NBZwQkRq/GbmE8bbzznW5UIpGKQ2R
JuPCs6rZ6HrGJPSOAuncruZfrLkxGR/Ao9MhFmtn6elQHWbpgGz5Ea9LRaJJYokqvArOQsLfZ75w
QnF/4KvfO+g8ffgx9wnOHubrM76jd62lB20ZCP76VqyEvQI84qzc9e8zAKEe0sD8hOEXFyXVC5Kh
SB+LvGuI7s3ggmrui5w6xCSITF2bOX0e/4/qNba/mOpdF6Czha/TmvJ4e24aYjw6EZ+ijXpOXrST
Fvtqoqopnt/fJMJg+JEIUMHG93wb9wxu1vO8tMeSeu7LudgHICoVDz49hUEnj2MkygYNYlwICzqv
cpmEbXLPsUyLgfViO4zsEV1UbODp9+/z1F8cNz4UKIxxrS+x+UtBguaO18/JPeVaw8vLAiEGTO+O
4sbtpBmc7vGscF37QzuksJV0EQZ3v77dCvTIyMHCkH7Co7Ix8O9R9t3/DmwWYEJrcafI1oQDPVLI
RJbJkkzVwcSndpKq3RNOONmfgh28MZ14L3jO1YtpJCfOoiBJYs2hsGPLxnYM/RkvrrB8uNYGkKpO
TFjBf23R0PUqk0QpNNFAp82MpUCNi3rREVHgMkPjb54vDW5xDzfIDsVYHyLAkJpeKst31dOgjixr
pv/h037HFQ5owRGAtTHgNrjtXKFxFfrraIAX1dLh+vjZiivKJ1xVC/fXSB18OZbIp0B3nQ58dQDf
D40msGRuFMA87/rYkLi6yquIrAGCOWPkLo61uzBZn8UKkcfxTQu+4fUsxDoxeJLd1IK8uEb7PDnc
mIrvIBLzmtMotUTRWNxpB81IXkYau8Zgqj6DB4+cw9cBpcGPjImif+g2IfD+eF/dqUUvuJVnZ1ZM
8c7LsB80VONwSilb1G0g2f5JQ9DI+qD3GlAt5Tlsch79onqcOlPD70jkwelwkK/Rhc2v9Hvvmwan
qIeBkiqRvgWc8RSGHlXd+eyiqg/aIAP+wMTWy3vfXyIHaEyPvZypo5SyUdR7jmGWDcMWsNS7t3iA
bX0jLGzf0Gf8PjgsoAvNxg7i40ZArXXzpIXf5GJhv2jrbmghoKmCk1KRCKAdLFh80Qzpbmzkj0FD
YEvspfeGk6tSBeUZ2KVnQt28aTRUdQn21B/bvCiBAEsYrUmFrcFy8AonsFzXAXQMbmrADzQHYJK9
qCRnxtwdvueguJ/DsIj0lNnMP7MA0lptd6s4LCElLfKYCK3qK0jLEhNPcoAN1ZWK6vTr4gHLEN4T
A9CGKLUsDHeOh/ErJRYGIKfuLhyPMOA8ahTsDwg056j6p4cOwgPseqfCj2D6nbjCPeYus6WmFeAn
tl25xCkLFpJJTOL3vx0ubRg2h3dMO5IOpY6qtBz4pxqsaSyZQfx0j59kDN+alDDvMvWgUrUgVfDQ
efFeaNZRXDLQh6Yh64/6HZZKn+3PvNanAHJaTI4I9cP7dmI/pjtck9jatfU+oPndMYBhoT/BAcle
fNCvabE89sE+4+h8EavqGrCiWm7G3dbtMk4SN+4T3j/7XrLOCe3bK91Y4dhv6TmAcWv6hry5LMwg
VvhkNSXjqkDQR/kJlr+vfVDxH/yV8bb7BYDAyLMs1ipLN76DSGp6lN6yZyLBbIZsUu0Xi3vbDvq9
79f3Qd+nAfVYjybN8mFlOfE7jsLj29H4SQX8F2rCwsn1JzVAu0MMFmx/Vc7UHJYGaWHN0cK3QGxE
245uMn2opAggd4gMKbOquj/dFDRozMM5KYprNo1cYL+PrOBGzCsChGaMhW2jwPyDepaPPMvm8w3E
DEPnnta8o7Ldl9+oDuFlLSpy965fGGgjieWRhHb6HbE3lsrk1ouh1UpRW3dEuc/9xh6n5kMas/V8
PCkKpa6HD8evgk/bkme0SAy/72PS5Ggd2u4kc+EIy5P3tJyDl7ji5g5ktlPUPynLPpwVWOg4sR6/
z3xEuHpWR+6cCCTPnAjeS8b+QG1eE2iP3LmajDRze1IO20ecSRBBK4VGUneQtwEyBPP2bz/ZYua7
gLJimOyZTvakT8IJIZaHrMwKAc3NO0L4rTE5O2j/bqnlkLA/o7/0UMqOOmZeShQxDASd9TOkDy+W
wa1kB34Y1Imj4QaU37QjoFdkDGRfplGkiQQlJY2lM6/eDG8EwfABSGWKiHPylKORqcVwajyNzZ71
NUND7ZHVdHImGQtF9H6h/65uNx1HsQf9QIbzP8RWH1nxHh58NMC9zmSndb+PjS2JPvfK4TF6MJEm
ftZj2n0YUH6M1E92shPEdePcaCEt4vlg21G60e3RIq6vsxfQ9dHJmsMrRX20lACeb3vQ0LDwkoek
/rXSU17ZMHWdc5/WkKD0+DK/suW2tnk1orrajZXPgdaPw/Mfre+iLJICBdBcmpOtvoyMgPnPqaYU
YK/AxAbU08hYrTT6wWB4/Z4wDN/YBju1FkMQnTyiI/m/OtOrmn2f+foF8A5H6W3Y0K04+eLC9U/F
w78hzCO/s+Ce/R+ow0sCnhFduBvgpRKePdMieS6JANGzWGaq852/QU5KF7K87IGuQN7NgGNIzQdg
rpytYJDHwiSsS6SdH77S3H/vG+DwbrCIo64NnX4LKal6nyJgIx7BwMjlFjSB4eXA96C3wr7BpZWT
2vHMRwO4YFB+a2W0W3NzysmLBVa2pNy391upqWmqPXRHRJO7oyvA+oQLQ5FSTbBFm84NzWxaBl6+
Gaq7dgzc05/UjRhVz4wqXyp8jAB7XO6RThT/BdB+++DT2KVSaSI1/87SFPELfoSl6/j2teMWiG9H
gRwv6syFcZ+NuHjMCliAjmOlcHAMBTejUHS/1FAfHYraKqE6MdzCnOys2F5ihfhekU3TNUohkJWY
HZ+SsWqb1An7dHUSrhNbhSXroDi38QIYAZoosCgdi3FNkqHD05DJcmpQXQj69YnHMvtUkBYnwDVq
6t/3nhh6y55blKxt4o6Mfv1u91HBX5+8kUdnp2ZqxahrnXSiEZgmCx5V/2zH65EJBuxcB45SdKqq
ABqVC+2r9bDahsYolG9vs5UNJC5Zz/l808NrhNqD0q9lUINSrr4mitVG+GT4ap+b+6k3tz0o7nkM
XEuKIY4zMit+YGfLJiRiD/V6zrnw6leJsF2ZoPMlpT+FKvUyUH8pbBRKoPhuHSiVo3eMlJJlgT/u
YHBNczH+QR0Wya5uG9WZP0hcKuUoJJe4KsT3/qcKCdupzDJySxNCXagsbkULzluNUDsVD2dpGGn/
6u4CTzfoXegOXjUYS2WNBWYmM3HIT7erKaQkqvI1PJbDy2bK1acJCagDRD3d3iHhk4dZ89CT/ANa
SislH3EH3tcaU3ZRoUrizMc8kC4kNqjXGvxpsmzZPv2ImqvaDKH/hJNaNSX9qBCJ1215gbs4uMvl
Sg/TcgGm/C9QV/PgghbjdjWY5bRmYElgTI3IXoiytcJqdUOPMA+mVYvbhNQuMgw8ZqQrHvL2H9Vg
e/6kZ2C9v/X8kbE8k7etmTQnR7xQh/ZXhk7ftCU6LDV5lC4J76Na9++MwtdkAetp9oxxkeEPb7PK
IWJyoPTTuphgXJx3duRBCCX4IpaRX1PTVBCPky75cvYSSxDonvHMokp13J/94ZTy+o4Fr8O0JD5G
PJ3G5e+xxXWMGjakgLuPYrBPwf5lMvtKneBBfCCpLi6d7Uo+hNHEF940ZaaAGKArsohtwFNJURaJ
4X1F3t9outtCpMaQft8qKwAjKB2TN0Qtjav8PJDTVj6HAO62nzHn02nMCh1so8awlyZXG19y8xaw
H87PCkzf1OE0MuX7VUCZGYlCiwsUOPJ1iu48YXHMraccaFfVLcxJi+y0PjP6208UgSsEAtZmTaXW
a9dbk48iEsbNNlMARZmKM209/csdf8uzqtK1AjMf4uvNizMW8AxNqao74+xTsxqg9PSNPPu5UB9N
f1z80mlHxto6FqrIEUIweuB0CFpJlXuZ/BfPMINczw9EM2b1fhEwwnirNIcbP9chqFwzVxcwxrTG
NQbPoMUibiFLpRS/Sn8xUXeJPou5ycXlgTH0ywwvXlPQfaI9u4K4LmMiG275YqU6xcdE7kj4DFtG
BVnzRuahUaoMYhx4RbmjKBsWChBkErOSG2IcVNdz9l1QGOy0uQXYA3K2BW1IW46dxOxiEmiS+TAR
ELaN3TIw62msm6LlLodBEj0a7dZxc9iDEUkv01GjAnuZXqqNZiEThMcVGQlLK0G+CqSZKvUee7qJ
z/7krtjJC+G8pmoiU4fPQkOFTzh+7QOTkzukeQ8IATnCjbi7V+2d+7h5Hlg+XW5C6HyiPo6oEOqG
ofDIOjIisAGmQuGWmALsh4yPui5t9gDC/ZxddmpGOaYrqQ2cMZ2VgGsEFgd6PUizd1YyCTLoRooo
g01ndrC5b1ulaTTRJuzooPfSb8GqajPXE9B4+O+zVxWeCGq1jlGSVaqQC/6azdtmdVm33vMYXz7U
6S3tb9S0T0X9yCg8MowdrKyAUJZRvYSer4ViiDrb//sLn6qSZavs0LjoOKT6hGqFOwWtQLtKpBuq
VGitU/UqZGIRCZ6HZfhhjJJQyupc3/uz4fXcLqPjaXr1kL6a33XmuokLZSXIgJTlXC0M4ngDxVXw
/pHhqXP9txnLyTBCOCb33v8B6olrmcFZy2Rg91Ag2WpmFTqDGKGfPxqDRnZn7gaqy3zDvV6pBGGV
FwW93lMnRS6kJSgr5pkfbDK3MH2PO9ozJRHNsNmyhp395wXCShLIfik38gKuD8P9AtTADvEgKonS
rYV1XcwndzE44PXhOAc9dKXyHySqo9rq9/M5zIJJ8TbvaGYxGJbSYR0SbTZR5AZeLkgbXg56i8Qm
+4YTFZWLsUD0wVYj4w9rfPlJ0cvfOkjAEDbNRIaSbMXE3pabMsePbLkW789ToDkCVJTlZiXnOe0M
K5Jalowdaf1qWG5A8Cwj7Bq/mFlM+Y9uEjWv1qhkrbt5u7poSIucggXbnqqiRRcAHCzvVjkBrlcY
vEQ5HqQJ8Rd620jK5UbNLPmSF7vwr0Uz0ZwUlLGkkY8ITgN2bgFY3qjzJM134k0IwY4/ejiv0R3N
ypt7rrHUHMhut4zOhr4c+ClTTO/tHESeynMFM90AMQz59ChFFDBXDIA81lUZ1jprTtTSoGNq1D4C
Pixb990qureo+39o8/HIuNvKNnMPWDWMNCc4Ku5NhwxHp86ic3nCldjGsZn6PpGYMwYMcn0pXfoe
PMuRiuDW3L1bL4Q+y+Dwn5KsyLo5IcYv06Kl8xrf4QMOEGBJ4RwAJfwbN4uYttR9EPp/Y/KdRVlM
Y00S/za+fy7j3dPNRKWQpzfz8yzged74TistV2HwxByWoyiieDgeCrpUy+FQrI0Pa8Dn02XYFaLn
TJ9jJ9BGt6wOtXpM+4HBMQS1NSF8CvBKVucOh+Cx3Ty5ldmkilNILJAMn3SJIVj/77LJwpVDSH0l
1gR87il8JN/vq/MUWV51mz8kBL9Abn2FtOKEjP17OYMe8EKpYe9f4+KdDqwg+lWgPPFYsRKw5yk5
OnLZbTGi/b2nNr2Xj7R6GgKZdnfNsHwiD4rRiwQD7SEYVhtUrwfSKhWs6ZzZnKSyUcqUKkGLKVWq
eaeEVxjMeRG8SYn8GQSKDXO3/1QxfVfOXWoOOhbvFs5TuUiPJ2tVPHSOThpxQS6DT70HFa+Fy33c
eEkvHKAr4sA0BbiKceuoByUk1D140968clYTxFKu+7ZVVPGERo7rpy8uMv/6OjCIlyvqBdjoZ5CI
GTtKSeB2HkLBZIPlPEmySpkKivZG/mlJZg806HBTrdxwm9drEIzfKQZ/fei7j4cFgCJyVh9QDFDD
bFDJs+xkcnVqKuRTReJNBXS/uYOfLIuCP+kdZmTVDv/iQTPes/Aji+5PL3QNB9bjT89DBJwOcvnG
lNY0ehT+mu/5YkzbEFTQYVhDVE7E4dqSc5VTR2kiebXHJXMaK2uss44PwjYlghmWNwfE32M4kn80
vcflaSjdMnDoTPrsguKPhaQypkD9lxOk52pFXnUfpBidr/fvg9LnJRVYwTxbXpeqqv9vcZseagTN
9qlai0Th/XBLbXH0hZF9g7MHGHyvbLVmXPA4G+oNWzqz9Soy88YPLixERkIbLwgPLmQCPGQpV7JW
yXo/usoetx86+gp+feVXb46rtyjXH204ypqfgTbRHCwcK6eAv+c2UXBYx84FUL99GNqOtkSqkc0t
ZNsjmGRGsmZ25v8gM91WP6OBrfe/Qwz39rl2i+9bE++Lv1EjhkXOysaEbdVRsi90HbD/6L/obVVA
SVwTKHg54OGaXvMw60kliM15PiXAoTcAJ6Y7nxNfQiginl2v7NX73I42GB6IQ/1yi0Sly/hfNg98
Re34woj2KnAiiCWrgvVwmRrcbhKBVCrrL6oN5A9ufyy1ZPsbcnjuEC0AYnCTFX3uhYxP+yQcTeSc
7NYzrHskfPt1NUyQvVRoSy1VwHqyyn9Moe3Ds4o0p6zhc8dAxM1iDIbnAmzo0hqK/wPaEdAX+Bq0
dxsiokqAZNia8aWIpoUJsmOhure/rms3Jv55vLyWbnF9xNvi1j5Yo/A442SNl+m148d5jgFFW++/
WS6B6vrLr5wdCnPPeKeUEcaJGeGlMnigsIlRxXjih7mv04SrED5E6JLrXIJXyz31ZYL2yvnMLz/c
In84XDE2rrdP69gWOe/lX4wmFNivCnt/LlmC080+UYspe4te/veHGmJ45XLNiGL3bxlQ80qFWFVi
hJRvjDIiUkkEYgk5ujp2RtYdIhI4X4Gw2tHFgKtIC/dYvMIf1WiFs/Hl4LSlpYigU4o0gP5/YAQc
8ySKzYk5KbEqtcoPJl6Dx/qPr814yGLZUgk7wg77geR7okeUOqU6Tdi66ySCJz4juph1INujIa00
GymY1kJuW/brwTpAXYlNsLsVLD/LLmGJ1COMz4fNEtirVzNURiljLuG8cyBjmp2wgh4SjQBnE/zI
mVXPO99kbVrgp947+IRSC/bx2iJdKNd+a/4w+X47w++syNxEq6MDAQltzYaiVYrzyr8UUNnMdnS6
z53nWn5IkWObEm8crPZz2rBDRn2NCKSZWFRyaDtfbaa+0KTPxtdq+9DXU7lJOnw8vuPfegmmzoCA
oIomhSdkyscwxXYdcIX7MujrAR7CYAxuoOywyQLI/FCbx2wb9ww2lPLdxlAehfa9JXG9SaQE8Bpl
sEt80Xi32TQLDKKdNBSG12ALhMq1sNRgVObgF0IK/VB/j5/uLiKeUhHOVtpfCqTOLbyacuVhHOnG
4hqd39rXSFZpJx0ajAgjVzmLWIrHzvT0pt3y6G9uXOoPDskEctHJUi9+suJpzAmvSDf/BkeO5PYM
oRGgzo8xXEJfwzTRHqFP+ckp1BsBAPgOzypbPxVdbc+Lu7L7IG8PuWbQr2AmOMmnMvUaLKVg49XT
piXdd68Ker/9e3NOdmW9JUjWnGHEBERPkI7V4N+2k5eepoK0F3AnbYSIF+ZCGQptzKaXS7jQC68G
kDwU9hdwPITytm9xxH297DoUDY0dKZIfpdJmssTG9EG8JOQjkRdS51RVOnEYfsAXudhTk7/KFGJ5
mVYUO56yTr10uFAICTf4uIS62k1wCiP8pvEo+DRc30X9TmRMmAHtHysm663WhfLwz9wr5fXNpzxl
58QHIT5n+qWzFbM3xtLicf3RxqFk2h6PxLTwPupfQdWAYkaisbVrJyJ0ZfHJsUDwr/srK38mbQFf
ug1EyomI3YTo1KM75Lih6JamyIPsr9cqTod+O0xYvKjpBZR+wKGoCYmXmhJo9nFJ6WTNd64MfUuJ
XrqdydDdyWo29qfEoADLOZv8gIQGl84nhHF6qkh2jIqtqv/g0i4tYm8OwKgwX8ed+b8d7jugTAQr
sbdWS5XdjhRqP0tMS2l11njm/wicxGS7Ok+gHNHeJF0MjT5W8Rv5hyLQ4JAtKY5GFC7aaNTpUeJX
B4hfTvrj/N5jkXd9dXHF7l3s274bWvR5XG/ayWQZ7Uh+Z3wcxNbTIQIYX0QolyP07//aJAa9XDo+
P4tqYbx+SIbm2psOmIiDgUxIBARapE28ybmT/0yhcO9o99Y9+6fwtNA26Lt39btZiuqf9lthCu5n
YSTfxr5lFgUIEfzf1ZomO2wemuMkdYoaBWNOoMJIFgH3pj3E+1WM8MPv4/hsDdEI6ApqaxJ6aNb6
y1V96u1djpgnq4KDi+Pg02X4xEx2dmXfJ9+9B1BipCnPGkRtdk5FPT2bN6zmud+k7kmVsP2mEhpk
FnFuSUyy9Gkvpr8RuNKMHcBi9XBQubxb4pgLBje4P8VYAhooO13DAhy0u4PNdOXbPWCbQ++rlaIB
75S/6HcBpY9VFZCONwrz5u8pIL+vzjbot1WygACCZ7CAv4mP6+OB1AXH4Ueuh4LHOFGTQDK1IZXq
nT7DOy5aHLgW5ilRLEb4WMO5Tt24xaGWyY7jncYMfQxZXyfBke1sXUyWanyIfs3Qkh22KIdgepmk
ltt8XBYMAUIocxYtOmLsFUW5w4YpFMN3sui+WjdeuGubgeAK/EmonfplkbRDakGR1OEmSymVsROs
gfv6Xh5vQTAgj3HcQFXW0cQLWCIVa+aNVc8kggFJHIRNrSLpY+fo9wch4TQ7UX99dTqMm6YPKA3Z
XjqTsm2q5k0J0WRsxH7pAYJDT/PRKBZWuAvvWmyYFdPt/BubYHUop7Bt5gkE0AqyDGRh1ezlSov/
3JLIHJOpFeCIPX+BvM6OW1AqLvvBA5UllrtYlfHIfdxXTBjbpU+b+lIzUXizNbwaWzev4NOQERsX
q7v3acj8C1oIf3qdjF5OHdX8gCQ+pz3c0bM4VGv9fliN6aqlKKxp6HOY9quwMkTAFBxASeywNHSS
oiQSzLKJcxa7FC9e0Y/FoVXyz/ZCjOKt41CNKOPlfceVB8K9wwPXJ+bUI6IQf2AmvGiKgcpqT8+T
6nAMeGsjaw8IgpGbe75FFSs1c+l1ytgEVxk6D8m4Aowbh69Zd/T41pNcTaNsn3Oa6d+20NJrKwX2
d49UWWEIcjNZV+uLyCUairB2OhLgEX5ns6Vy95Mx/6NPu9GhTOGbN5ogCmBIqTlfni1yrewp1QuI
IYphSbEF2mOF5smwduMIwvJjSEmSS74kkVRimU+zTfIuh0yBhRoKbeW24G0Hbf/aOwxX6Qn1WlVy
WlQocHYb5R7ofIS5wgYJV5BYExB0MV9cdcuoWtwOUjVVQ02BKDoNUDZ3TWhAI+L8WOMZfpyXtjpP
HNwdGSxORNxGni0uuPCiwk3k97fELIRWKJ0xTuPJC0+bZ9o0rZMN2r1gC5VhPoExwU7GZpXeNuVe
+PLI2zYFnqBBBhWHJ4eiVLOV/BFJ46deLZlSjs/S6ko8SZw2EHPMlRYHOaPMNfYDg7Rb3QGHz/Jp
ZcZISGRNUBrcIiXCezad7sbQOkxGy9WCXKTg2ocFjxq5NlCWo/ha7+ZjXUfvcnIea83n5mO/AfD4
xm2ve/tbjiXuQyv3Bwi6aYDMKZ0q6M4izEhtX1MJqUnD3Js3Iawbk/jbUyA00iPBwV7siMe3ECXv
Oy4Ae1ugyq8jzwKVxdEY3JEModXM187fHnnqJSPmUmUgt2D4iyZ1OKpHBc4OL+6kFn9GUE3CCNmD
zIf9rXq9U8Q9quax1bsICMUAmctOncA+QniwuhBhsuMKzQQV6ffipRjpZCThJR471HQRN5gEHLRR
XC262HmDCfIVo3fGwf6y2KGRlqhHxg1arYS5s6GtaaEpHlj4jSAyahLKHOyZRhb9cAjt6ob9LDIj
s9yoM1ayK8sy5LGnXfYiOQhOKI731vf1wsdv2wKPNzPppGliqzQ0v7Zx1Twh0x2ZbslHGZTGJSpu
sTaWcHadtBC3MgtnsM/TlSr7gUI00JEJZiBquKu6kUcesquBXcV+u5iPkwLbclnbaF5uIp1tnybt
2OwJrbIicy0QINc8BIgS+TY3isQBS6CpbH3Blte2AaALcsn1sUWtmit0JFleTfbPAFv3xIsEaBmT
NMpG8mrgAfHL2JG0XZolM27fBQefOb16nIeluy18af8L+GKsli0QsFvZhFHI7sJ82ZV19Hd2riyO
xEIz2/HFxu1Z13cp0mxooG/K10tTI895j5/3cfGffCNebPhA52bWlURLn02Lsyf2B6BWAvOtlS5q
kMtS7OHfjsKNEXE98x8zmfPpqCK9exOzvsPpbC591Ml6M9iKBnPO3o8BPwRFLSwFtMrUwv1dCRJ1
SG8uoDN17cs532oOSYffAqFO6fvWSkE0H8RzOSO7T4WXTasO8eZ5QaFOoi4OGiPxU3KzTnfP7bVm
2GxBsCHwVk5gKH2UmCe161RrLiGcqcUsGnKpiuI4eWCP1e/sKjDje9nBHiO3NSD64ilt34tet//1
AY/AqnyNBBs5QbJJP9GHGyTp0buoCBLMBF0mQ/tgsdu7ODxebdVF8HVHsP3hwXAANF2WoECdR5rL
DgmvFoiQMCinVLoBZ/ivLpsPCLiJaPniNpPZ9+KefGWxINhqwZ9WQprTkL92Leueu9ndVLNiC4RU
zIM75hKzod8EJkPPRkbiOCDdCfb7OJB15xmnzBL7paRtKlCTvRX4nIaHJ4DjREZrODSA/IFuimSR
scsGLqe4vXvO3nB/B8kKOzQyfV5YE+nTcuRP00k3rKXnAW0w9ZpwwEzojU4iT7rCp8d/zC39kjSI
tpiXQB0m2AXHWwIMzckfyjtZe5t9gCz2X7RU/qdCa2bePX3WonHpEM+Tbd8R+TNVHX7yM7m54t+O
wa/gXLi2YM0iDB/LW8jDtVMACoHWIIZYGKVDPls9R5JUO7uPtAUcYohieA8dZYBDZxkzLcxlos8D
Yvnv9DIoW+xuDmCwVyw/E1aPHcVd65rGW3f5chGmOvDsW04z0Ih4h8BBDDDDtNjWIw3A9Lqz5+tq
/VJLz4UPYT+LqQyemLF2k2q2o/9d1F3LrwEoPMXvxskJnsQks1VZHQdGAz+ympKKhA5dutFGhfe/
7pR80hkBenOaM4pYZ5UFXd7Z06T0STpnxn7vKeK3EFEqUYfEcmP3s5RZuh8fkwl7ZifEEGuf4/Xm
2wzipJrcXI7C6Mq9McNplKNaJGj/ZWFfFVJ5v3h/QksWYAQeGHTCtVIKVlur3DZKhS2FlVRPEC/L
irO1zuCcpnrr+JAgE/soJlkQINqnDjZYCxYgKqKsePuIRzC5lB6rj+bQU21LDdzlUZ+yRABdjG0+
cvgZBhKrKL6SH0ZpKXELzgTrRAbz3n8PUbprgb3yFEQ6Lka/so0CIPaP4wj0aULN5jEhWYeXyG4v
MvXjCUJdco9CA2upqvmQEgA4uO0jAW9DUtRQVkRkQmsKmJ6WGx2kqIJyOuyGoU3j3OrhPRK6qSuN
HD8lFpX68wHyVyI8vDWhMEtIAs4+CKjr52Gyy88xz1WfqB4E6Nbjt5ahofp9x2UadUaxzV4qIzbp
r32K4B+hRKvFFrFWelUDhbta7lCUf/N/NTUxKYkgZ3goR4J1xLDsQe4lU0Ao4GuZIJwvweHwrB9v
5z0DPaqgEnX1ggjrL8SpaIQTiUDYiJHFBcvrC6CjhQZg7MKVBu+VsUUV8+lXz7t2aC95i0rOxkks
+h//hI2NvriCumd4GCGW0hQhRhBba+dlBdcVgpH53rlEfC7Y8GTge2IcCIInIYHlfypHoQeyI1t1
bcBKMgThJtikJu6HrQdKe57ulvFWEf3tcEeXaK3sl6sHmTzpiu5g4rKZmOeNp937G4MVjOawVOEg
ptmQiNjHQ0Y+HO30I5UNmyD+cfghTYIjhTXRxIRmynP5DBkj+1ptaWdk58FVA52y9sZF278uZDpK
qPBlrdDBk795MeqXGcxK6+8Jm6gWT/DIc74MPzxeSMl1fHazX1cD2bEJ6dcqBJnBu0TRFrvOsjw+
ACJ3xpiPWv5yAAtZiCmHyiRqFQ1SnMh2xlApWyBT4CCttEgwKSPafYQa97U3SHRt4dC7xMg/DC7r
eMSyDfdO/OguxDsiOlwvsjIVu/54nRfkbUyA3HmFBiPpzSDgj818Vsbg+Hj15ZnqexujBm3T+h35
zkF41NSv2fGg8WQ7NH/smTT6omg8zMH0A6TYWFMObmh5aD6CZtUCVEdEMRqmSrDmyKXr0wJdh+ym
j9+CMu/AD1+1qqIrdDEGi6gRWg0qQGeEDVK1rF81h3eiAkZQ31jk3IF92QzjW6yGjGpeQxG6luId
2mGws4ihw6tY1+jg4re4ustNQGV51Osu8TQmfP3LQQ+F6QCTZM/A/1GDDrp97AspvzSA7AqlDVsS
UuOHCkWm1eh8ZvlKInzOA/v3MkUCX62vws44Ia8OtjHYMH4A4l4lLpSZ4WLWen+zt9cGfAKMbIok
psaP2AyP0IEuHjOAbsmCOL6LvAmaXq7yRCjBGQwWjj7Xd3I/87gux6lAE50t0eSVI9pYxVWAIXYd
qYaIlc08Yvvdoky52pz3GtVYbqrk5W4iLd85FhUM19OwU1I/DsKyDqImd5dZtaN92bp5cc/W/TmN
2IJgLM852PBHQUncZAr4EOf8UDZVRfqu99JRH1xgbHC9g83f8iFRwq71kjPrUfHiouZ8pTfwCMIP
09f0Myo4EaIH51ntiWx/lsbxTa1bFx68mMDnk1jafm5I70Nfe8hQq7pN5AvfEKVbvz3H3HQmtbIF
/hkevS6UriIXAANKhZLOMgEDKv4DF9xm+RzAZDdtPqAvrMxvtFcU0/kht224Ckoftk9o7o57JVqI
UP+chODrq2BBduZggquXxrcQp7Y5ch2QmwgWjDCYDeqvvStI1XFH1CehqxFA9Uks0HRaY6PBjdTC
wJ6IcIo+JeeLA6ivAkiBtoZqWDfeZvC3BO5C2FBdWwOU+p/AAQN+vT0BvxFGbLwXrXHHk0rlRyba
Wtr/N5Z6wS+MgSpof6ZdyUbnrEIK4sEMN64o5ghDBoK24qcoP52nFfPnsT9dnGJ5hhS8PRogcbB/
mRS+lzBZ54RMtB9zpWJpRuwbmcaVViNARmkP2sXv9Sls96BbWTQcLi+nsPISv2FVV5lwGTXKRDUG
k3I6hYhROF7dhXyVeq16WA0J8MKJpb2wQpLP0eTuwlLYZ3KZteKx0e8cRvYcEOYklP7tbDYASj56
+T3g4pvr8noKIwNSzqANQnHbexIDPuVFvxuExPGspGMfeX806wRSEa13+XIp0sKFCz36xqsIeYDa
3pDXXiI4Hh1brfFX1L8YNRvIn5BftAd6dX0e93RkD8PNtIDm4I9jG2OWd7nKU6xnhFMOFUIGH7Vn
5babN80Y+YqnijShzDNP05GttuaVt9oFXDO8iLc+HJ/2hIyNiVuB89jV8Gj2nGc8u1GXbDuu2Emk
pu0cSk7KzJ7nHJC1Nficwg7sUXDZY4jI/KpmLq/WDkxI26K7WrkXag9MUQNOszlwSq7fDUjI1dg3
kXyDxJQpn1OBOMTqoA8XsgmGMmSgwERdw/o5uC05jSn4ASArPwID5mEmQ6o/SZ01b6e3awrs+kAM
0t64qBm8J2DA+NbR6TcRoRuf48OkCLlsR9AX/HCmdT/SwbMQGE9vq+/0czGX0BfCoQz8cTcuZzdA
+wyVorlKwlj4Q8W316CuAQjUDMdNthEvzlnt4W/Xj2hHw4cXwbQ5NSytdG0xHyc9D49JDmhFZ9Fl
Nq9g069Aj/2OZL5GeBHMK74pLeobvikS52QFbotvSWxJFaKW8X2Y4tTZ9tGMUZ8xp26elsouT3eF
ePT/QPtc+6JSbG/aVr1zkE6h6668XO/fDm3AcgqWUKH/AjWmGGbG7So5t1pWZ1y/ro1fBqGeZo/W
m+iiy0THvEv46c6QehlZ0HNLlH+BaKFfFlD9ISN82pGCFM6r1LeaodOrgm1f/cm/y9Ek8hlM+yHv
cTgK7YDB+ZlKNMp0JwZAfD9zu5TcTJra2hAEPRag2SE0/l7Z2S1ONmAnfff9LJn28k69q0jRzkwu
bbIJL5gQIbnDzd4K9BppF5k/m+AjtahZmfZBHTvyzQH97epbXqvrJ6ln4tuHG7ABMGdt3hdlxrkU
MfercgICU6HW9n9CP0R2UdwGtG8I214IsVLo6N2RiSc76tgATRmtwynaTNU0GcmlDDjcy9XyueXs
Yjg2bgqQ4vSoJbXnwQq4D+mTygSmb5eaTk2juz30CeqVoEYl7Eh+1oEemvrBdn2PBRnCwtKmJcF/
AEZK+PcCIR2JJW+qqkkNHnNqmb5S64TtQ3NFK+OBUnLMOqYsalJd/l2mYT92W+ngWTGFHbT7nLy7
NFja0UQuoFnqRKEmxo2nHJQ159mAuPIsNg9B1D6qysSRnwkvT3PsIxcgkAWtnV74j5Zz5lL87AYd
QOr7HJr/jb016sZQGliHtYiyngGhp9/LHTEs9haqXzOGOjD67hK4hayp+jOCwkvD8PNIVzYa8AJx
8UZkgd40avS1x2QTpFO8rbydukvhUsGMiF80zk+0mugq9xyJz4gSJhaE1ryseUHP//nikyhxD9NL
05gP0n3VuwHyZQgGXggvl6TR/O3hSGCqSLUXArPBh/nhZb+hm/ZB9tl6yzS9ENirrv7SBheQIt/R
p4HUiC5f2523ahJ4cconRDj/wdQiQbiVrK/0fJYPswZerj4B+uf+6SIay98fKUH7XUx4gd9Kj32s
YTzNuIJMbQThrqcKknEydDptxgLY9xOugKo2WSgEqTtHwn7EZAE/XhkibWPSNoEXqQfkigYKA8OW
i5SdX7FmV9jKPVOpc2xcx889i7I3CvwvQhDqwADVdf0tLBNuGs+YZM8f7WHn/JAsRQrL4O1U1hI0
6NY5pyMdVJGuf0o4+f1/OzmO0e+dcAEVJeAcSgjECVWGyUMQNW9vtpBKluB0icxJLhQwgVDnqXNR
ofXcHX8oghd+eACNwAuIqzp1fdqwjd25Xy7hJEnyD9SV68lKCN2AmNxr+fCsR47mAgkfuLzKugr0
Y69tiiyxb+ETYQCevxcZKOOIV03uoK1Qs/hqviZJM3cUXQmgnGEepZq5eMol8Uo+mpS5oXc+Th68
pYCJLmFa7PWNy37SOUr5xVgM2We8DyoubwHEERlYlKI/KbRFNTVKZf/MTqXH0EUme/PRgq+2xcbL
wzNXjCDVmnT2CFrPl9dqlkgN6lQig6kyJBtv3O1tqAZHNWkKrhZNhJxp6snWg5dUjpPz0/+QeKFH
Gxoev/6Tst3I/Pkai+JKS50mCgXn3pg1tjVEDFQQLpxA1oQEQjgkYiE77iK1tyTCmcZ7A0jRzrCG
RmH5k9UAfgEEx3ulPiAHuqtrSBkpCU+iAWE6EkReFb+QuYluQPuH2Iw8vHXyk0KPDDM2TKwL/9K2
3/M5OpHqdvzwxu/EoSokvI46ggGENbc5fAm4ZFKZmk3JLTOmnzZtWi6n70QSk8ArUpBQhgS2OtlR
QaLSSuiiSValXhwjT2wiwztnctGjeHjJq3yvVuXJbX8xwP264u3huJr/By7t214/4ezdzo986TqG
9nBlRrtNaL/6cHQ6faFdCX6yGyt4JxTE/NMqjMh7AuvuDw9B6NULfcB7KrnTqtvTxdFrFfZa0PvI
7KwIyOUDlFJxSXj4p3NhCp4yi1TO+pu75zu25Wm9qENjLHkJSYrjIyjvhUK4hwyXSTbOwOKvTjcB
bU7E0rCD+LRcjrrJzMAzpblT/GtIFnw1YXPO7jM+6uxha6UXT4V0Y5+lOiMzxSAGnQpy5+8Klpsm
sqqAgozwTZgOk3n1UCz7CFYg5N0H+sUMFHR/UxJdd/44J4AWe/nH9/JyTVp6xVuRskHFAWaN+iHp
VUYGwx3C1msrk2LffC3DkPDT71hrMTPul6HyR7N4jFJXKWPsh4TgABDXhdP/kvQ4eAyNM4aDH1DZ
919sat/s5GOwI3VHumvvsAJsonDnkHZ0AVwV+3j8t6PhtpxIJn4HRo03NoA5FQMG0StfLZoOcEMc
74kKKthkBiDPaLNRcCeO8HXuxQ8ANIiXf4zrXf84B5Zfaa8zuGJ+wemrXq7eGhGwFo2aKlhBcUzP
Eecg9m7jQ5MgWQG9VWSpHD1E0M/GDg3CDqG/nultosk0Vx7XCj3WYvnUeL48OYbJIJxqqQ2khz8e
YNj9RBXM+hGjFKPeZeZV1QkeeW6D0Nc9WlFDUbO4/xY/aU2DsAKQngpXPkr5Zw4n/mDrglFqAbcf
iv7l5a1k11yD1BpVVNSDy3kTsMuCk8DXdTvEB3UOGLY7yi33NxKvhPkUUWDMDQ8zNI+ymOGyZm49
+uc7MxXwTVLVJgHE5iXoqA9PVi3iTdSXJVOSQJGxtdUXxWvgnyExBa3/29OF7+J8NnJxzF7uqqhL
bagZo5uVuINmWcf07h5PGmGX8JvpukB5VfWk2VOF0q1qhIU2MG65DgzplxL0MEcgUZ7Br5twtpRd
rx1dtrTPFg2/fj2D9NfzDBt5g4+q94kkOnWTpFr+y4BrAFI1xEkcshSzjcqpEb+DYJgT6+H65M/i
7B+AMTntY5AIgoN9bUFmmQ1DXrW/GZmbcuYGF+R7UYLLQ04pcRZsJMkP/RfLzOVtCGeslh8bCugs
5MLO9x/pnYzVotw4OHzb0P3fTiYImmPDD/Nn2NpIUfUrwL7fONUH0WJa0pwG2/EHZfI3dr4rocOJ
ivmt2+INDqATRok4ZTY8g8QAs4jbrRo2vzlTVC/7lnBcEFmArTaSRlRkYRhWyXdaKXlrrLMOd1uS
g7CKjaKWeMEyM2G1fvSIQKwu1kC2k6KhUQQs0CP2Jx2dwr4U0jGSwv6MAtOgEVbjZt+QRINZ3BQ7
l17fgMxDTAwLtlgbW5rakSPiT+lXC9RCrk7VRfabh4o1TZ/1yS7pdnAerGk9RzrOxlXtmFB6iqVK
9CS+GzGLNkThYp0yVhsXlnZ5XU6+JOHF2GMBSpoT13bbt9srrPv/Ybc4FkJFpo8UQ1EdtVXUhGeg
m9KuSbJ8a0bQ7feguhOMBV01xda0A3jKUImsi9Tw0TpGGee9iSdVPNrza7bnXd20Kqzp0iWmW7/6
s7vdmW9zMr0MyuNWlRGbZSMTqJV0HP0q7Knjd2zyhE4i0JDnt1i0rTVuHQoCL+sx8BReG4g3y2Ra
kDGxLCLO2BFvALcndKFnqSMrBb4S8CNLaLftSaUrN7h1NL1WsBgeavcbPR4PyX2DaBUdKIHIcK6P
GzJ3DCWO//QG5RBxNXNs2S96M1df6+aKdeR1+8dB8bBW8p/OvQ5OL4y5c/kC8YEtDjN5XETKBSDU
wWsLX4z6k/j/HxxeTMbpK/XDZVO8a+mVj4I9eg/QAhQ0Hbux8AW0EMYfnjvXdWnoE4boWuX9g7TW
G2KlrQjupeXm6IZuXuqQIjjK9MFgEfnh36i+br1ofGJ9Y5JDLldZ7pb7QzaO2dalQXJ9xtbqjcyH
pn5MWBAngBkXob9++uot9Dr6EeXM+9SbbQAusFiYw0FCDbbfLwaSLJDcYxN9FzFOjPIKrCR5Y5Ag
V8DjkL22H1tkikbq+TXC4B/+pfIwTZwUOAs0K5hA+b0oYQ/ZSti+l58NKBcfhU3nRa9OOCoMV7OV
X8BPLXpisYbYuZKKaGSm1gfJ+s+4PlfQcvpqcYejzxnFFCphk9VXwm2dsn4ZVik5OO6xVynHht9T
5xELhK5+wYihHpSNNCqpHpaLaTBBpkoo4rXWM0yUvsB70nzWWxyDcN/NxYT6IyQGn8h+iYIN/Wk4
TN5NmkMXU+48HkhiQLoimjeT8KrwvWlhCoIvfsZJa9IDdev3bFjQQQEMHesAadXLVeymcAdkCphT
CNLD/oR0nNnTQq9fe5kUW8dZEqCzEspw/R9iGs09ilN9xR9WZIQAJ3oTXK575YB9u5vXOa5iAopC
LtrXsgwerrhNx66QAW5HAq92NvX4ZlvYiVEqXjS50iyV/92AhrGFIFcs6BXialoczAqjztlQyxpb
0lGvCViOJsfmVObBO+oZqiYag1vNFPYUpXL52PczGOqSDGxDbeAfZGGugFeV9TGkyb/Jq9gVzKc4
wddygdBOUvA9TI+Nurp+4AhqI+2QMB+HovN8VVYVvHK+wgDb0HNKoGDY4mHxHajvVvAPTgLjE5lS
Oly3DEqbhg7IzMAhp7/5oNRy4kf9xoks++zOcKGtxlMoH0a4meOCPzxRrbpo8VKuRLirt+8rncSY
wtOjfNJwdkV5q0dtawFWMStDshoBChjxN26w4iyyKI9Sn/odCOKMGKdC7+ewS4pa6XyQ0GFsr5o9
M5MKlaqEwCEX2QJCrGD6RZ1I11+LnQtKiCtlOqumXeQTvKHbN/hAhvWamUU6L9LctgOGAu/6ZBH0
WPyoASecSmDsWHEAG8SD5gzl3FW/yZoxfthgjxHAIAVSrmFgsG903jJbzTOiEWmstPq+vyVrY71a
asK21TBo/Lm3bYmbLf7ZpMyTeJxNa5s5nkZZOgWZNQIIxWaAY2tcOiD3nJmZ7RY2IlGgbw6tVpWx
C2O3osvahJCb2lVcMpFW9jdE30+lWlW9VlIxH+ETx+4rIaSQ0Mjo7rPt0se1JkgatoHAZNQ2wa/Z
2iW2Z2cLmGFGaaFsKIq1brXbm2vluz+IutNMt8WUgJFnVBDeNK+9kCqStt8IEFHzGkoKxsOLb63m
71YNxzD6gyVBCVGMM+sPe34sMe8VUdCAf9hgDKLTRb1w7ScHh1ACiBTQnyTJM1vkN8bcGoxUlPxQ
FZXqXU1mhUVhKbwEhIGQl/Wo54reXgWMOmJJbM49kec0ptyIlCZXqaBIZ3FlI3h4XdGYpd7rDK27
8bwLW2VWH/U2nS7edPvCjfe/dKWk75s/57qywyOFgpIBBsiaShBDBXyR9NfZhhvAs5dzSdvxr6lx
+m8v/+PS8ZwqRxBj090MVIpFhStgo1Gu1+PO4NL/GhIuyANRDflnJKwM+kzLhO1uAuCjbqE8T06n
4iINDzBXMlnv9tZ8K3MQ4Nv/rYibRtXEhijcyog/ITUCoZQqyzgwUfS7SvXg1kVKbxml/Ss1SYJY
GHNwrIoDA048pDZj+6YB3vmdkKCg75H6vcsDbLmV5WDUaY82jg1d/yfCbQyNj3kYJCZf8Jpm/uMz
Jt3VW5SyOfcPgrFKraq0vf3HoLugp35WwlgIcoSSrM6pdJlNeMc710X2nnWU+AJnLt9NgiZiKz1S
+4mxjbzDxyW+8f6JJc/EzsCoWoyXVRZHstxaotuEeCABpXzajxLqJwBZPs2KxarQojmcaAz19Tcl
OTxHosdRkn8e42VS9ZNb1KHdLb23HdT2OYWy02FVsQe3ZV1WhPVEz6/b47Z7w9Kci/F8HYgqS84F
a96dWaD5YPoVJffoqnTx89GpJ7emgm45vzfrymxteRWkUx7wyq9gv3eHjDBhkInHD+C3wsb6xA2u
5VmA27oLgFNoXyDFCpQc64qiGLX5LlMr/A+UpxTrlEhDrXnK2veE4rnNs1qIWGuVqDCSeqyzAQAd
A859yYQPGCWSnLoqvggJWgE69Hs0YVlm8529ersdhIgCHbuQvDWIuKGpbYcoYLFFLPyC5pv6ubbC
mly8goJqL4jWjpMHBXG/2fUP0RNMJwZ8ZqPexltfI9Q5drTHgdpycu637POTUhv4QWhVwXUXnPOl
mToDL7aDHh7cwZhNSvCBNhISGgtdpFSxXfW4ePqy4+++Ora6TXRpujX3SQJMonCZqTBh3tew8UrA
CuHkFmjoX2B+hjhZb2xl/yzVXyOtdRzua9Wvlnk4vZrL7L0Gm3NYj3TZUmoOekJI+RDsKkxLv52f
XYTQiLQn69X3wDx4TUxrnYmGuWrYGTuV6zv24ljsEnh8F6qQ0Vd8sJ4QF3hP3SN5KbqMP8iXG6LI
zaknS9yD6OiROWXLBydfnaegfE2w5kTclWq5Qxz3Opbrrs44zzrdZrpNBQICv8LIJ4CJ5xU8LHc/
0rLyhtWuh8y7lxtSGblkZLp2pjCVyI3iJYfc1dkClcf1w67PmgHBRVdE/6yW+AC0QRbFWHtrU+qB
qYYXYPxeksVKyRziqTS7fbENVFxMDzjxjd9OP2OMe0i4wFhnUMW9WNXgl8z0AcdXSOKV2b2AnZHE
C70s64D1k5v7AWcBvpjqaSWcCFsabX1WBAzqZ2VJnlz6zwnqp3MgkTIz4KloX1vN7DM30FvjPoNe
Sm5FbEyt5cpBOWu62eW3GxPS95Q7TWnVGhZk7KMQ14lkJmEtB3LPPCGKmSOMqLAx/1r0aux7WBia
2ZFQSI6dOQJTOWE7luRC4O4qidKv3pkhy7OA/YJh1h8w6beAnPcDlX6okbWECDxcDXNUXK60OJXt
g2ZRxb/Sdi2N3h7+LK4ub67jcu9Z3BItXZ6GflRwLF7dRIX1KLVaP05jFEl+mw/3jcBMJZTBUbMf
LrJkWJzFJA8OLJ4F870rRSpFitxIV7Y4uTXfYoYSFRRULxBzFEWoMkcTjz6HNFQm4ALJlnD/p+dn
lvF1BqGlgj6WvmzzZz3DdlkgmryJujLeJgAssVVu3f20tiUJYNyGyaJ1kdQ55uw9DYu7MkUnBRtL
LQ15CQoRZPorSLnhuURMrVRSqUgPDiju1EgmgK0KXXYDcD08C7MtSM7LmAMd1n1iUWissQUKGC11
9mJYfvq+Fy/ngkSfpse+Yy2s4hmFjiDbXdpXD7DzEKlyJfe5625Bj8GZcY1h33lC+GwgPBNN9kig
r4iygnAirWdEYVHW2l5KsKwQF6p9NF687tBKLOGpbYtsygBfYGEzpOERe5R4cEhltcuA3MijH2TV
Cx3DRHn7k2JoH3U1VHpYAHThL4HmJ/klFO+VKjeB+KFn2TyUstIsYpSDawPKpjgotxaOi09JvHcs
6tOko4+eCBtR5/YFyZ4ebVOFW5Vt8Cl0YqxJ9sQ6XlZAfjDM0Lzpgm9J7oEF/4r69SNUVaeM9arF
DUvZBQv+LsM0i+d5CkCigZQvQNtTGKVVlbsLllrk1Fy0DcOsY1MrgKtX4vzDPLfB4W+DVYZoSN/e
UZn2tNWmJieEL0kWvtr6qSnE8y7/+oL2VcTWUEZzpI8zxfXH+5/Gt9A3F99AtdO0a/YidQKi675e
AxR/A+35RlAgm/nj9YJkE3uJD7N8zXqeTcZLf+1Y47RwVT6zeHn+CPK/NrMQhbP32gwtTXhDV+Yb
ycHcWeShfUSCgQtPNSYyjgD8ikHLk1C+MSx9a+s4F8G8mezJxl5RpqrsnF5hvEPZtyk2Mm6pb8QU
Zf0pheqe6jZgMLygK3yx9Uh+9Zc3pFgJ6bB1XS4XwiP+w/mv8niePQPst+7AXqoANh+I5TBa+bFD
E2xHk81zfiBQVHhnRpJtNTjb1oxVUVCCGaX8XsowAQQ8CEa6PWDLqrl+dL+1ZD+5mSxIzeJ8JMwm
JpIAc4SM0fZ8a2NVnPCI1BV5vJ1vTQ51pr1CSCeJyHJ4NTgSPaT2ItXZYL/wgRJ5BaZ5SWlDv9d5
tTtQsf2GwIZv3b9TCuvvsUekZgusMLuA2Du4qRFXy7sHuWTH9rIoVzEv3orzLpyh7Ffa4E7fmKK5
uaI/+XpLXVaLRBlgwX0Ovm1efPVnJTiFgX1d/j24CXKNqTzFczs3xlc+PXka3LgFg7CLTF/+lnSo
3twZy5HAMzUsPOws+8xQg/oyMD+jifurSNHUGEVsRAkoAzFpqVSFbmdQDrackLVHVPOaLFqnVodc
aqacXoT+PNvX/uhdyQLojVWICmWJIq2mV+eWDiWyCHWisbTcszGUz7u17RrFhCMDn9zE4kICJQan
8j3FoLm/KrJRxEvCiMCWbP6cSJhBn3LlZxOFl5S2pbcgUEpKY7bAU7p3CS5bLECl2WoLO32Qq0pX
2XjcfEOVbdfSb7o0KN9H3TIv/Wdabwuir+ByjBIBUnGb9N9vYdrr1SPkg4ffuYxwRJeE/ejuzLlr
VVc7w59S0xOcwAzvhinAwbXmgnwvNeMmnNdICxYudIOuOpHMrJc3ippkK0tB2Fxkx55fPT58Evew
rzNHdOrDzkknO2Ox6iWcQcdCGMwhtjjJtJfLlU+R2yD14Ii8QnOVy01zscfXdkqqaSuOZaTixjQV
lWQq2t7ghuSu5GWPzsWtrjPokKH5Nh8VbxU5C9ULLKW4M/ewhYY4G6oua7xe5kEMXz5haPwCKTiZ
pyQIKKeNQJNVf5Wyibg5nI+l+D55MoJ28kdTm4mJuE1v7sXDfsM5msJWt5M9ZG4vT94fhPI0H9i7
12DsEOkA6nAbM6vt7TmZOwzs60AFwn99dAhsrDyXD1VzXUQQVP8aCY1UnwVKmcB8xdRhy3v8sEw0
jsfKB86vzDkv3GfGyiNEYbXpz4jDfGOaN9KSPYUhpDV8fCc+/VuBBEgUova34rohdEGtTuDoTpCW
yVFLijKdCY3ENLmuxqi5cTug2v0yDlNc9lKfMyp123TCY94CHWz5GaXGZeEThnAUwgdvebot+iiq
hf9zuLfKp0C1WzFvFaSbOfjTMXSDcAQyl+MQjmz72Tk3VWYgx8Z5DDb+OaXk/PjsMNOAzEoRcy4g
GfexnpgmHLSnKl7xfV1soa/r9a5ls7P78n978pLiM+Qp0+GiMjWLGAct8OvJKLr+L9obM9RSUpff
grZ5auxhKN6I6VTRfNOQyXG5gDU7TY4MszOxm6od1fon+jI2k41DbzJ32+shixe3fJK0nM/MKPsU
2Bt7hYue1pR/2W+lCgxj+eHKNw/WEaJ8COi9l00DsXXmeSp92Pj60bGpkWYV5l6CykB1O0ag0XKk
qlprnFrxl7vn6yJmqDOzACtVRPui27HoCC/WDcSDas9kFwrjRT85TI2L9vs5lnbrntUkGb0zbuDC
fxj0LVP90Sc7uxjg6l3M590OqI95Hm6m3jkAvOEBeUq9QTiYCt+yFXI3/v1lVlAFY+Kt58sIUA0Y
RCs+YSNZTl0A4/NG/qJbvnp4Qsh24QFDrC5QaMhohBQrspP2HEd/6rB89aVUQkkaq3l7KAML65be
cPtoKKrEp7xG9LQQvCPrdsAl1HbvSQ1wL8e+jDfT+tHvJmlf+i44UKWw+jq6sdtd8rnvOSHYuH5b
WUctVoiyaq59OuIzncopcXCQ3yyf8cpNWkOvAxZ+ZUpYZQh+ELYlee0pca9DidROPoQI1WbKv5Vg
/ZuH52ljjhPqcQf4HQl2M/onvLWa+mpHrKqCA3pATfhDCoZSnBElQkCVW8MAcBPpF0Xzrc3rTE8g
rtgkatAeJEuk/iM/NCIxjurXWzFgN9SfW2j9SQDC6KbFM5f42zix5gHX3FIqbjj3M1J3umvsGMzn
jEunTJ8wLJdmd3ZD0YQuVUP22CvufsTjFXXuGYVi/jMJ1Vps9S7Vb7IGUke+IwYe3qDHuXU5mc1q
BGtkT+PcXsNDnl4GdLxjZIQ8qn0Z7UbaCJZaU7T1m+RYqK2wXQrq4QYblskHyRKV54cBD/7mDBce
YVeYoi1aaTUNsVrN4dKbSQeYamYSykIOl79bxBoPyP4ddJ8qbycCmlRGI3WVyurv04AaPArbXBoh
B0YJWd1bV4+NAMftQhAQ4cbtrcNz/vbZ1GoPXWmOg0+CjgQu8o3vA8Hj6tFvWP1Vu2RHqQ5epPen
QlyGc2XYFmZRJi/MHYKGiQbuJUXh5wS+uGSdSaXWGwMVpC4NLmiT00mtxugwEXX/bMgHQneK6rp3
TRd3eXQRRpu8lVHHAa+ejFTpInHLZjvpcSj0avWxJ8eYDNquREf4jKgewnjSiwJNSGzR+Z1YzvAF
VL8wOP9Sb2HrFrq4WKdzZ6SHQxfG6nqS6ET0n8IeaL7UZ8zBeMaZ9xw7wAXACCDjcrAcqspFrJMz
dBeSMqjmjFUKbq5eIYooWdBmwSz3IW9LE0otYRCCLWCztfiuxikJScZvtFkGdP7rBEgf3OP3hEMS
XtbJkpfTFQckP2zDtoMhuIkgykmlBTSODviL+YDvMJseYCn3p9L131JLLaByNYO4Q9cKl6bjiiS0
UFS4C098fNgV+OC9znMeyzCC44LjU/o4eBTEdUc4//uXoYWZokkVMuuo+yvJEV/S5mCGWusetosY
I61CnNNC+b1ebXAsqNm7QPFo1664DdFa9tdAe1qxbJyc8bFcaN2ej51zvNUNa2ZyqrEYNI54BYe2
f0EwGEm4hkzqK8AYcMPIilkbdQrr/a7amXCWM2S5x55hv5J7iV5Us1XRsw6E8ee+T8vdWfxPvKCz
TyLfX+KiTlMj3SRXD21w8KViOIXyzuoEV+HZO8gTx4h0sg3lJ9KHpEKlDXFozkGT4/K8woMo/63s
bhfzrMt4FCs3b9rCBENQPehZFmYetd8VDjoX1jvzHPIagBitTAs74ZXJvKV6+cRcpHFs8YuFnI/i
hVjRQ6reh/7vII1o8WCsTEBmSHdFRWu4H7AFWXwueAh5Qak40gnYO52AF33BoQN0uW39eUY19plQ
kOWw5AJj7w1TWJEDnLI2Uyj0/gToRXaP7sXt5nmWJ7BEz/qKYp3/TGEibqQaro9Oh51Hr9sKoVty
XUCQmWGnxmWb7UQhuxScnSIPEcOVUIRPLvA7eAr3bWMIN05koqxqWo4N7nQ2NYnMyQPord8QpCV0
lxpjgsZwcJ93w3Qinf0XVd+kxtoP676HNm/oyGHAkfJtuSUIcqwvC7jhryQTK/6QokuR06VlROme
9qhVEbLVQC0ds84OBaXSZCmOJumzWPBiPFNE/ALEF9kdjHNMIAHC5LGb9JVvUo0HMTdfeHobOJqe
8GUUlbk0ZWQiYtQJuaw8nTHT8mglNIOzfOK5UgAPZXIi1Afyjovp/v2CFgvS4LRZzTyoUOrld2iJ
E0FOZ6xoIwoCi/5HkJXRA3FQm6VIWTaeli80fHrEpgeZEGW8OcuiVKV9AVe2WLYxUuFlipJ/KCoe
dB1vosILM1++T+l5j6/dEAF9wJtE1UWeP90IFHa7t2FncpWup/VQviRHWThtEVlcocVWMAZhWt8K
L4SBKhT64dTVtqH44NvX5PNAO+sJDMq6yZB87Z8d2B7PDW5S95bWH6Z83rjCiyPQ6zQGdW+dVGQU
YFCj0xpY0H3KKT/HzqGoGf8qiZW4FbsgRp4/E6oBf84ssy5CYinmIwEDsxydwL2TkmJZ4n1YV5IF
8DWMNduO6CdDOS19VdQhVuQf2vk7riiwW8HSL8JjxO1nDHKpPAYBX/UCjon0qbKRlRpJHBnY2WvL
L5x1RhcM48LjlKLJFDZtyv4B7y0ZK8lJK3msrNtFciNZFNvGX2g5UtQn7IqZm/Q3jbLeLVh8KuMI
reMpGF+GWMmCPILCbbDHZbZmnj+rZbgzgVlPRvFarTpg8mk39cRC6sxftJY/EDT9Xs9b/0fb3M3R
rccxWCDvOzcnFEjB9vYQRPBnM8egY5ZvKpYMUYsYnwMEQHQbOTnY1IovcWuBKyGzFDn6P+bIxu8D
Jxt46ZQTtttjQBc9by8nwauIe5+7YtK2F6vjbDuFVcHNaz6QZkiDj67GcWcbDOJ9+H/43J4euWF9
XyQmqNiGHr0qpWfu9BSF01jof+TUcr+cafp6ET6Z2IfHbLRMw+lLUoxUDNPHPJscbVEDVGVWk8Vl
atqtXlAb64LYrdiXN9QNY0nJsz+bU0BzC0Z1+lrlHQTxDrtk0GiSmf6RjTlz3511zW3iB40C24GB
Kd5p0eQ+0PBMj+4PD54/collcMgIE3UhS/0RepvpJgKjMSKf/95nCxoUDKYWRypkBIEsjKiMEz6D
5Vi4uV3SKZyXw4Q3mh3ecxu8h89Uim38Ioxe5LotZ2zAG/VcPcTssqf8+AAEevn+UeFd/zZgCxyu
22ZwgTsxGW0lLfG7YTFAh4VgLrWbKjUEFooqe8Hk1YeOz7MDhEmSQ/bvYvteUAPub/10oUyJst8a
QL59VliMSPAuIxMrRwjiHaG95tRxZamWS1C8qj4YDLjVGmILp9MY3gySCaQKwF7oo9cLi+n4Q52B
ZDYVPa7OEs/F1zN7OE7DDaZd2Zl2RuKET3OpAxyHPuN+v2kklBckREqFHPN15qhQdUwa+b3T0rxw
0Eu81JYWTARHj/aGAniKzt+v5TYGfq64HeV9wIpd73bnW2IOf/XKw3YxYGkR8S9V5RJNsy6k7aSc
BaUV/zJBgQUVVZwRotNpT9+gI2PsovzjQM3kPnAjdZvwrMv/08Ey50n+KvhaSuxX7PQaAFuU7VEX
4IGLeuvvYYvCDI4mOz8XXiaNXZmBR0bPTRZcFJmHKzMWDNTHi5JRHYYaYGEOo76LfxOkEJpSBLkg
4V+QkxXHCbX4WlZC1F7xc6nInAcd1HGuceMsc8e4XW16wjq98y4ulLe47wyqQkMTjo2z+pK3NXMt
g9oMOBq4YBY61sdo+WnHEJ3oqAkcFzdmftShWN/GA7yZbM6SPp5CGaDq6cNYECTI7XyX5VBqb6Ee
Sl37ovQAWQKvJDThFzjE/tZg3PIyvW/pfLYvi8FFs0l8Z6e/yoz53FoRDzGUca3s3tSCZPBaRKwS
qkMwTs2NVOhf4BVvQDT5UgBkKp9QZniGprIQ7W/zdBxsSPdGX1CnWMwCFmblWnyPikw5VeldePua
b6tWCEsELgA35TI6EAoKLlqmjdsuC9kEmv2xwF08vZwUts0J0DSvWj6+hTWRgYLSuYcShvMz5ste
zEGR5cM19c/J1a8fJ+oEtjiNf9CvNe/65aohsQIet+buJj8GNDY/PjdYuN/BQP8piT4lQ/2HFma+
Vnth/YJybE5GRCoI8YbqYyVJ5sV/YW1kaPT5LJWbJ7dEHoaS+XoYZEH3EEccdvrfhXYdEq2TTKdZ
s2vjUM2jJwOmIvuoXlXDPVdDo7LKa0XvY2lse92oLYfOpjmDZxpzhbWTqYXNRR3Z36JO/QLAzarW
Pt3JUmbPevaTRY5SwaS/LT51EKPwzjnfqMO1wZw7LTcjcEWhyoPPAjp/TqxF+2LGa3iGEBXYx46m
1RAFz3f2e5fNCgEieUjTjdNcLsIrznsifj5X5YnbANryeDpLpNlMD8bdLamthjG0uVWMrTa5DjbY
DxE98rJfXvniyFG+/zZMDEy7/wpz1lcCURvbknqy/ub7FQdmNeK8i9WDK96/A/VTTjmExM5IYwZj
BcKlg5yQHadCQWumeoPAc4VBVRR/bi1e45lRcjLFTZ1U8VhOhXGtm10rToia3Lr/FBRfapoZhZP2
tWTUQofWH9eWhTaBYgPzkwjnt0CjzQMJmnJkdKo776I+UfaZL6NpHDsmiAUPQ5yB7fL7GfaRqaEE
hBg4GM38FgPDTigyijnbz5PmHdg+NiY0vyJaNBpRGvJ9WgixChWi8mte7snpajmYS04wsjWDzzwz
QRtfGzH/8atr7Kt8HwiaZks84Zi75mAelP5hJ7r66gJ4uCf7ym5Nea4OHz5Ol9d63AB+DO1QGBaL
noekEw4DuFmZhCxJIeWz6P/CdCcwr7BonWauvtOYDi59IMyNONsWIuZdJVcLIaSlTflN7WKho861
lb4gXq0Bkw63xpC54JRe0P8BsCsAKkYrjGgetn9FT96z3yT7b955MFrWaUfcQjgP/h/OEas5fEum
/WTJlXq/e29GHmpxUkMaR8kxRYgCJdrKdqmIIZACkLirjaOof3huFC6xQ0ieq/eqShZTqYDCbN9X
WWfShCrev9HAqu5o5468OU/B7G7OiBtLpfk6+BTKgxGINu1XwVch7gUxV6jUVyugcbrAqzX3M4uO
3k+qbK3GHl4s7jtkvG6/IfgxwqnO4kfCglo/Lh8Ou/crXEMA5BFBfhoThTNqAeATaEJMtjMTIwE5
2vOmxp6aBxUQ8YQ8QZsbU8FktVldPkWkmtun0oWxnxisBCeVJcl/6Q00Vm3EvUvpHo2jeteDCqtT
N0wsIFoLXYwwQKB5akwxVAn8qTcnFAzfbRKdTsYuIPlo91YupRRBPCOGAjCCUsuPzrXXtNSB7m1U
L9OBfsNT7O9vBKOCIrc/WWkI+BJMndWmvORA8FZsk8v8JcHhbHdUqLDu5PEWnQ+ikyCjDpoOnvT5
Y9cHdh6L6NaytSFxwgIgf1beFCIhNIhxFC2GHTVJTx6VLPti6VwjSn34448dOXTveis2HTAYYm9p
y7bh18InWR/2J2ioJUJdglRXWg7HVQPLMSQGpjK/bngkDv3eUc+3pQSRfwHYRED28c5L6YWz1Dc8
qwdqI5qA0vPNNRqQ49VzBMfmRhNZ48oPybQ+blccuC9BCa4LiMptHPA9j4jajf0cPV04EHjaY28M
TYa2aANZklZw+0PBmOac5c7BMwJBj3wh53PV2Z+HMEpQ5cl5XudN857GN2liRWaWJ4Vtz32jyc/K
4ppQN3Oi24yzy6aDTQK7IxiGlpQdrb9qrSPvzboNzHqYY6GWPFrZmQxVVO0otNAQDPS1ef0eBxXD
N3NHzyh2NCkgmKSC8wiiXytj5+mF0/zaEL2BfGW5BeoL2derNRmuutBEqC3XSiXsBJGQvBMQtIew
ap2bteV3wphcsJRxtYvBGpBvJbvB0g3I8gfNsgEgWAGJTnpfq/mMVcVDbIZVQUg1Mf7MtD51MDyS
iIE3zXpB8r9TsVSPeKuaguGpxgwkKsEJyXvwxM6XpCHxaQEQ+Hn12njs1+4QTyIgigDGtH3Niwz2
7pFDBglj9ILYinZZj5lzcbZY6Ntiyad3oVpNp1BIwcLoIKdJAdLQ78pMRwkwTROGVKEGPs5Fx6KW
hzHLGA5x9jVaJ3AYfGMuebcstIjKIoWdZGaZND4Me8FK0y3Zhim6P9RtwtDjphgfnAl2UrTCuHlJ
qhFzoWOxULoRgTOuUoR9zGu/fop/b/Q8OENg+bNzYyfcHCeO0IBdeV1GSrsnwlncQWZ/Ezr95b7f
1msv7K72+kV07VQIpk7NfIl5FcfSCAzKKODp3cK4i9DLdsvjieO5w7YaGStDY/yQdhv/jS2hyl4S
/vjJZ5S/1fDPQKKTmsmi+3iLrngmti9XvNRWLauiFSpBxhu22iw9pPGBNiiNm6W/T5XwCyiRNlJM
W7z8bt/w9Tcmpy+B0ieotbiiqWmSsbiNzceapjsPahSxBHDa7AE43vaFOIRMqnVKGAdHuJ1It20g
rzZxg867BTWVlMS0JkPKGBF06CIkWBg1AeudYAuNd9iDzA9DqAJuu9an7dviQssg0eINIvFTHDnD
l8X3ZX99OJaQ/OR8LmicdR6VdPjcesD7InhOQP4fH32AaJoxHD33strbHaeJy3bUVBpcLH2Exb/O
M0eUAKKw8KMh8f0FozU8YL6SNn+j9wRhMvDbgSUIcT1sYbl/nAf9MgbAlSyvl8ZyaXpI7C0ZQ6rw
kTplDADrv0wV4IL09jgOIcp0lo/gwr7XCeYcy2ngxgoNSC1nL0L7a3gdoRZ4Z64SuH05wa7bsprg
BldXR4m2olq1G+3X/s54a4v95cGlnOlo1mg0MHoHww39scgImKx2F8dLEgCgoxQB3VZoI2sVlCKI
U2o1OEG0gR8DRZRVQ2ByxlhswNOe18Zd6/jN2V5qD0X4xv/C3VVzvLbDgat4Xq/NmCbJlJvNKmxy
J1f6pTTayFyK80QbYnWwqZLrtFO+Mwr6faf8o26KseXEEkvjdwYPfV4T5BN0plkmpf8Q6STzjCtq
Z/9PgbFNGQ0a7AqFlVwDbRF+BqctNMJ48MmzcYWNNnJK8xX6JQlwHvJHRO+a2RVw4IE08ueSDAr0
gPKjopteLQajOr66gh4jqDs4PDtVgScb/0Ee7YQYGhdiDIPMRLGg6f06xtfM7ij9LcUAJhBoOxDD
/zPEvONgamHR8akwnRbyvTOVjPPxiUvziuOKw+OwU1N5ByqmPHbz3Ygr9MVYAncYThPmSEN9kh2I
EQdSDUonYMbURbigpRRmCTETvuJcqg5Gvabz8IFW9PdC9eS8gbnpFwHHZ0JZt2+47m/n9Gz4RGZX
K21yYeeAqVvTLLUu65ei70WcrRIcLpjlWdclh+DvNiR6suegjGV2LGVBtvfQjZiabCyqmE4N7kNL
qGtjBJZCLj83WV89JoDIbATT/Ufrja5mOxj1qHylTrKx4Bn6E8exXs0BAgo9A4wDbmuAIg14pI6U
dOJtxPkVQvsEQKFyS+PdI/MTaA3o+bUSjMCxzGU3JEqRTN1nNTlmi8U/2CYS5GHxDLHrcxDiIdgo
t+pRL+fuk9Ne7aIUNyMAoSglp812CNfWEyOOSUIQgFZoxACfYi1QQxylzYWksjLDx9W8WpYc5iHv
gYJ6vUvigGIRh/7lSg/cVNFGfhzM0N6hsrMnnCIyMwo1IKjzeLFYbGZmzqzRCxSzaSMdE5VaSoD6
hRGPmkCiSs3whgXV2BEKuEy5QkSD8R8Nd8YIOlp+1fOvNcO+ZopUEA070ADzKz1clBkkpB4sWWec
613XYYbvabNDUgpTFcOoc5llEGqwaUT9zZiwwFlKjGnbBgt7dhatYiDZw3SeJxgIJ4SanTi+9LHi
5xV2/3BgQgDv2EexPs/XYRa6Q7EYdnSgvDpc98eon8o5wvZLR5M8bujWL/Wm7n57ijgeLr7kPqYe
c756v3DOB+iwLNoQ6IkFCpqUNYdGeVy5lsyNjvrnVMuGvjQg/vevo8pzJQruxEHotQfxGTefWtV1
vnuJjSVfM0Pk9bnm095jNOJF8c5De65IgGpXhI5wLXnuPtlmVOvJg+mRe4sdtHLzpTPgavPjCG4i
aIhCvZ/t4I7idxkTM6HLniIp8pd/v/djDj3/J6xpTDUHe3FxePDO9FGKCcuNz5jj4Ure+vUid+KB
JEIq/xNZkPmBOthdRUPpbr2dYlRgmcHZqqncYwnz82kI1OB22C0+NOmUHKnojgMYpDDU8YFmYRsW
TJwg26DWYEKeacsjkr9lqoxNRbMZIGLtG4fWQnaCgdd+WdFnJ+ZBa8dLo54rNHyCVlAVgBLKyVNj
MZtm+S2LX28snWQRGo5ynt3XgocSAHOLfaem4ro2RYjwduZ9TajSyVsaWoHgqUbfI/Fv0hpa3YAe
e4+mbaaKm+qTBdia2/KjyPfNni//KYTPK4QTYDQ2CoPF40y3bRX3N3Mtfl/y+GJCI4KHKLGeZBvM
Lqv3+BslcrV+Ki0oroRfYd8JN6a+hSL7/93//Uc35/e60vV/dhA1vgYhhcnti+O9SfEJPxXitPNq
QXjOu7RZMmDb64dCGCNqKaOfC1ZNum1Od2kqMWDI4EjwG2nob0/amEc35qqa90KfkqoBXyBfWYYJ
JEVF0aAbCky+o0BpBTc8UiEaXt+Dts0sk8XMrVgnp/kqkXEuGpTCtto6giSemaxrGkxF0SGu6bhF
4tfsJ4/8+axW77tYPAVbIdnLn5hMi8lfLE3wKOVcOZ99BVVOKIJg7KzGFWLOfeO/f9Jbp7hanPwI
YERpSYRFlEznFqRnsDS71NlVVMZvJoR5b34SL3LQh34VdUxnp6FyrIIFBicGRmsnYGdL77zkKPRM
/rBq+Oj5GhU1T44kX4W+qHFAzCoAG4G8/FYmMnWE6jT/x/sTH6cm67trJC3DXQ6Ja9DcZesTJnYl
Sp+cca75j98TdpoEAOAd6k9bn40jNWGa4gONSJB0pv1jOEVjARLtlW0efLMauqUOznFAOQdfQiAS
0zmRW4rP1+LxDqAYSsZIJ815wH2SNMTTtcxq4rbFZCd1ZRfBVdviM6C2wC8LmftNmZViODuhKpMi
4ufjtt6KOUkhcZUHdgoep3AGbA3xWbZj6K3LvBMVbhSNJS5jGKj1d56tUY5otK/DX9LfWWa7FQv9
fnJJEJg1JmbGBjQ53dKTPmY3+ez9zGUL4RZ+u9uZR6/PKkububcjfP7T9/1DG8oT9Ya18l4dhWK4
I3MsQrOkzy+QQvsWI+pFs/Gzlxpsvly2CnRmxHBEu+Pxi3y+wU9gToCUcjJawioBGdzcdooxDQpX
BGFD8z1j4mw7N4OOcdp1QzlG3UAi+dlSPQE9874C7hL9E36yasbTn0cSZlAmlXRbzH0y58Sjry6G
k9Qn4NGOOCevSSemfiOQgt9NqZCnaLOTKsteB5Fo0iGKU1Wm7o9gEmwzDjsO88U1MrB+Sx/5EhLm
wBx2v/MBhh2JC+RqyLnPF5l4nryUSVkyhhNILbWdSkA0BfmxwgrxN94Vl6r7OGEPNfs9IUA68Iko
mYIpjHQLXrSePzPNHCp4Rw+HoWxgTjykw6oyFFwwjpSBykOjssoQLr9wHc1DSwlXfsCWVRuLfdDj
A4rEo4H98cLoayujZHPBRWOBYmoqrkhyywP9y4b5RjlszrNF1npgb9iyoSgPMdvf85WdhsULXHD3
Ejar/Wzx+PKtaxPjRku5XsJEdtF1+TZWwKVpNia9EWPhO4zegHdM00SBO8Qvu4rZWX1igB73oP07
ZJWbELCl0YvRzhIrdwpU3Q9gKlZYr4iRvdTQWfpuLDluy9N5fdZj6jE/BAAr2YOOnNVDzKmA4MNK
gzzUQKHXYyDTFQLIEKtGRjMObHaSJaPPuTbg4Dkf/nWs3VCiQyM3QR247qMeOCttNByEv+jqLfpG
IlK8YT9LSUDo6pXCOTL+NqjTinSmw/weSqbiVz9AG/Sjuv+VFi5TB5n45CY/yZVfdDeBh4d9ZIcR
JowSksHwJNd9umxLRKYpfdblULmgoazsrbcSV+wyhXXDfgtXknjtDP3C8VYt01DOi3KinfGIZ4wS
qc8Vr0fYhZJlIESGeJ8ZSg1R/gsIQLfLONEaIX1NIaWw5XWuuNj0T+CPQFDAGZgB3CJ+0KtTOjdO
Nyxc3wKLbirBVC7tYf4N0ZayO0X3t09G2YebMbHWi9x99b5lQhqjBVnWzHDJGPFbgZm4qIa8KR3p
yxVpTVFKfwxqNWA7GWdF7fJ76IbbHv6JhpFwzbMQ4l68wxoZLdsAm31lffi6IMXVncJW8hn3wrM0
eSEQuPmo4ZF4S8gnFIpXSD5bes7ghuZ4Zn4fME8NpLn56FWvb3B0gafNRmFcZ3c7Q49hDUuGdfNX
0dOtWe7PotG6q5UsnKYI88zz8XfTXbgyommLCaj3G0oLUZtwA49HYbG2N6olWxDzMy8wtt1W11fN
xCh3I66Bl0YOpEMaK1kTYQVp/FF+tHM/oB9CfXyCV0mMcILPgr8KdDpuN2fQvSKXp+BRyooEwpQ0
XxvPIoHmK1wvC1EHI7Hx4ssqyZKQ0YFq69MmRqUXBa2xxpCP1sYh8BSlk7UvpQWBapE2XCRCwVIh
9+UDZszwq1ED6fZnOTtr0vbxeNQZhgpChVWKGEGdcbcHboiqY4md7fcMyrCrgSE8gJFHJWZ74EM8
ThxnjrpvGzBAj3FDtsV2crrFzne26oAj2DqyyIXXGgft58W1/OTGYOjz1h9D6wecZRfuzzTYnjcg
58S1OOBcLgLDJnj71fNI7m3ZD+Qls6Uy9XeeqKoPUC5ljL7q40fl/E+DU+p/gBzisDitA1Ji+wP6
zwCkHHM+VDeSS1fy9a1VdXTeEKmza+u3MjFXkSuQx67tZ8YTPIHJwvwgcUsqRgjvq1nbUZo+9F/Y
xjM+Waagu/CKBTZoqGtWiVJ3/TAuolJ/ixYMwIee2alzCKSpxQO42T0NY/KhSRg3NmhX9Jo/gWf8
AM65hdgZBRBUeQENrIZtS3FngWKePVWqXIYxCw2XQc0Pjtr6vLUP0RtrWi+U/Whl9qAfZJNWm5UG
JOjhoIzV/UaIhQDcSHtTYyrZE1LNUlEm5P0vBuGHxDsenm5qvPH1HUNkJcSpaIHPNrrT7IePuadU
CuB/IC83W2EjAD6dlkk4KQv74Xn3eU1u8N+FwILJ+aK+ZCx9VQWVa8gjLT/KXhrG+Us/psIkbikJ
d1mEiBCU3nQD3MtnGspMdMtzwctZ+BWFpX8EjneYdrvj2LI6OBb5Ig5QurntMNujiErZYbhN3k5x
z61IepiwKJFOLMu/3EiiRU8582pFIwCupZC5JPfrBiB2pJ8VbH2Oo+oDJn7xTe9yiKtXD29LE5dE
W4LDEgoGDW26l++IdTnXSq/Er6RAOIIYUFutJ52s4omWBx9TPB7hcfl2EJE7mEmxBPtMhQCe2IBZ
hj0QWg4m/evE9pRQfcQmT/VQUy71ecvAk68K07aXmhcqAKz/ENUSzbmReihETNXcgDpuBmIfH1oG
vfZTFPeLHsgRYQ9UTdSyM6nQyoBZszgKOLg6B6VqIVo4fonI0zVoZV+HxYofpPFSLFj9D4qZIEqX
OnZru/Ds+WvpGehn+Wba2TYxlvNohT9OAhd1sOUnlGmPIGC8VUR8rO6xTArJfdMNd7/yUAbkmjEu
zM6iC5PL6F5Fj43M0KVLKVp0kenr/NL4azVoWvScSiNvULnOgOq0dEeidaN3mPgquq01zQLwmDxD
SkuaoDYFDHt5+9o0gETBGfnxObvnFouWQZ/XfMvQ/0hhVbuA6u+aLrqdvBHn86N7LW0hWupl2qur
ieh5qzH9KPQJno/GdxtuUIi70CDjVgqpvyFM5s40Z6j9n8bqucBUI5ryfhFUbqrEVGwalgHa+PNz
J2K6aPX2DvZZPBIks048fnU6l782dMiHyQ2uQgDaiMrhCnDNWf4eBCpDCqQhAxNmb3FADuEwY1yX
mj/JM3PG06tnB9BV2UlhscQ5ZPebjvy5zX71O2CECQDa9Qwodiz5mQ0ZP7czYRjgSJPCJYQcZjFF
ldzeikyKRAJX1Kq8PW8CLxspF7AqLVfgiVchILXWzO3Ce1o8ZDj45QbgoKHHyMl1IvxCsPxN0kir
Ib9gEImCDdMzCJAhTEkozkSbWxWRKcVg/OX+17P1NgcWLCvARB7p5SYK0aNZJYGe/KVVYUm8Sp5Y
Q1wPO4kq/fC8k2ne/qEIvow8J0+e/K+CsfFhKCuQqXp94c/yFrknc98/clWhEHQYxyzDk4jpwBdR
UsvNC11s+DJ1M9ZJVaNJjWMHAB2jqKEPXmalWesWXYcO8qA4VWMRqWIbmWFf7tv3lX96v3VP4h+p
Oi55I5XCCHUODKOidxDHRZsEnp0LrPPqhraTdS0TqhWFXKaFYfRSj8Rs+bg2slRuH2Obv0hjCSiY
xTIpdY9Xw6QYe1UocSjmO6Pc0W31m8EW2hovoF6opELb60JhleVtGsHiQKsgRFJYuydhklWdC1xG
/4mZjk/+9M7OGmzFhWajBQTHf9kS34jN3aYRZkW0I515+4X/X2Ox9DQ1R1v3jj50dGQ6hzD2o6UW
dEP+j9sGz8Hw9nJqfsaneX0I3jpUwWnFbXEU6YlioF956I7HJcj/be2sUkyxWv81ZPadS5qNvQeL
spqPCMEQPK8/hxy07cYUgjUu/A83wzDMc7SOxNNBA//AK4jBzY9nfEyiXcz3xGxlkB/Wzk6MxMBh
voSKDnEXiF1wA6aD/idYpiSsvrikLra2OvQnw222E6qyjz1lY1YoTRvqqDZG7me/ipVS3NVX1t03
FQXNnmzIVZceOPgEKjIcGPTXUcLIJfpGjrcJlamCxE2G9RayzJJZFNKKQT72bDWCza/USTm+Iww0
6UGyz4osHzPlZ4HtfWbdVIT/jiVNRWiZJS9mAN/tIkaJKeTCNq9z45RMdolmNpBPFcevxp/Tu7CR
4b1dJn1aA+36bbc0lyjgLlLcSoYIJzwQh6lIul3wlWXt0BCbcMmXH+MILRmLCGDCi12LpTEWpC9V
0pDNkn7ev1sSjuSJM6HWZNTfwM8sZbOfflBxvj2dAl6f40vR7GlVtVFULho2UBDDoQVHXdEEA5Fk
H7hsiFvBnDoKh7fzDPvwYr8cq8w2UyMADZs8kOGodzhUvJf9TpU3QN283MPY7HiMUkfGJaSWzZZ+
yMBmtZj8MK5LrGvdYXizA9ldqRgPGBhQhfs58egbfgOM/k8JbZKPAnW+BABMSifE6HX8zTUi2oIH
OxcBDWSkMMcqO7XjkFc6e5qJg9etEWWppteqY7uM40ubk2DoxHxVWK9QhTV8k8CQ+5m3Lu3iTNJu
33rHqXrCstzbzAiiB0/9yq5BVJ6J/Qfy/Amzx4BF52ti3MpooDh+Nu7hYauvQGzCUwoI7yOFZ5M/
A1WaN9Jf4wkReoTxzIH4h2+acRlUUyapB1wFyY8UDoitrTSOybTqQ3eVtePtG/oTGpza46LXqmPr
njqsI9acc/ziyQuvrcZ/Cyur0x+3rR7DfJ8FAFfMrfoXHP9NFAUn+v1D3JrQ5ExQzE3BIXy/Va1S
fVy23aF4312b/GTQLGm8CVTqqzUfw+1XNMArGXa1pw3zd8Dg+lwdI+QsWLCuBc/bqkKUDVhfjJQY
Ju5QJfw9puf/+VPDF8NJB1QOrtQ1/kMdp93N/E82AziUA/TAMc7jvi/4YR5sJHlYNcNdYm3eVUaC
0lFe0YWUb8SLNvtgRHTeTaC2gyzm75Y4VLk+PMiagHFdcYYk/+cZJYygPvFTJo94yUJJCYPg7KVh
P3OHVvWRFe3yxKSBl2lQofJynlARkm9T6NSBMiWe5Of0THaXkiKwmQ/uOStRRW2W/AONcVNJT9SR
rO1TQjgdGDA6wBlsSXOs0Njw0m5619mLqbhNgBL2gZniHCSzUp2wKmFxW9jrTDlFBGIzC28IILXR
5yUum9oERdqWpt04Rhg8y2I7A2neZrxbMS4gP/C8ned5ic9fILb6Nd//eZA+ZT3Dm1VoXLQftE2a
WwdMknHDeY7dlECeCEdadkmvZ2XZgazRUPgh+iJ3ZwjmVETfG8kprEgx172hAUOgJCk0v0KLA8C+
KJKhWhTFvJ5TO56dG5QGsad57G8a3BYeWx1Lu7KbLSxMF4JmHycO29JPyg9XoOeySkO+IDDf0ki2
i+S2pIP1F/poz+45ziB3nFJvcfyAhlbAUQiOg6QAfpPkkrrwrhklCKFFxaJThsCK8Bd3ewXZbxvu
S8XmL1jAPUE3JOS6nzZYmZ9soLyS9O1HDhT1rZQnJ2ExRJ825J/kERTMi+FcVhvaPPr4jHlOVNNJ
kYwBc9iyciqYA998PVMfekYgNpsKCh7I9CBDrdWX1CyDZGUMYHK58hzPRcEh3PtyHoWB7aZKad++
QcAbKtyIYbyQdNsobRaoJKhS94CTKD7W1vQ/p+n2nDKqg0UaZZcH0/2Z9aE9J/iLhJE1UswBsEZ+
nns6tS8jMe5QKunDUD3vMIpKCHQo49EbEFXiZFk80iFH01c9LySBlb2iADaFAG+lqU2IEQQAfIlI
lWqF6xFtDKGXRl8y5AK8t0dnKHQBLlpAtD4wwqcrDtATwbc0MH+f891YDM2LNkdkO6jt9HxNgJVy
W3tUQ0XVUpZPIha8c0t+MDBroN/M76WWAmpZucUg5JeTEwFYTyTcs2czPn3rbeSnzTy8Gfr4hSje
XU4LBhDP4RR0Nv3L6NBm1d9cs4ZYWzcJNJSBZGdgc7CW0Uy93pqS1p4x1bWFmaA8pxTOHG1ggWA5
x545pmKDsoq3N/xqdwgWGeNt6Eu6JX+uAnO9NgZAnrzS5PXXvGfDNLSoZ+vcdbXV6KQlxOCGbr4E
J9Y5jEXAnOKnXSDshjmYAV1PbnArFlziMSo6gNqmEuIRhJXqVGb7wwH7SC5PCtlVbHanELRA0uio
KuIpVCONs4cfVgX/396Y38LWpi4zuOfaB110jLbeiGennqYHZgO0pY8gHcT2MC/UW3vxM9CEvRNu
6YsO2wrjngbE8eTFEEsDnRLnu1C6FfSolg0/mVd0dp52h2pBqUFvG5tFuQTs3VNLDW9Y1yTn8IYu
HK1WZZrz2PvUNZOfVFIuqQ3gQx8BahiRBENsyjHCjcBKWB2fwkJkjKrYfKb9vqNn6ZZpN6HPpNns
jthrMinDxOvXQR5sIybgt6LSfYyV5fpp5+s6G1axjsYJ2ybQD8/KZIgirO8DYRebNTT01LS1puRv
SFXV/TFbefJnlTHsvP1TMm6ZTKAHYCZ/m+HJIZlQCM+P9d53XTqgyQbZeJhIE0pUrc5mNpfaK+rN
p9dMZPiEwVvyYFq7bpXDECSympDfHVbhb8zQUwVy1Y+Z3nF4RLkACLAVb7nUn0IdmptcM8b4J1Tx
c1cCxlmlyKTFg1gIqykVWWCGJUyQxA384G/2Rk7oHbUJWUnsjkNXdLipBBhNzMXPqTjDzdxBLTRn
pmzZkIsTlXbcet35NALNQerPolPsH8f9HM7fmXNsRGBdNPCNmoXvCeUPgf9FSvTxAPRAD88Vaiq2
vKCr3RPSyR0S14nciUoX2VFM2n8WKjUBJZSQyaYf16vrkr8URpkv47YrxzrPpaI+fDmRIzg6O5uV
t6/MGSWnCeYEALNXDlnAe1eo0Na2L7bcPIKunOHrR0JMAZEyhGE7t+qQCzps6WbeGV+gr2y4R9RN
KTIKWPrdA8VWnVvhuT3UQd5zglzOk4N8Gcytnm1WbnYKg+zORCh+z4EubPvcZUhmmUFIAsypWO3Y
wYmNF6adv+kw5aDp74IKs1bf3Z4kILHbgUFKvWCILJpRypQVA5VlsJZhvNrpshoVPBOjM9RsMP73
+jy/ch8D9go+pxPG/ZfqqlWteV4HZSXaF/thkSyHIQ0K/jIuhBLTbdf/SZTQNrQ8qhVevNemxe5D
0HAp6OvsnBLTo6S54TwuRUQ9UXm802U0mNyuQWVAiZHRTAMmrrJ4luGpXli+gjoMJzvRCfKNOduB
sbs0hf2dXrZHyDcBZjhTY07w9IaG2HZ1MwDlocHxQm4Zp7YhJ+KE0E5Cf2nl2tL4LBrJ8UJo0loe
bQTr6EyWJRoi+3zPz29IXK0P/rvCjIugXBigZbzmqVt3dcjQhOefYR+n/C/QTNw6Lj/Wagl2HMMZ
yj9ooYNozwTDfgg3kOSfL7lfarGJq4uiW5Rx9Ndwcct1BaRss0S9wVUIEvde+pduA+IKKH6j4iyw
q2ziNSGnQ9yEOPs9JNWCCbH6WECXYyFEuf75pgXpSdd5T1smVluA05h4dguGL5sRH1zoBJg0NsV4
C3piFz49ZQzcQoc6tA7Bil4b3+0BrjPkt18IBxUSZeHgzU6bQa68tT/UM8U6D43+B1ualJBc/xnW
qQQfAjzEBW/qEsxJEgxpsBUBGkMcB93sdUkRozlx8HNOdKaI23uDy2AjmQ7DDveI2Rl0Y0+JzVWq
K3No6mJrDqHpXCjfYwPHYgdeBnl4ZfpRBcJAy8yAiwACC2S+djwSYZ1rDPzQPQy8/M5f2zKmrEtT
IdyMLNfE1sBctO/F99Eflph6EyYqeAX8fB+y5oNiR1MFSO/kTHqytRMZcJolun4oH1uMVsVdT3mE
7ndpbTOA90FA7sPPAXWPR1iEJ4G1WnBFUOesTbt4M1b/jExun6rEBPKmFp0GdyX7gR/s3/C2jNhE
brw/LHE2Keyb3gQuUk021Dqs+K6CxoypOJXEFoWPJaaNj1sngfM6ZulsfbtKOp5SZ9cFj86jQ/J3
gccquJjzDZS4u7uytZHRTxUeEzVlvnGRm4tjlB126dlOYdj3HU2BSSRZYxq3kvd0TVJhbEw9bFx1
+CFrzjIqF6Ygjn2w5nF7nFL5T7faQAeEXS/q4wYP6Msns60kW+1TAIRiWXLl6S4hkAF6aDx6MX3/
zABf17JKFEFIaScTLq8pzAySBQ4z1rn3inSmtvlo3o110Y0/jl5KmTEfeI5plRweoTFaYM9XRDy0
Z2cvAFFGtZtEd+NYm8UthCxZ5CqmfBFUM5iYbL5zjiPFGOKLNMRxyHagbWos1gwBrWzqbgBiUR63
XXjA860DVClcNS0w+dd7BIbRXdn8jwGJIMCqr5ZR3QXLdnzihLP2SYaMLcteeVd8RFO+38luj/TF
plngApRLOo24Jp1cEjFz5OaMbpc/yzuz73yOn4TqnKa33WMcqe/2kCFw5E09awxB4fG1KJ64Zu2k
H3/ciMGx632PBwhuMvWCiQGtDQyWuAFgjyEdCmo4EM0+LuEU8/lB64F2Ii64tZD6LG8BRuIuVpXK
iaA2WODB3tBUurEcc6XZnTIHKgJmVvU9S85qQEhfTe+G+Fu7hssF2qjJjL9YpryfkRhYFC/cn6eM
/vO2wgwGsb/tE6Y8TIo1/natA2heFLag8/eCr0pqWZSLS16KyRLQkiuaHCWeQzHMD233qANSiYnW
r59Q6b3wn05IXbuxqVAZH2RVw9/2fYuOLh3U/rkjetyxgnoM/pbzaqxcpmEmKFC042FPhbe4mr5S
AaYZRZOJecnTxH60Ppo6FeNTbQmIWQckN3p4cpyQA4pka96NAqeHUFEVCsGhHehsJG1GcBhap1Au
LU+GIuYGfE+ShL3kh4tAi2Nz5yvR2Bjva2/M7MfmFjKXdGZZD7lXmDu6N+PoYwVGOWYBJkcAhh+2
7O5TKlYiD1+xvoYbyjW+C8ZQOP96Is35WBH4rBrkbxrPXnrvGBnfmOU0pV8OZXkI50f7GEBZVETl
qPh9e8NiAKg+gPJwMzrvtKqxSwtCl1Scq0ON1aXsv5t6gHnxXrlsDKw+LAGTVx2wTsPJwt8K8HVl
oxLvVpJYGwaZCGRMBALiYh4BkqcRnnW62cmQ0HuXy5PJjbNAc6o9G+a5oX1QtusvooGzd3Q/l6S5
iONoWcBy0OFkE9k4ssCT4IfaTaAvVdMtqMmAB3VedjnkCqMPz7qv68LXF3zm9sUoQsg3m0ewa7Kl
o8/803sAH4Cp3GAeLfE8EMxD3+t17wlv+ovotlUuOhrbeHRXDOmJ0nGV0KUkKGMtwmERDuRuq9Ql
96bDY32W/Fw43S2tp2z9aG34iyJk/n0D5GugXU4BHVMLeSENCGl811aCGOxs45y/Wm8zINS1amux
YC8CJ8HVWsI+AIn17lhhEGSM34VTcw6J72PK7TZ9oYLoixXENFy00o4KqfdOu0ce+JiZP6ChUnL3
49h8QoSVXRDVFW86BgkyxcYNyWet4Hw6rpbaFy2mb6jaXUheiDtL4VRk3LYMF0sRgCcf4s93AhBO
4TWG/cOn2LSp7EOY8HXfRc7Lr3Ae5kgFMw+TXz+t0YLpvvv/n7iM05i2wpP+PIFCdpQAgC7ydLXG
zKkj6bg31O9oWpfug3u93HC1tXqaGXF3AAs/FNeKR9zLGl3++Ys+wfl6wepjIoNEENbA+7yABsKk
KW8lVXE/EiFYgIErOT7p78wYyEyo3cwmHGzt+gaTgjRgyptPAAKU23sMAea1iS7bbm0riL0uD0vz
e9PdKUhmIu7mXHAPIJyUyOGYptrhcYxOL2956WSP4e1eDXsqpXszw1kvPHB2FA5DgrcGbaBeIzFd
H9EHXx838BHrfOYY3lq/dETDGlDULUVKM5jwm1EcDCVILaISj1ogBjWveq814uFo5PBboEzk/BVN
0SiuaEyp+SBqEzC+6RPYsCyDFnn8OesUFmK5pKP3pbsachTGAUrjwIXT/9m7Zd2npAxcKPoLzn64
GKLqR7Hnd2XR43i4CcObbXqaOYv5jBKMhFWpw172ZoFy6fZscr7aBgMHOUgjYDk7R2wmZ4vuRmpT
HvnznLq/9D0UuDBvyePvC1yL9JmExZoiLpsBfUJDeyUJRogXYEiTz1CfEcnv4lcZ4/wv4mxgAFw1
nsx+2/pnf3DGAItFqcKe7VMqhzvfxipllhPvEJMnq+M2AWUBWP+qzfpZGI6q/Zz6JyIU0RzinE5m
M4Ze9aJFY9sPEWTLP9KkNnyAgbnAQ+Ue51OSxHhmvZjKoQWgYhCUJwHpbFwpJ53hhGET2DECgZXF
y11m9Xcjg4Ne0a889E6GMsbzRPdLT+tmVRFDkHcXf4CaJ4vIHQWe0wYwFoOr5RB2Pjb6/NcF7oxg
qs0HDslVTNnHcr9One3tjSxwpunaTqUHjKeLLuD/GlA6Z0SdIVQ6J6yleGaizshmXOS/bp2UCq/B
8WwYEnbhqeq2rqsm6xDFZHwr2kZXrNQnkZgroC4D2UvzAVIIalLZFCfbSu0Chq+77WtyPl9jowwi
9iX9DgldkLx6zsQQRrOqDJYkR8LLB1MERtLvMD/5utfXRHQlFPBvzWcn2iY9cHCSAafi+c8BkBtw
Tymr2alOMKMuUNY8yNBZgCS2SZBCRCTvWpDo1TkdfxTK5ihPND/H9lwLCtoaRoi5Ql/ZtL3NHPwB
3r6eH0keFpx4Wv6WkgfANm8Kh6jMcd74aoDchhzf8R085TBeK6PmzWDizvLmweIEaSxsDilOxSL+
EOSAXe8DF7X6rcKMaNbl00M2RK63Abn9SnggfYoyjcwQIUZq37MfckEyMuQ/wDlGy5jvkm3yJhH8
WOf6jl43SXj8xQqD1+ldkfSRXsKemJhhMCZk7yxO9QIf0kRERaLUxu3w/jfbuzGOn6mkIaIuzXxj
BPpzbNY6TBkwSJWBc67M7LBFpXTu1PAR4hQ2d3qPTds8LwgvvC1dFH9T0iD0+wdlEW+ck9ZZddBE
/p78qgcxoEQLA+N5b8E8jDvZ4pS8irZ+zTQy0OsRocoAChghCDBm6db30+dvM323VkobNvPKqOSs
Rb64vCo5bgQz+LdISzpcEkpOrZVeS0wa47YjTPsEkOCU0v5v1M4ggXuZLAc5dkY49FNeGCXjNUBF
vj30Hvcfh1xu8SNaM62eijN3zuWuHP1EmUIz9wXv3eUSKTOMJZzbOSZmRbV2imYfb9hdSSRnXSym
4wtdwV2/e/ob/4t2cZ8oqQHO5QS4SMSb1DHzm5p2RWzRpD4hWBqWypYtnhD93GwINZGLJ3YWvJJt
WTiir3ztqWfUxxgV2GuT7Ljmt9sXdTs777LzaiP5k+U1/5GgLG2di5sL9EgXcTLPcW22qC5Uliz0
rFfZuL1guPOVar1yZ9pLp72hdEdZV3MudfZ4skuD4P7uepuOhNyi2zktxrMsYxIzfxmEPz64wpTX
2CI+nANAJDI9GkMVcfa++xh8N1j0maOUgPP/R74CrZFNnGgiulC6WVTKhDCJxIsg/6aatfvqKqlW
17B2+CgXOYO4kREYupL3Tm4rd8S3nrsLaUR3V8zQTAgmInjUrgcsbI5WrqiHPTtk95FF4WJ+9J0O
qfC+gfcWudVrNUH+jNunmwEPBNOboouXMUAA/hZn4VaqDq7MWGncz4PSbixpiMMSdpmnb64Dy3pH
9y8//VqbxwFq0fj6BTjYlH3h3i4rkzeYg2rsLch89EJm9ewerE8qxhFEEBcbindymQWxTXQmoFLr
dpjV9HYMC4hbDmVnuL2dXxDzI+xz+AjNmHOk2GJfkv/vEh3fGqaFgAjGCHTXmTxk3e8pY20Lmzwf
gqwbwG5yd5nDYixnnzkgJ/wNDbzWC2Y2rD7FVteCmJ33iHC3fh3DknG7GYB9ICI0iPuhi/nG0el5
nWZWRnzFuY9Hq7HGUEgjGcNeWOlItqjQdTdBkTFq+vo2WOhlSNTnCy3HjDI/c8oH+3M7WADAyhiD
7fQ9u+YTYcc60wsi3QCSyZt4ggF8XL60WOKMvMNQR2oDchtvfi/28hhuBi2JMmKry7I9OfNCdbQZ
cN9+DY72yetp+Nj3CCCiQrqpvEBZZp0j/vPxoO/k3JTagvntCIx6xZUCbewJUmoIycphP+BQhFWO
igAziGTZqCyheLjik1lWIOpP6oCOr09JdcQ7VDFh2bvSH8jXjLLVNx1lqwsdOiHj8DcgcmecuP0J
8NqbmM5E/syDfGYZ3reyz5kH+nxRzorv8AUtWe/7lLbGEoeL3JDiA4YR34uFn19YviIYaBK6RPhm
M1jwBNziNReMCxQMosiyDNWDpekgcGecLCjeivsyhaLxMtvYOeZpaxRo5dI05DCAWmddiCLHnPdE
ZXpEVpRzjwva5RNuUCUAak+5K6+BpAQfMj8lAoLqzgkJHR4uh1CV5ymIkxk8zt4y8bgDWuaYVnC9
9p2bw4bJ/dc6PovvtoQdlSQEC2SA+Acu/lQqMwUdc4eT3Mz1fOGbqWbxPsAnI1oHQMcqgUIXkV8E
FLC6rKEIvUs6wODBO3nGcKcYoAlVwg6P4O3UC2vQQXr4CvE++bLozL+0Ph7B/5mGpEe4XNRLslj8
ElKZdiJTRcTxWhXcbY/rGb9kELZeEoHnGjGEt7nuL6q7wDWpkDoKzAjhkh2XqJNyS9yIamUlkx3e
vs0lcCyxXOEJCMkB7bk83uRu5UIR/M0OgRv0j5VWBPLKJbtf6jS4dAaWFz/X+KGscKKD/6y3AomF
Xdefx/DNWXnKW/4OnSQ2L4iGAtnLNAUjXLHa9sOBcIws4LxDIbboqi4z89yhi69d7llvwiz2ZMFr
F5w7sKDf1UMyABUQgYKsJLpldh/CWpxEr3XMmlD8c3g4AvCLyyToySvqThJjVaTMeNA2ITWs60LV
TiZIWzrk4LoeYBBB7+8Hg6d46HT5NDJ2UxUpkDys3TFFJnf5T8QWnDeoUcYcpNhysXQg9g90eexI
E03xPKtjxEo1RTHAClFrCOH3WQuM3+0B9Bs78bb32rpBGA6GondrGAuemUixubFunXGlBCtmArY5
p8HzDb39+6DTnqc6AHpn/IkBCs7L2nvvbbihFFCY4tazVqXGGXD1Kq/oxQuiyzObOQ8H97jpNKVr
gQAYWiC2yAXDee2usumgVgMvYyeDHa1UJjV/L6H53U1azatli69fanGdIjrVHkleby3vftTtD/pB
rd1S0vJAUQAAcjzIgaX6/QISQEDYqhU7X+ZJ85BYqJHeXKzuS44wqapjHJcjzdmt8HGh1Lhz1NG1
D5ewBPQxcHhzgNhRG/7Cb2l7ghBU0EomwtSgdW+uDn1Px1PDOfUQRy40HkGsXqbaU6w9seQ4vmBQ
y2xuAjAYfZ7WMMQNnteBePTjKDkQlL8WF9HKTN2PbTNhRq4z4shdYDmrpQiSLv6f730Vqkb3rBrA
Q1JWZ3t1XE+G6bpFShtwM8In3xCj/dugbLZBBk4U4ykmrGQs/2oao7JUWA3rBhMiswgby85uoodF
4ahFEtLiumWcqGp7Bfq3YWN9ySvtlcJ2xJTKU4BK9sfRAiBatvKIb0/jS9MTSRYLttJ6mT4ZckkQ
9FnNuG3E3uzXNMAPOAAiZnWVJ3vOo833d1e+Qn4j8USurCQMhz/GNq5+TmfBQaEQTFZDT+JlUafi
tqUJezzdDR6QD7ftCtSb7GYARmKr0uaGVWYvg9JDE7f6lJb04Oed/OS4Y4lXepVyOz3u+lk0t6bm
Tjbx0GirvA5B1CIH38a05sFrIULfNuf9w005qpwZFfrovinDPooX5a9EipE6tzPaCnej8zW5/5Cw
d6NpRhGC3IKk0AOHF1zZt4C2DVb2lR7KAWdQDaU9mifdHPTnAbFuoSoKo/JPQ3vrpJeg95YWgQ+W
VgzU/UBAd9txhwdE7GfUrPAodYNG8WZzi1KF7Q+fmfAoYnCE7MvkepAmx/l3AQlhfnjr9G5me63r
g9BCRiqwnE2PwP8rbg4jyd8hYyOjJ5KWVXzemWHyadiot9I8rdd4MkbWrDBXGhYMo5UOeZzYdm6A
WgjmXEM+pv6EI6ZWxWdhW8oP/TVcZIhgVWnlwg5C7RCQ3rDwW4MMvfXEnvMUgKq/+d7o1hHEXC8d
VvcTuqaXFuFvXPHTepYEV7o5RVWews7IJgOnUCnsrdLrwj8wzsFycNKsu98VgKbyKYhZDMK2a6S9
wYNx5QaEb44DWVDJiruvrkSxR2LAe5lJzZyzn1ET9KfsbpkZwrRfEWTv3zuQ5aeWyCE47BZC1N7x
sEq+UYQocGcs4GtwkuHYe8Opt2wtjMeU/2cqscnXGWuZiFF4+k65tOwN5CdGw768HBb/nzYQfKbH
pl2F9rPoIGA/dLN5BRsFuo3JCjaqAKGTchoFJu77N+aGDbZYuzwrv5KYkigBbBXS0grUwPCwjKIN
ePpYEng+QemnDAKj+Osferw+msRvDqg6Bejxq3ZiLh0ajv9/B6kj7ro5vXmyiIzopYWNtVruwc/r
C9OHswpOKp0pXTPaxwRnZItUhGrupzjngjqXo+0h/Se0NA9nKM7YYUvv20cuGa6xg/1OoIEpreaR
O3tWd0ykKeXp7g1M4UHECxHaW/Cfg+k93qludz4gQ1UMKSSn4Ch+UyKodyD0vsUHN3vzhT3/iN9w
HGCQ3lda+CeDbM81jiLioQ/Sq75wsRW+F+q3fSjaa4dbVPPe2F3rQPjvTgM86uEf4f6ZpULt42Fe
u3/LE23lGQUfr5EUh6oCRg6Y2xvW6hH8stIHTMKJnoL3O60HSp1YvL/JX/Th6Gi5vXaMUsPNqkhv
4Vqlmvwryisc/kNsJLZvIYm/tjnJoi/5X4feBgtCjS4+xiWI4ydLWm5Uf+UoEaaCRzQRhPrb6iwC
fYe62+4EFMB2q4A6FRzs9nifzYrtaR2cTXbYaTxd9LTNuWp9yT6vxmht4ZrSSybdkEGRh32Q8Y/f
LuquhmJvKK+u0BvIPnxz6yDkoRgCKhCkN215sDI4V7ukfuyQNG6cNvRE6mawL8oVie8gpqhEQ9z8
G3/m43UuLDzzDhmfDSfVX9ESRy82KzM3g94e/rCQzUadGtionWWWQCA6HTMeJ+DsrnIC8GhI3epY
4tWWSR3FS5Z1EOBquwSfsDzcIay4aHqjkdax7WPIkkvtD+wBYx2JB94olsyEyOoyRDJklDgCHmPm
7GrJrMkL42e6SoOk3ar8F6mNHqWIyOtIH4Pio1GdDZy6qQ8hX+Zx4KnY4FIE8r7B9uP2caBx+KyR
Yh6K85Esfk5R4WkTwUAUKU7sPKPaBvFFmNxjL9MQNWGMxVINtB4Xtbu18RbaZ35vZaijB4D9rlTF
gD6nKmT3CgyHhVOKxstidjmwjznIIh6OFckR03ugHvPKNNX4E1pkBgl0ZdHIo0iXnp3q395SmvcR
0XHr8wdmPDHyMIoMf5p82luysadsk5EWTP4rJvXwj2epEACLUM4uq1KgjRMEDVkpdAF5Xj7UUV1r
IiEhAgnBFQBBo8+bDAWrB4/w6Lp5oG3qV20D2TEsxIHSkoPq1CZ1am1ndv4JvFiZbxPCHqBkETtF
mToBUo1fYJrabQmZsQn7+vK1PUSLvdoMYodQR3JgFbFOa0EG68h/l2pbhlesQwF1fTwMSLIZvKbP
LiRPwY4Y/s/fapTru/ItXANMjvifHuHCd3b0k1xKvqhqlFCdn5WweRElaOlQlAeBloSLIefQOYsa
B26kU2fSlBYgb5HPy3KYPiIuzeIW2IwgIbRnHdIzT+dlBQF97FDYZuyPVF8I5GT6PpJ1KbEdige9
RuueieivhPTCR9KVHVfJm50k0M+7RDFVpcdI4aFoPuv5B1Ovd3HJbxEbxClPk0loBU+Mw207Rl/H
EYicmt4p1vVP1Ftok1cb1VGH4FiePSAag9MunA77Kv7ph/bYL2Moa8/RPnvpTguSIdcbBQz5JSoH
kNIcsdCmbMat9zxTMsPozeRvBhcH8gmgmstSQsuqXaWVCjyXQP2tnfqwK6WNdIxiA7SHc22b7in4
u8CNlr1osetX1xF8G9+tUqZO5rxv5L2M41iglpovZqnuHs2jgjk0afVOM6ycJTJcD6F93AMglLb6
pkdgCJjnILek7cSliJrRuoq3Khet6TlDYG9yq5whR/O2RFdrbC2l5vqlNHQKvfpOEes7RbSjDW5F
w5NZEGVnXP7ojfwXbvyPJ8NyQUf3SCkc4WF5hOXD9L/E79nRdVdWLXBi6R6xCP1PIwj4K9TcW41o
bvntdWzU6y3Shx5QPARiEj8vnC+LdA0JPEdiYmWh/kwWoPltI4V6nzXX0wseQiOQ7Cfjm1fYBSUb
aiYhDcDFAHsrPpqNDms7D3CpJdyLtCcOY7BXv3E0Y4kYDuUvsJb3ZdqcUeCqq1JQJ8NsXw9HIKO5
8SrmJSygp/pvNaVS6eA11am3E76UOo9rVdtBdhGLJlUbRSYlEtw2pp79g9lHfoa+aG7zZfsWyJZY
q13+zOvhx80RT8qNfTyfWXCj194R4Q45MfuEID2pDGCTJW58KtbtwDK5yoOZvvTV8f7B30gpc8FH
54oGhpOn3IcqtXidTbPD3TsS8j7dEBDoVZW3j1QDBTJDLQ98AYtqFrpTgKEuANuLF89c29+RN9GL
UfgkA5/y7e+T9AnrWRRJ5MIU0HAViBnYLltLTS1PCXfFS9Tbx0oRzn1k3feiRV/HX5fEugXUbesu
NzMzaKB9Ft6bZA4v18AIhfAUUbts1/n9PsvEGQ5294CcKtGbUz9osts8Bb55Hz/ou7JNq7YzQfgf
43Ml4YG1IRT2l6oKthzFl8USyjNEYop9CJPsW8mIPdkr/T4qbGbnPmw2D4plzvr//oh3lEFUR/uN
/fXhi9oeeHYXkM19XecRMfg1s6Z84/L1nB1nD6q48/Mv7PfxA3N9ZK68EP22Ya3nmkQBSQYFa5RY
qq449LD2uWRNxmmNyYWWgZqMJ74tJ3zsdUMllpMq3aEhlpEQtlyF5RSEBJGF8Tt2bq9gwNzp+2hd
H6+Lr6c78hkvrcfIWIJ86W+gKKPnu0Z5vUT+GJURTW8TuKK/Wh8ihLHtjTKeaBqSlrA/5BMExkvF
z2DmkHqua4KBnsfYaUdgirRtvQuZVqVtTR80ouk+BR5XwsGbIl1CU8i1tMeTz/KGwx+R7lqzDPmm
NLGfNBeu0jxQ0fQ4OruFj7PvGRqGeyTi03qtZXNNCixjqyiRXdONEk3MdcS0Ogt4rgHOhMjcm6st
qHAicOoHqfjZ7QaeUiFUb6joogroc4p84DHlNYiZ8oc+DxY1T1pSpQO3pt27qDRI/OfRnlXT3lk0
ghcx4hSYLDvQgcpapE7UQVRgLFTkfnC0awGscdfpYOkegBnYs6h5na+6GJ6sG/FJKTHPPu705w/9
kroaANVdOfZt5FxmpyzBm+WcgiEqDOiekfVHPshqxyQJesxYHw0W9WsUFZzVkQ9MIeYHCIB1srlV
li7rdTuMF4RfqMogJRj9hRbNY5k1dyFgwRrW1I72wV6ga/XUIF4m9pqIfonQGMf+9w2R0/qeF0f5
y+F/802FvZbnSpvzR7IY80EJPmNJW01UZJzxKzLj3SlV93SqebjqgYyQov3q9gtXagZuHYiSc3OX
Xjv6/E+Gflr/tas8HhzGnfkmLMOer43NVd516t2AX3bYiAjBb5lPrx6CbgnVVfFo2eue7JQSTSWm
24AOlOUy8hQfV6TXdT78nKlvvQawAewqHAkGxgclzBMb86Ar9vCBNCVSkaf37+BjCPOGINXmVZE9
UoVi5euqEfUF26RjfLIjVKMdobJei+Uj5BEzdoB6/5MK43Y8Peyz4huMAKdqoIAuCFA3ZdRMDSdu
TFcRxP92D3B9stOQFL2brcctz3yR1LqXlfngAADxionDWHz14rfHR7Iikq702dsgS1a2y1/bKxOl
fHWCwUpW21zFhve863RF4uh0u6gpy4ueSRmgnezqWlcRlUD+sChCL2Ot/MGkdRnD1c8xYcpZ4g6w
TbZj51NUX2jvRC2VVOxuo8le30prEEVV++Y9DqvuXDqktHuiUWp9STJzzwkXPKTKhpflAu7c24Tp
s2WykTsrI2Os3FqAMiAtNfmSFGBPwRUcoBOIprp4YWAC5z0llIY5M7EZGbBGV+mwnBTMfzXmF9X8
CcadZeNMsWpeDGTS1KzbI28P5qjWt45hj4nppW5A6A2RR2K50SB0zgD7WO2jduu4VMVZoSiW4yGD
DOdapNsGFarPa77z/Nan1eq+kw/g2eLnxJFTW8KIk3vRt8DYq1NrUu9s7pI3hovoRN8DQWR91a0h
Uh8zbDoaluKvxUBX5g57H2a39HIAo/u/amMhwk8mh3htZ3kdZgDQ5bEbCokjl7fktya+QSzpWBa3
mdIfTSukeMfgVHlqx2PvDzSsya8y48B2fkBndl5MbO+DsUUphp5uIs9yaQnB/F0l8b1kMUsmIe0U
/4S0S+/K5vm5wMGc+Hsqz2WyFTK55QpFX/Cv95oIRbm27J7MmbaPoK18TG1GISWlSjNR5QiZUHGz
y7JJ4sOEVKmxE1SNoXlEFq78JjgME/q6vzZPfKGCXekKkTH4QKphGyvQsL4ll6oB9yPp4hyoJOTg
+Q5DoLPGw6TEPgpugIj6qBhw4wipo0i7IIRgkAov4aQaIxagoTCHqW9VYEupOtEEHNYk9FzheNBs
5aWG6ueJfTbd0Lo84Bwdkv88DEMgc0BRjcrXRpieqmKe5N12KEl5MjubWn1MMZz4lU92zs2/Kogj
Si7JH/234Gcg0A74vfxnpR6JFxkx+H2hXOuDFO2pF+nOPpPUD6evS6cjDB/BwXE3xzqwRPR6+6tf
huBKkJQppTCJhhPZ0aBcciJ6svo9Ma9Ty4KdFopGmufD8xcEXWTUHQx/N9Abvm3ieTDyBtZ3wiEE
3JrA19OgBvOYtoFNO5rw1WGuQhA4WgXsCsYiN19DG2UESy1FE2Uwj73CpCpkGV/Xx8IsU6IfRHXy
loAiytc4x6zx+h+MGfLjcrdkB2xDbbx5wy+i1aOJSXOw6CKFS5DVFy3EpYXHiXsuBiolmt4k/YQB
mJnWtehbKCGwF1Vo0Djas3fdyfFAddKdvnmFX76wdqESYZ8ud6s878gl9oStPu7kBpE9cDCbw0lI
bMGgQwfvRdtovoacJlrfN3+HSiRqC4NU8K7CKFJKqMifEQiYzDzpEELt5QwlKNfAvNrf1V3BFuo5
7CZxSztOQNbbIpSNQAA8DnYOcEGRiF69zIGj1InLEutLXeCoLcUnqObFaJzXQnUYwux5cI5FQEB9
HHR+A7IsZXql/Gm56OtmkLH+qsUXmSd8Cvg/XLIDnarrHO/uzZU3BhBNONB0Gi0SIiOEcgjvfT05
QsrqvVXDvk7PFo5B1jvkHLMxfIxD+29La3/qaFgurhC1/7FkUy/jKohAhKrmuiSDvB7Tkkrn/9yS
7h9DhthqmKUwZPPiI3QXWzofaHMU1x4J4iGPXkGBLSWEOin4XB/jBJut2R0ppoHKQb0yIEZElHup
RqJIxxSmsKyXkmOE1TD0Xhl5j9FLG5M0ZjnTFuUKYVPwa68l31ZAAhfZinc6rsDNQrHJCg8py7f1
kT2OnRutqvzsugPWnO4xsRu+vHl37KTamARP5Q+UOoXf+Iao5BDWAM9N+CM/IYmSxkE8z5Zf5itJ
Yu6CpDb1KY/nFPuBG2EmkI1i/Cuc5K/gzMjK6N55O3pZNRLYsqidCc7BOoS6zoBi7RGoPqebnAJ0
tnGlC1ApIMdwJst4MPg2tve5XYcGP/qE46OepdURBBmNIcEH/ZsF6Pp1lmr2fWwnu5+rYBkybGml
26WriXZ26kLr6IDnnCFTdsXL2K6WfSLIjdVevGupKdh2BBdZlcMm9yQyiG2+KgbUqQRJHG7nTQtH
CCPhCy19FemCUClOrWb9rjn98/HHXtq4uEwAZxM/1UplmSnbAicEPOOzFxgtzQZ/Th29uapWfh2O
dFIgxMq1yOEx/hm1GaItv6vlFLgnAjpI7X0HfVz11kaQfm7ZDhVu3M7g6WDRX/9Q8Y5PpF0Nn48G
mcrp3/wqDYca/W1Mtm2GNYcaBfmnGW1hGeZ+SIzBHI8Mgt6EY6iMbI4SEbQnDtUl5YyzSavjEZqQ
H4/Dprqjh+Fs3ZUfGhfop/+9GsGo8noo5G02cJog87P6WdZo89ZJUBz6XRx5KejNy6a9TVv5C6xU
xOYf3D7SpBSaK8EtNy8ZVt9NGLUhrZqkbS80BPNwvqrpUaZnL8sisW5drps22mlkInQ84RWTWrJ2
/rkwDlO6bbIsNf5SM2KwEt6wS4EUNQoyVx7AtJXDq9Ybyu1vxnSgg/QNTDpbe1j2bRPp5NbCV3ED
mtqqmaNQSuMJv1UYNdfPmNcJ99brNnmhuyIlRgvlHhEFi89dZvA3P76/YU2mzTz+/wFAsrAAoUSN
BIQGiePdoNGz66EpFvLCfaHJUifTDH8IGLa3GR22AIm8DElDBVflf+cy7eP2NumkmGxRxJsAWhYn
YAQ0exjO8O/GAYJ59FReByPtOXWu9yjma9XFXErdXbX3M+g8DtmTcraYH6oM6jVMN1bcUCOqMBLU
HRYvkhmOUhkFKwwvbj5G7yqYIG2gGZ9UkDlUoh2JqoiGpaYm5TOWJtxAIOADH8mDO2fHeTjpNNtI
oSKC8WLBzRS4QpKBojV3vSquoViLAvAs7pBGTMQaJXibhE5IPZYLd3ufhSp6NU4KpzYKnk7PiRIn
1s+Cf/nJGE/cos+E0taU84jnooZ58BftxfDmCIqEJd4pvAaIJq29bh7XWr9DDpF54Gml7U8JxXqU
0nP1W0if5PGyfB+AzbuG4ewmHkymAjavYnHTp3TwYVcmID3rfbySIFhHJZ0DWahNhn5kTn1SchNg
GrkEaY+Y1iJZhchJhZbuE3gs7V61GNZNGbaI4tDKBix5mNm+iU+rTFXNDRSuJzvVofxMmy+EYuLg
TeLWzzBDL2QqQhoJT33JASzI7catO/PWlvAPmopvmHeUPled6yLihC+d/pnXzOlMspGIyx/+eqKp
ZmPZwaY3v/JSxhWbwAAm952QQbDjk7JtlEzfHIuYHPVTTD+STlpbTI0PGwpdNTnnqGt8QFdPt/JR
7hKPawo/KYZnrM38FdiJXnWHQt4syCb2+Tq8uSHU5W4Iyf2G6J2bbDEahk8xhHpOLsudZl3TGtiz
DRm3bkvBQhoNO6Cd12cQVIPGwwZ17GDdmb0gTxdaeFb7lTBK3rpLozHz7oYs1DhiQ5g0fSQ9fhIe
YJI2Xmq6hvxGCoUGSIkaMEJqK7V3m85hlSK6KQZo/GFPmMRdvyZ3xWJEd9BR3Kn2xzYkvvUB/rQo
pH5C8JcSIEULcmpsHgElCvJxYlNoFERdWmYjlCJjkDoxjNEliMS6txq7A9tU+X7qfiGUWsIPxaDf
x7wlNYKywZV8MHbQ2LUJobeKzqtyRDk3sDVJucyJVWAn/t9vR6AtrbSJ02gtHaP1mACvbKBt/Ktn
ZunfyFWqyuf0vZ0Wv5YOFOMxVWgUYHUdqrbvBsaEHNeZ1FLiZkjKCydITlmiJv7fhhXWw+SYIO3o
fFfhL/9NbF67A4kf0YMaEr4y2s1jn1sEb8TjNkn1Yuc8aqz8zwyGMZt6srD/IwNOGvVKdn67DrpJ
AJ3XWEg7JijhdXUh/H6IL4lPGU1OXwgA8t//bKUGCtEuzbsQQd/kyQX1cfMTISEhlkYlX/bulhES
BOxiqJIOBDpbOHr2f9tESF2dRPbVnjuKPDs2pWU8Do6RoBPKw83aMVw2Me4AckK/YkyQFaFS8pGn
BTkf0o+ykNRQZiSJJ46WQI7hfzIHEeUeta7c+HStI4PZzq1QjBM5AGN/fA64FjlUP8mOwxtxWKHm
32cUqtTBYZ8ghjc6Z8PI23ISLJT0i5JUP2y/rXFl7T/WGFipX8uEKV3+5b3vVeM0ZfK3O4qEtWHk
un1wTFB2pqtnk6BpGrP9m5znL1/bIgGAHn2vcHYMeOjCi6Ih2FJVCv4DF+MuF2wKc5wMMx2dNrrF
Fh46qVTT76OIMTeB9w3oMIyTPAJ9Av8GXu42zBgolq7IKfJNiVtaN/VlIL5FNAUlczXLCNOg4v2M
+Th/VBXtM6IsCrfVvETPbmisMTFcvMU70Eub/E6qgvfDDb2Y1oalFCpPUhyWEfi56qORugThWo83
YYamvi1DReJAi+b6Iv5iIIn6Xrsv0N8Fwz1QYLhb7zvSG8fN3cEQM2cU2K7s19abRLh3hE7s90CT
VTzGftVJHcOSGeDBACI0B0/fVJfiLJ3iBCgPGN70NOCCj7TnxGom8sy3xLgsAn2kN3s7lrJjKuZo
54mEujQLoX94texkQkbEbidDu77Ggym4nTG1ko4qQwRvWMcelowS+JFKGvaLkNYc+eDMlT4d055G
dF2Cjyqx/SpIJ6HDYR5m05vccri01bDvOKjxGS1u2QMYptIM/YNTASo6IufWZxblGsMA6wD80pGk
GqEbQasnYf05rE67liK83ykzFrhBm50uIC3VaYU48UHpCTLywKq7X2bDNvwa5ETvbYssFslXiR6w
RdE4x9vLAmkyojdA7tMnGnPPJ5lEfadde7AJC6wSwHOb3BI5jwnrphELVjEQSN4BKBgA65Sp/ka3
FG9cpWLxspbK8fiEtjZgknhB2kFJDEqBR2BTD7hfgCLMSuEjVd7O0g9BmjpTxgoNhfxrA/IGj9wQ
dYyTL6xqSJkI0ruNZae5NRqQw/WYJ95W+GcBOthZ8PBumLZsQCCJ3MDYs6qljolHeTynitpBYuQ6
9SOcbr+E+sT1obTkSt8ZRVSLeDY+XNIhGqb2HHbaRNVnhtj+o3gFSlnW48GKqdoEOL8UUk4o7Q1f
3wVvCLyS7TgyykSW+aXcl6DrEGDaCHnABfne1jbb+qqoXFeLy2xni4PMeZj0vpJHjAYFYwiGfzRN
T1nBZExWwczcEOmYWAEbbHYxbxt6THiuHpEmRDQSclGidxH6Qx3IfV7MdgqYsgpnF2O4HJRFLIXh
YPSB2Yli22qwjST0YeiVqDKc2xzik4G5wsE+Dr+i+99OdOc7+ftG4cp5od+ziNCog+3DXncA50Hm
0PDhJrKKtnsRE2tVxgFOJO6UeK1xvgXVp1ISVnLwYWEM9RFy3DsDJOm9OJVzEEe/0fFvL7CjPl+l
UodTFYTkQVWoxU/CkgQJ5Oj30rDHl0TPC12tSb5e7QRYEGVR0aS1W8FN1TFkjIC6QTI9rv4KixfY
aRoShw5zv/Y/QB4xB0WXTZUYgrKN34/Ih1o9NFLB4KB0hP7SHSZr5UEHlLg7WHACu2UaY5iFI00u
VR1USrW8KVTTWpSjOyFH+0hHYoj5AbVLIrxTLpQCKXjONybXyCBmy75ymTSYmSAOL+xoTlTDmJl5
xdKEqEj1sv7VGcwKXYY6to45X29EqmjHcp8Z+U0GOu3eRoV2yYm97uDlsYdJ2c4cC4hR6KEGNdeD
gcCmBX/5RQKiMVbTopLi3TOV7Izfhyg9mqc2a0m3nrbVVuZI6r+CZSG+/uHo1leVBtgcr8TihEbR
NOC5DmQAkfaMTjy0TNXVySBoyJ5r1cgzCPt63ICPtszWYwjU9ZRHoWEEK5pNSvOBs93DJmN0vqxU
CYJ8KjpwLLAGzcbtJxDCi5fxNJvvV1dBPe0XkYWsBw8IAl9xOJbIXkm8eExvepm2pPgVF3ZrIPxk
laymZJ6cNY8KtDu91qIdGwdOdJIs7ZdlOs0URGOC99FAyclaAdX2/dWP2UYHflaOrbBubp3u2cgT
o3MD3RoqADIWQF284s4f7s5TiQWu4FX/Qgpvc7ZIRhmpQ7LWhkdiSqGzfUDIAfuho4SENFonmUzp
btEY2DOVz5VdJK8yw8JmSEZJd+7WXVstb8WlnB8hx9esPJPBqTm/Zfu1+Vuc3qWQmgj5re/o10Pq
hFfvOlR1gvne1gZ8bsI1PyhhkzgbCb3SQREpz1T9kp0MILluYfPXTf/aK6BHk3bOWQrHKjhJ5yzA
aR7u+AK5XFy5P8LxP9OAU6Hy28Fx8Kuu7dKOdL021toQveCkunpAB8xfEPu87DvJTUslStA237jY
jTLQIe9/tKwT4T5dWV4oM/9U1yV73sk+ObBcZsisPmUtfw/PABvP+alxThvw8ZM88YBRmoKuYgQY
YWTZratrVfOi/8BRtTLddHA+CQxadz51MKNrjLjkgNGXhTabEQRzOLugQrTQlETh2k5eGFLV0Xmj
NXTuziKTq+oD+lIPeJRNSYX8ztoHaCvhiO9twTdnwq6gCgbgzv/xhytDg3rX/ZoWMrZu3N0T5yUR
tCiXbkaO03jNcOKM4fGqntxtrx2fs5m9ZqAW3gagN2qajnNMBzokZykCpAP+f5uxzOLajDs6t0LG
cKQ2RcffoaGXzEGJZlpCPid2jvei83m+uoVymx5smwdajqTnEzD2BP+8hzRU3C/FTOwQcgHEBcHa
HdLFRC0r8UTf23hPKNDPSywyHb6YLZCWjkVSJ5Ke5utftqw76FmMfP4L0U6OoEPqmmFfSyMm+TBx
N3z1gT0xdSNRAB5BVaxepytzotWlpuSIW71XPgoYFwsRoWeBPpKN1wLZkccg0E8a3Ib0zSB2S8sd
gOqOr5SHwfskShvLYtd0vUEEJUK+QiKQfE89G6UY0mBUKL9ivdMEs35U6uMG/YxUqBl4uAvdhzsv
VPLLs1GCM4dckRrDPrTeBloQ1Q4MhLHjyZI7DIg6U2yuTEcXtfIDkTXUCF9860GhdHg7IeEkRGXT
vRbsUxUUXBR1eyroQMuVw0sZGONYmUG6TfgM7CuDmO2N2yx403JRZcX9xo+2ALqjNuvB4T6aI+Xy
Rw11a0A8KBHuUwWfFKbQGja5TwIETYgIDqT/OhjuvwpAzmbkFz/fcCv99DRS3vLcJsWi0mPYUcfJ
/8l5eh6kk/KjeRVnVL+P5cLVOkYIEmc5SmTQqaYBxKDkneeYjfzzly6vnmhn3zSHtlLHFHmquwkB
d6rpiDsoNs7Gfom1ZDKsgpjDIi00gkRC6/JHW+gFAKHduSIDkV0MbXojZ1wem547/tLEmY03WJTj
+NcoVW1qp3fEkEEgvJucXeyqEQjoQysur+kGr9vZzeZ7QuJCIX1poEDngpQkBbR1FVyhSfm6XzX0
0zb/CyCxstZLHj4PI7YIIq+A1BEhB+gLf4pgCF5i8Xr/sgnFiV7JrSfhakDUx7NGucb7Nj5xtsF3
F0MKBxQjZ0JI23Ym0aG6PU80hMtQYz8NjmDz5Gk494WRX7lV5+bXowaLAm0zWXu+zyKAPNbS9qew
JvynNFEmRArKkvVdhL5sK1aJsGeneTx61TVvQmWPrDPAO3kq8SE93JpM2E4mSJ1G8a2Egv3fP/o4
pBhpYV47L2BzGDilVNBEzsiCoOjOzTbbHXUXO94BkVkCmUgj+4UI/VSVTxm1e16WLBE9SAfmkvEr
W1V6nFR/o1oG4vrfw0z621jkW4ljZpy2xzQRkvEKrtHS+jvqBDIcA8bpS6zj5rlB5J/JRGhRvzJk
KD8kalnLfYpdO2nxmqDEX4gCS1hpuMpNGshVajUW75FmW9L6Va2wI3Q3CSFYVZcOqzu8gu3GwYyI
msyOJN8ZJBMlxm8ba41BK3EvSDCa8wddvylXMtXUFSg+vOn1CawuTky1l48b59YdzN161pGboMo1
180V/ikC1evs5alsE6KsNUxZNdde1Y3nM/Odv/vWfa57fNZaPfLyh2BjMLYVT+JCUbm/WyU5dMPw
GW3rp54pxdkC1Lj5CWr9knXFYkdFjjzh3ryzIUGz8JcPvmbME2krel/82qsvV6AIMz2078VManOI
ODTa+Z4hS25HQTk3EFCRAI/Lu38F+YUgTKzYJsFkANeepP+ZLif3E1gEVbNrpPEuA2OwCSVv1NAw
vAahy1fK8qOvfhadPzSQKAxEqifF/yrIDB2NlIYpJ+8GAOFyK8kigoBB2L4Na3NsxGvJwr39u8Yg
X/w01r8ZuGilG4QxQL4djduijjYfM0enK6PWAtvGLtCYwcNZxABQCGXQ8wYgaREwZQFEA6qKR23Y
W54Qt9c2l70rhCMnSKKSWLYX0NZ39pGkbUEhx1sV8cUq0GcET1c6u/vnkkXeKuP/y40+ZExduCD9
JHiOiNz9+2eTFrHPB/1wESSQ8YJYyIpNFhkN+pHD/lZFtjFrYXj/azc7kldhGRvzU/V/PbyqPGTM
eNxsKLmVWVsrW7SceVLA4gRKy94d+dMiipBqEynhKHDNmkxy9E9KHJNmrvyLXAusfCdknrQQZbMk
lB7Moy5WBRnnMjmISgTLRAsIsdUw6n04BUSvKqB3lQF6VNpVcHXo9vWE/UNvK72q0a12Rfl4chiR
vyVT/cc6IaZVRuQwJYghDe278ERDLSddz4RKklX1LDbV7yGXiJc1DWtlVO55nIBXXyi7sOjjb2Bo
CPtJ5p8OPg6b4AR7Rtwd1Ca7FIS29r/xyhKK57H88XrwbIddMLfusJ4hwsO8PdyKkpAnD0kEyoCo
aJhvGumfGceSieO+HkONviVlPnfDxQo8P+ZhmTxph2mZSwr6fL3sZFRuscf9Jodq4fDDCt0J2Xy0
hWl30UzCYQLUTh7rpMDJDWxUxL93s8WD3vt9gcd6KnpjjScRtw5IXK5PPftrnlRuBbwt234UJ74p
+gRleBOXd9PvflxkOKbOzAZhW1oigg0I6kboIcPMhizX2y0r9HccTAOmUVrJV3LLajNz5iD7TsL0
pfhD55g73nRbwVJ6IB823Imrj5nheAi/x0xrv0SMpWQLhIk9aubC2e0CB3g7G9DGrv8je0ltysYo
lA2d91QKap2/oclQWm4kiPQscPNMW2o/YossXEG8irU7WVGXfdHtonJw9FWPDuAml3WcL0ybzJDF
j54Z+WnBCSVli0MNbStT4aZKs99Pgt64Ur+aOdpcU1YsdwlsXWAHEdkIK6CH0Pssj8sIIovT4UHu
H3ImZPkN85SQLWMdq2ODDZral5dSDfDgyY9C3getSMUYKwXQHPyXRdWPFZB9zqhsop5voShDsDR+
KKQwfMT/UimulqXcaFKvGYyjcPXcZaulJsrUOwm92sTaXZuH7obkrcrHk5QlXYz9OTv2yrTp3eGw
MAlM4W3ETPr6fXUhMgmQxECs1xDkhlilM7nlva3he6G5AG3E0a1KlOmWE4AcoObaGj/ot2+pBTqN
2GVSjqGhkkk6AiG6tY6PNgLA4PTvuQGn/fQx3q0efoQTP3hhl3zcWL9b0NNUUs2id8vNQenG54rO
gqcSZm2UItxF1YNEppu+6yT/hViITHrQ4efAC3IzWMBtGa1XTeD3wXR8FpH8gykr0fjP0zq7dFHt
mQvjsLEB2KUsc85/k5yMi+ihe2CO9Yp0/dQqKQBaxPnyLuBQeoBvHSXG7NRBuHdho+tfb8IxDjKW
tNNKQ5ELt6OP2pooSYa3FsuNPP+dugv8u/QRNL03rdRjV5m4SL/LBaobhfZrOvIfYM2Om9CBcXAX
b/OESSWaPoxYRuWFd/k5/ysTj7YEWV333MkWY/PXBvUCDCHNsq2s9tZF2XnBrJ3md0RwAQez2ZM2
5m0OvgVPK4ajMv69pzwB4lYfXuVzLFyOTxC53sh7HcevIRfIVEvU6OOpSdZNLdhernNFV1ce/Ogv
0xwxgR2ztdfNNYE43FGYJQF2o6GTJPzG7j5WXxP8S9H6coKo0+oBJcTMdYA6vIfveJGQCcyAXZBm
APJqmirqgz3dsCgze/6OGANY7lkr4l5645gwVzziTkHq4FE7vma0BCsx3D8NbNe7k4ff1bQ9v46e
tfUl/42TiWolWB18IsFBIJ5e1XB13hqXHmIh+HqGr0IHifhwJJAkq2x4Y9I8NwNCiDpGWPZfK4gW
JZobz265NLMxBPqICyCGlmTJi8OgdaCoakVbOP68ZXIF7gSXE+CZw7dlgKAycWaTzOCadl2iFHA2
IE6FikOtcrDOAuChfAiCJwBM5Hgp/jNEszpiQa6WWJ0T8Ve2M8pwUokkoHU7HYUqcmwXxdqZ5j69
iK247WnS7YLjkoTpblM8BIG4LxlWl5URRPCDBppDjkATqoxtqLsxtQ2YCmusGVCC4bBjYCq2IwRP
W0gqQEeSTvo1eTwwbDTkUX59DQ9jDu8zfyqojwjgX3tXo1xWxcNUCtOgZNX8liP3jmPkbMzSqTu/
m/Q7aYCs38RjDMV3tSroZe3OeO8F84K8CPH57UcVd80qhuKUiwuBHW/NVFnX2RiMaLWQpNgbnx0Y
409qwEJwJ9xFqvkfSNGxLiGkYwQHTJiPeRyCEdYOSRW9dcw1Vyet27YTfLKWHcphjMtt+vNoX1Sb
mEjvd2GQenivUPV0dyDU2PtKx0Mt0FGT0uyNYaldEdhuxbWWbLLpyjpSJDB5do7OUaFCKYE2Cu9h
qISel2c6CWDiyXLO/ENLokdNwonYU0FeMgnWyc893W8h4iNqlqFduCYtR24ikURKHt2ET63cTer8
82m/Ehru22afUQyPcnHxtUAE7oZOm6Rkafxq48ZjnrLW3RePIZrgOu3faTjVvrGzeFkU8wLXsyiJ
PtqMieShNLk/VGfDmksFH/rImJ9Rt2HntBwx/ZeiGi2cnYk50DmwAay/nKmCzFaB/yPhqwQiv79T
sRqYIoI28qyxPtwoRay1/qMGCF/LiP3/eruHd0zDTwhecQD5W07/vayZrL0DFMuN3+Zrf5mTplPQ
C3Ka5rfjIAA8WdMvFKK4Bo3tG0ASRo9kvSju1tmcoI8DMU3RGT2txKjfYW0Wsfgc9j6zEAPVfp8H
pLzG3F5oB/OexXkpG8dhnPbHtf9KpamkUWoc5ZvKW9J+ZgGWZwpvtqxdlO/UTDFGHHiGCznATgnL
OvKXs5yXOBQAAf08w02p/oNGFb/sT58t19xQ6IIRbPo9QWADD8MlPBR/GXRxmgR7WPhJccarh7Ni
U0s1YbwrsNHigLPoS+mHOkpq9peFs2UX4uSxLOGK01zelRF24VJv7mk5Wllg/hcvASoO28zhkaoO
yMTWLhy/yIHKur+HYbLQR74RBTx/ZEyZBD26ChtnjAPv/r4KplhVqKx0kadGiMNuGktmHEHC7tnZ
PUsrC+LM4AlC2dzdHynyPiLZaXB5MYcKjNEI1F+QhJU4jmuXTY/gxoFLHEemYA2uFtXEfNy5F7wE
p3iXJr3rHKD6hT5CMLMM1EmytQo2P5siglwxh0y1NRfljpkPLtcoURGHqUO6rLVLfL1Gsc+SsLh5
FwVura3C7MejYASrW429uquGbM1etHqnsgxBd3zv72a4px+c5uIHEfZe9XCtCoLxaIPRUCpPPfDi
U0gvgV5kHJj8XVMWdxMRxwxBosHLk2gRcM9QkBLz9VFg5BPTwNFF8XW9O4KiWLFR/HBKAtEWkjOB
fi1ZKp+ZGTD8R/yRLsKJY0ugx69rF2VWmqxLDI+iqgtSyh8CyOsPVxdaqw7lHH0T9UKhZVSF5Vf3
ONzeSCrMEp97KS3hGGk3LnTkSbR4D/0d4p7K7wsMgXABCD3vl3it6jJhE8uPiKoeYp9CKEzyGT5v
wo7f0Pq4LUptNneOoq7mTbEC4xteBOlSzmJ/RLu4l/g1kQQUwu6wq0DciA+OTERSx4Pz6ob8LeZq
RXuJVO8rrZcD6dEH2rPhUBqNSVobRUfOxvNTE+SfKKtBToke5wLdNnIUl3Jo7ez2jpY6tp5iVn97
DH0a4L6D9aXXpbKaf1c/XHSm6m9u0EovHpaCYIS3Zx2NcXZiUbYnTOn0apAqCYEabQ+Iq6O6gb82
7CzXt8b4uN6m0G8VQcTOU0FVC8JmXG9osvswqnaGmW0cAXTNej+B/7D1waj9Rx4xw1CTwQbWdJ9N
YZCc/H8j8oOLZvzCR1xnjSYGAyejTjhGdQy0KmLSVXrxYl937PpqNQNNZFqv2yu8FxcunllaZIzL
cyO6IS6BiC5+I8vcED6KctCQKgfjUKUpdCd7UMDqaR8Fc2mqMIuJLt5dEiujwPGlmB7FSas1M3PM
BrxxNK+z4NrCX7oNXnVDX2RH788iw/v2MHdGkc5NpsLkWrUEspwnekNP+4BhYqFIXSF7gOrqHxOa
sFMS1LfjnO2DiBzOU+dSfQs3iaClyhhZtA65m44Stj3JQau4FUKnuflRseJUlfWohYQV71n4deAY
Vp87UMV/CFVWW975qufQIrcl20vqSqhYRo59J7KxFkF6Ufl60xlpghOIIA6G2fa4n/cDwEq7uyc3
1ejaNjn/cmNVTFFicbBAHOO5vi8BXQmO+PsrC1ltp/6q+DNycJr4qUA0OUmjfAbI3hcucv+Od74S
4C7kHZ//BeYXJh+lQ9zvttAWzbO/0HxjMwenMWd3qJ7/Q/nvSOs0mLgKvaXon7xQxWqhYhQntAFg
8Ts7Ogn9eybGCHzohv05xJXmmJMVRugu8Jo9AJ6ybBNfukeaZELrQW0prshve2mui+gkTdezFs/7
a3Hje6sMAl1PfsKzudTdC39r4r3tHyr9E2M+tCtdmI6Fya9LQ8wRO9PXyjbG20eNQrR0lkZLBwce
q94wdCb1yG8zfG5NjUZBTNUFHoqtTs+S7IMuLzjWhPpEhtf18fJa2apfTLlnr4CFwH+ZvUlil6dC
1nJ9dyus0/zFVeprJvUB4hopBfo+zq4PHZhwZri6heRO0g18Wfp0JxePhQzREyHtZ39DnCidfJn/
m0KB5LqO6k2q1GDy4+aykWZFnD7Q6VMP1d/Y6CFy5wlyhS/58dLul64ImFwyC5Y4OEJgUqNBvYHm
ED0k1LAw6k+1G95AA17d0xk3AkLTCdJGl1XHc6pxx/kc7Ly0L7cnyhBuJ6UQOH/v4bveD1GOcMzI
ssvr934QNS18uZU340yq0+oC8nHqW3YnmfotDOTmh3CTD5wLWn75uU2GitqRs0IJD5lC77+vDNQd
k5tJTYBf2bOMKPxtHiSLVgzm0k5mTGZB6BKPG7ntygsGmX2b+PpLGHKFvtwxgAO769ahndAQxqn4
r2TTR607kknvdLTXLCbskotOQpPSqv8Drz6xKJhhE1otttlMiaFZZ+e3fDn7lNzGvpraP2oiruYM
rJPgpwCWxwfx0aETlvKJSmb1tH+VYlHxmH23hLocULEjjCtbKg2KacyaZ+e+edVGowXwyONiwCuf
+AvPHzUsFxDlYYNim6a64C1T3hd7K7OW6GBFxBQ+A4Zwk+zUeiK7c83rIWXs9fpWYeHox/J3vYwF
Tw6vk9bPc+v9r9uk8H0mwEzQZsz4UxZ0q7E60f94b1asVZ4H3sbsyzZYZ3uLrdfLIdkyQeIw/BY3
9fZ+1pJGvun2mUz40nqAwc0ZwaafSl75tp8eZDL796Y1SIc9fWy4WEDWYk13kH279GvB0B3EN1hJ
lABGHsZ8ibB8fAmlflVcNR5iXOGhFmHVWGNWex0fQdShH0PcS+k32rGctJCBk+8OdlM8hUK+sLTj
4pFKPd/x9pLOaQG3/P/POO/qfM2CdWoFYZSctgchTNIeaf1vbmVdKGrGIJylshPfKBwT1/uyIM8T
E3ERJsbCfZ8r/4MBQBXuCw9HhgRjunnsUmvCWm4CNUSeaA36ozbwyUkNHxNYio6dDi3onNq42Nnh
JNM9ARNkj8qbAshCnED5ioovXHctXd7JcRVVBYuqPlFZxp94iTHvk7UoCwd6hAQLalTE54AMPQ4w
m2G9M+w0QlSDvzu0di8Iym6bdKYUyOQRH/Fp21EWLWV2qhd3HEirkctEPP2wFpLYz6JsDyrZH2HO
7FLKFVCHw+QpGPLgDCTPX5gtOtmTfNnTWunEySy3T782w8gMJ/HJFSzmFX4FYIY0OwRDEMCPJvGW
a5hkEi4B37TZJ+wCEkpGQB5dZN2Ju3dmRaa2X5uH+Ihz8ZvgWJIXGwGA6RW6qFa+no+R4bxAU4qT
UZHhkVoPm5quL7OOraDPyXpTO7vz9202GsXJO1sKsms65DJmol8XICTgIK89Z5kfga9NW038o7EU
6vJ1ywoTCDlUYVUhes8DvRkFR6yHEfTaZFtrmkQ/Ipgm0pF8StTV1QpRu1sbsq8n+LJo0qhkJEl4
hWsk0nB5U28KOdsuh2bx51bRSPHhkwDjnHO1opKqIkvfQ6FrdBFZsDkc+iygkVEC7jcuHs/PuCzO
weY1fhYyzzP+fLIhtUFxMs2MPIF/fCSzQ8oKpQx3kp14kI4eaVQuRWD7L4u79HniC7posn0oHGtG
hAXFF/BYPA0fBrkQsd+dg0IuSAlq3ZH5IWrgBMeO6lmtYFllR62lhYHIVW/iRUu8k8BQ+mOHvWmO
3lb3IhfX1Z/gygEFRS6vtUm0dBaQqX7Dt3It4ZB9cSC0KbEF7k+48s7WOel811MHqbIkVxxwclzX
7HE3++odz5BYahK5qoRtgJ2kIsAaZYjFJxT3oRxQc6gb7ciuH808YhV7uutOZXFcsj90uMgzDBo1
yBuDqHHUSQW11a/qOE4getFNp0iSjW1Q43+SYKqlwbQ1bzoApnRAq/ujRudc9tCdBHGrJ9kAmF9j
+/m+EBw32lrcxAtP6Du9Bsj6qQ+H1vm8JXwaVr968qPstX2rjNm0wN1yQVvDSc9DuGx9Wz2paPix
6Ck2AfAp0kA2k3acotdJsiEWrSjNU49z/6jERLqLncjgCdDDO0NExIX9NA0k0p6SRGZvdnETHrcm
yGe9P1HkXTBR9B7cUrHkC581DaZxzYrFt+zgAliU+vVDOaokKMPmHVB9e6A+FAAkBQ8T5tEI78ON
+oZPAV7HSkq1Vfs/B2qgdGyxhMFBchEyuzJWWrsBZ5esmYJwrWCXlhs4cMnXNH2Ir5M1JKS13Adb
WsUlpONemWqEg4nc9l2Agby1YAHY2PLGhkAcB2XPAIa2gckvYUZ/elwRZPIf+hOt1dR5cmtk7v8t
MCXbtGJSqiJGHKQ88G8k6U2lYr/iif52NgwICq89+V8nGuZ5WbnS08LvJBymu0BEao/AzfwUzdwc
VxrLV255SadfuO1r6dUbsFOyZFGL8RfDIhJj0wAoLnUa0d4xaz4LP5An6fb2Wx6Hzis8zXSYgr4/
vWMscs4sMPUdRrVlbZ3+7VYJ+qn5q4DS6ZQi5tA19Szbk9xa9A0AGn/jrM3RzpRzYJolnzIbdMbo
Mt8t9NCOJ9S/9E+TmAeMhKj9eTTFp+LL8WHd6+Uug6sXrGj/JPcD+HNzk0nEcFPJAQZrrWrydSlj
4xryeDxfEz/xr9d+xW3aVFVe9uVmYlTbyAQlmBPjsWOtGVwnIBM6xPwOiWF7HyXQHZvBUWDpShmC
Cwgo6rIW8/cvi1cDDXSB8y31FXnFdbW6eNSXAnM68GhaoX8kgKbQbIvtELv4UFrHt2YiSnGwslLh
jwp7ioSmOYOXNVfsSkHS7cJOsZ1VWSs2DV+L/5WN8Z0vPza3t+JpOi0Lf9X4fbm1NEwcPQaxV3nh
aDnJCzU2ZpEwU6gNLPRjLqV2xwwNRUXp3oPXVRk1xooWlS5Y3xiWjR6OdHSArKYnfpH3H+aMw+GO
gOHvX0G4Tr5xbmHbHfYNqgo/0kC1jkC/tAgTcCdNsYO+34AcaRF8otuY5sGhUmEPeOOcMnMmCGAg
Qc+5djnM2eJbMmV2/CKN9NwlEkD1SOKupcKBNCetq2LaB1hxIyOPuxHi8eJ7Iqjiglhv1fXm3V41
t3i+duUZSiY2e9CBwR/iwm5twfIGU/EvAurMP6G6AyJspLSWPKNoZee+iD1RYn7oo/lkE16vuvSh
o0sKvPbQad8hK51WyY0OCOH7iE9ssBdZIs7tUxlVANmmpt7FBuWUD+vvhkls5OM/mOx73u39K2ah
/vBeNW0WDrhb7VE2W1GxUljx8XO60cTeWWjhrjef/5laG2AqyI4khvMrU7xPvBZPemlllivHJnrD
6qaDKdDG+YHNlRxcjA0+am6YNFm0Cu/aPhDvUjYEStjX7DhFlGME/FH3j5810fy7oieAIufxu+wK
9OO3uFU1ytLIKj8FSG1C3YSeduBZZsPcxqZGgrgeb1JAT6PVZpH2u2X+U9Pv7yZ2NxhdXKhxUxWo
LWnR9G/IaCJ3ul4Uq5G440KhSg2O1hOKn9MFVSGOl0pvAh/fgZYExbOZn6ETEDDSqlugAut0L4+a
N4V7W3gRt5jhBeWraP/T57nFxiYyLPeo+A/rQd76LD/F2Ds4rjP58moRNX5ayh4Hx2gY/iVit54W
LXB0lSARyD9D63kyOf5WYuBJwoJWq9xevasgOdTiDW7o5rKwxEEAqdJyIlvre1RxztMrezlHPQBA
5gHvnYQnDFoB/Dfz/Fy7eU14z7o9BfNMKok3IESuUASnHQnM1lCh/Gk4lr3tv9PMhLj0QmLjuO8P
zUvmGQzSlviQSNro2s6xVPHl7lxibBCiAxmmpcmFR4iRdkMB4q+bxZK26VrdX7hraVRuUprsUfbH
ledRExbOvX9gQEkUX7vyBh3zJNIy42KBXT8jCnKs6YdoMZsKK1o1xrzLuwfacbt86JLRhk2Xe8RP
nKVBdGI6AnY0F8h82/nMbQjghnRmn0LodcjfFJJWJE9Ikas7mpUK9B/EXcpLYm/RTaIMF4ufMlop
19SPsc+1PMJ7gq7FYpABls1SkGjz5rM0TkbJ1YK7SQw0HL0Hj96TKBRjMFgT2z7hbW01My6AHCZR
Fub3hB7zbsvE2Qo0ieUVY7IUP4uPhud4gwRZMJLDXOJtON5SysxxNJji9Vf26L1kJjpcXIqSNOzJ
sPzsbXoNwZZl69a9h6M/cxR6gwNYIPFFfxi93t9kvHEE0c3EVOc184qWBUX357ibI8NtNRllUO/2
DHYK3CNRVex26OX3zeN9SRZOFLwfVYGDAF+HU+mSzTAkup8Yro7ejhsOWayhxJySvrSYpKv0NMBZ
pbFHLczFZQwdBIZs9VQugwwrCtkSGesvwnTf4D1nIm5CamPPEcXsrKRDGSie3RaTA1xpazSKRDpg
NvgqRILTBgwWK/vhkQr+rHNvkIG80n35twPBJx8BBhas/UOOA7IshwLJcLejySmiVVD348DLWOvr
n45oObIo3LI748SRNWR4Ic7DgzvdJ8xFKzK0tkeZG/tPNIfHWrrnAB7UEcIoP37qxkckoK1l52ZL
F/WYoTXZBiQauMouSZlmvaSvRcpMUWd6JP1a9Wv/czSqPu5WVpDWFfyQhqop4vt1xl5Fc0J1ozg3
jPm/kK0AszUbdHVI4oGhY4BjY+BaTP9H3XSrWqItww7BIBSQbl6j1EaRYgjergnEPuGN79Si/I9p
lUuMuMK1CrRr10RPj0Ys0ozZHzl8JwJWIpT5uhx+monBAQxBM6lYDNVRqT38APDj8ZtQLf3JoV5q
6tFddbll/lI2LXS5BmJB8V4xUMP84P/7J1oJyZ9L31R1Ay/te21FE/tpJsEV7gWWU/QFY0l+thgh
yP1LLDXYvqiCAeiSH6j+AuD5NgEopq/AnQS6X+0EKEzFSeWNZYOpDIOReRUjSUFJXD+EgDDaMiQr
FnZaXyPQsjmanMJu0vGCUxZcQS8toCB7eUFMhoiKYC5hCSdPz9HQy7rXB0oskrK3loHL9C6yOrS8
RdrLmBqYDuhfAGQB4YiYheT43+wGteN7zRneIy3JpM9T8ia1cjCgF3Kh/TN778TUNQ6bLanZHK4l
in3hisUdTcGpn9tP0GWks7AJMSWUqPjmApnh7Hm6HWjnBv/eXM085ZiDq+yguteu3u395HpXEPhs
1lE7pLraBwA05v/0r5GoL1qNYcVwEKcOw0cg7grrve/eo91WicCb0235lbrpXjlqQiStv2RBzzSl
bzCmOoFfQlJBfeqbJStGLRKEAP6Wa7NRIJ81avumlFQmPfU3ZI6ULrdNnBPca2T8v44RM4I97Pe3
DM515rq/KVVqMxLD2V2jRjQeWFsaFPRiLwSDq9EdfFYPFhmWlI8f24k3ihFlHD5wVceLIVEczTvJ
51tyFiFhNvEi5Ry7olvykMCY+XHgTfLqPNY5/yLUCXf5pO7oiJ5Sn3+5Hz7jZ9cQYnx/kN5DVvSU
eZqqV5Kp5vfX9MbBRSbK+ER9JNeJbfFBSZFrEQjJW3w75f8ua+ylBGlFG+Ymdo0BR7GgWtyTp+tX
zOcUkO+mDzXzeF2aMfSIqH/1xee5oNkF9qmD2JzyeZvIY0zKdN7TQcIGZbAgt9sg5T7bORAM/y5Q
SIrbbx+i6W5UTRB5+z3ihMbtMXMfC7MEiclrQBVIx0+chwHnG9OZ4f9k+HbTbCw39rPDEAJQx4qV
cExaXX5eYG7YiU6qLYNyTKBHN6c4CBuxIy+4iT5m/VwcOKZEs6P897qLk6H3Y/J0esQ4WLIdg100
zvnHTXqgg1/iZ8o5yWaMVxbNa1cDl3s+lZb/ZfhAmrdk8YsqIsTRyTwPHURAbvZ/w+IlmEjPvrDa
YPprNutXj2ITpDiA8SnM6BzdfNMsxibvZgxrHskNAJ0HDfqOdSlCWu+leUfmZkdTaiOEvTtWLjWw
aRXl0CwvlP/sbbuL8lty/8yEPKmDwDfmjJJdBI9Hu64RbGAf4B4APKFyenAflubOwic/1vWNhkO2
JcGKONAJv3ECHpUjhMdPik1LZc3geOnKpKsA4lCe/0+bH9W+lF3M7w0ShdTz0z/MHFkiVMi1y9TJ
mX79tLhagGRUWbuiXnXuYqWCIt5u1vgmXSLvip1BHozZIn7xc7UMNum6uhXps/ovnl84lHUlBtjC
AtsxaI873ZRrRcwmHMc1ui2OKyUDg/KQKuqcftwJuJL6SYFOVLKCr45cA9Dpd4uVrJtbRfbpNDdQ
q8uphz9QegxmOJ40eMRRVBps/w+0hwaIl/V8N2mX8i7u3uUiNCK9nqCXWIgKR1AswIzGge1wU+9V
kyMDcKaLNF9gZZgX5vOlNRKG/6QDZRlFSIUbiZ8f+d4W0bjQYEqae6ar4nrP2ihpYrdZPz06ifK0
JbnCwI8uq6ej9LxXQKtuTFqycJlgAugx5xnWrqOlao59uqsZH7IHcobHatcHHr0WVz4ahx97OO54
UkVAxPt50AgXJmosiKnhApynxuAmU3Q7wCHKMMzbeq/2saut1Ry14TBGd/bXkzXJ8NpcPmNi5HrR
SL8KvUsJce8di2rRFRHAzUI4DqxVJg/7ZATA/z4loLI9lu5rq1M26aJlzcEJgzf0/ZAhF2ZJz3uO
KeeQh7KJ5oZ4lWxS+XUaG5WNv3Mp/HH4+5OTCmEQ32BOAikHIsn8ZtKP+4eCElSEassNuesUW+9u
NTnye7ubqTURycXCrZcQ88WYgQVgDgq/4UzOt6gUTgM1FdYjB+F19HYIZABflRiECD5eBimfP6zS
2dPKwjyvUQMNAd3gQgQpvN5p4NGdDJzB+i/vOPX+/tt9JNq1VLsfIU2F3Zc0GCcBfaXIAjJp9aRh
84oiy5Zcr+cBAtRLgaMf46LtvCIBgMxda7kH+pBIghvU3K6DIz5b1oY/sTH+79MjIRQkwiyj1CD9
NTjjlxbb7nAhJuAlstkPR6uNgLhGcKWsy619gHq1HkkdBE8P4JZz3udzxmvwd7NA3/xKGFxj7tTF
Z/D4mCDGDoqHkJbBhaWkfsPDuzabCsqM5kNVp3t5veh1nhZnXBMYH0FIrBFXZvAOBVUMybXz/Zk1
eIIrKacPK2TwNVmoS0UYOo6lXxI29DiVCbPlfjPuyIri6vQSR8NedxF36w0TqpDalwFmqrtRrkPh
BU4LKssB7sXo9Qc7tBWmaQLEM2cfG7L1VQw216khRaqXn/6hQvckMGl/SLl3YkKfLpq3Lfx6R+aK
0HbOReulwkZaoLFRed0FvdQMCwNV3p7WhVQmkiuU39+lj9+WKnDLmete+K5lX92QtDH5QSL8OSN2
c4gzoacCDEqpMckd8+t73g2+XaX91oQvfjXh9mPMXv/qAmx9S8BGV4OMhRdS9V3rhBk/+u41hWqD
4DIVhRY9Z4keMoWwoQu0KrUj+8MhDGJrWxS64oj91Z8Ll0Gtpy1mOM+ANF3wKHZBiFkGHf73MwaM
KtshCVHTV/surVP3/bNAOH4wlkrLveO0DLdih5ag74NEfxPmU7vwWOg7jU+wHgywo8uA1dTolpOf
gjU0aoxfo/wihlfyapCBZK5PtOcd/NduwAfv1ScClhFpJPRtd2zBk77BxTSVvGWochry/sgcQvsb
VTuFnttWwlr5aThk+TJZ8526YRJdHVYb6gWc2mJBapssHyosm8/vldWvzyqLqF3bx//sshxrn4nu
k5BQ71/Z84fkUKt7ZiKim/mOH3/u80eB+YTWGM0Jxofk4oSlhLSGnRuRyL2fcZEolUYFTTfeqQuz
eXjg5oK4BDwvPjRBogLGsARhyMVN6pJw4GcAXxDMnM/JtFjbZHbQoXrnVBsboX+h1J1GMVxY0ySN
+YBnilstbqnQ5ucqIkZtpeVOwvpK91WOCP2UN35Hgyyzz0QKah0EtgV0XDyj7Eg9GkNUipK7qAQE
/JXY7884xzbM5aa9x4pgtHmIVoywV68oSmPsl13/EO5Ojn5KHSc5V36gXI9NnwU9BKOdqD1T4gCO
0JiE5WZaWHSRoG9sSADTjVetmtFQQOdPxT1Ak4Gs2ohObjcDqKcfuq3pX0xwItDRrW5IalVJfQBv
KVqLAH92lXj7jhvVc25xfs6obb3m76Qe/Y0zrDWwCTWjHWc2FGmGdpmXfrMBTb+hHzbfVk4nlxiX
ysUusuoORnfme8RFdychvFfDJrFW0I7ldW7tcyksoEadXF1V6Mb/f5rYZ1oj6piqqfSXUo4n7W4q
u+Jt2i9ns2KuopH+Y1TaHccHGwPA+ufCf0ccQOTjZKYYR9JTbR7gghA5Ls+pJKtcAkewu5T1GXNY
UmSpdRTcVfFxFbqhcsysFz5aTzN5k2WBjosCIn+gHyY1gGYZYYxtdbjIOC2RguJqV0WhRxH4+EJo
diZpv6Z1wGdCUNwbFDNijoPZNdaGtgEUw/XfwrCkGRjsuGQvBnBJCDnISb3Xl+dno9pDAQo6q/u1
vl827bnaQoTDzMUfNCuObODg5DeX2rtHsN0SOGF7XjkwcYvKIav4B6UQmQCDE2H0mEG8O+T+73qi
5FbdD5RKo4H/KFSQY4fIFER+lQ2EybDRpk5vEdPWgS7wJASlJLBwGAGHAB6VCrIo2/h1cVrYpJLv
QmNMGOAsIbxe+blCkJGKs6rvAU3a2XT8laCBSrnDCwMudJwJ6ddcUTXiCjg6LJBPELOwhh6xrgS/
AJb+7zdPX0dts9Q1BzVVJltmU8sk9L0oFxfaggzSgFPGlu2x4kxbmTqhA/zx0irdMQCoLRZwCZCT
1vBWZ9mbF763LxgG5ko+9xnlm9EqWCKQefu8j2+0j2Y1km2Z8NE1Y2ZSfsf1WUK2y4PPT4iRsZn+
+OzGaw9Hjt6yUnfhrRy5CXy0ZCmmnNPoute4mHrDWLDaujCYA5JD1ZAVWsR4FsJjI8D0z7NRgvKc
qSqRUHGUfvK/TBhxPluXUoLR2wQ2xoLjTyrmIbpu3TXIteUn7WZKA32CrSr3r2TKN6hf7aPC34iI
mcNlsngRzRn16c/vuMBX6B09liCj/ZgsJehv2g5/ZWyqxTPc35+yX7pkfrup68XDAmvCihIVCPor
vY/fzgLkC/IZ0fzSfXwzkh5PfyQkwkKXmhhjUUX+jBBu96kp6VTslMfew93LvqM+xkoH1xs6R2KK
W+Ni03P3sPZXGwnJkSMjwlppoP4RAZBBPL3fyUsKfGIrGSkrzBBVnVReP6QdUCY4eX1eZFJzSYI3
ky3tJpNvP7X5aRl8TNe0I+s3KNcyQOnG3X5B0OfSUVQtkn2KWnLLLzyHc/pcVrIObuYndHDCLYII
rdAj1ih/Yn6l2I6fTIkS5xSqnaMv1KCdvmZy23Sr7cXFP0PdRBkXNr1taGgAQJcL0x6tgnwfPDDV
+fY6xfObHjCq4G5oEUGd8L4dBY9FIMfQbCx3hAO9E0LWVCc8ASSmogpT3HcaY90RF3tw8yk7H6gB
s+WZRQLB4FusBzkaG1EOnZCk/UKR4XMxnovZIPAOLZ8AJLdZFVrbPp4Rl/aC8T3cuiPjP4syqRAc
uXgUE64vUctKxtXswnfKFewrUrBYET8Wj9UUs94TxSIRidpP8Db59PIxDIZz6zrkrM1HQjORZLYt
MaSbcXatukVeaYqLQukZCDD6rnYJfOAtoi7pH81gup6/UZEaJZhVXkV+9DaMsgBpRUuyflIJfkfq
Z0IXMxjMOhOlvzN37pHmMjLsHZoF1mQhcX56IIFQld4V/z2XR+LPyhM4RJg0b+6yHasLrzgGFEki
GZOM+VoXy7NmPiFr+7Ojk30lGNvJSvwyVfD27jeTADpLUDv79dwkWdug9cy8G7tbqEctDxjC7sjd
t4VojF1xSDQYWfnBWYmQs2ijtcqHMnVfUuMAw5Y6iER9OSM/gCOAg0bD83A+G6iteX5TY6XmFbpT
CdEBW1FVEQ7v6d6zxWiy60AKjhxzT+KrpyKJOI8cvekYqQt4fG1nLwceeVicyx/dZYBqAOI5n9rn
DGc4x2FXoztxPgewnGVtm4hxHovnFRcLEJ6Uqy1XWoK3FgyU/oM22sPanCMKynqwkDgb1oveuueD
oR6oRR6ahvDpQCSriIzh27lwjxwZMbcpAePokE87MW0QdBion5zqjEHZ5+6IoVXChnK+VNPM1I+M
chh9l569FZEBlQRgmg3RcSNyBG03qL4PLAcVS8MOQVpfyM1QK/E07LaqRi1uno33pZZgKmxD/1w4
3f3im0ehRoRAIioOHJeVV7diAKiomaesxGxUBX+tMKCIvHPcQ1NRXMgDcurHmchJWBZRRqhxJi7v
rX6lYFWIRLgwsbVkCUWcw/u7ugzmKUfzhJzOaxj55qG3KnUbt0kCzptka2a03GcoDG/m0RRQDpsw
GN0WllPQ3yKsjQzLXCSULZvo/aAzh0gaAoZNbspWU+VY8fLXo1Zh8fakDmVK5aRfQITCu2jCWivp
J4XkkQY4h5rdiE7rvMC7p6EHpwWrvta5nVEiugSYi4U/tKKWsIsDOrN5TUw+ftZt+vwrHTIOitYj
5RipLK7yOQF43iM5Q1uILP92PDnMbIO3CgyvqtPzuFi7qWDVkj7e5ik/hDU3jyPDru+pjPSdLUj8
ZIdzzlz/rVSYgen+k2T+ZspEGeasEadAics/T/QDB/IY1aZS+flSYmH+JbDQ2CwisVw8BdRSG0Y8
A4hGxl0lZGY4Io3cmLnlmYRNG5UDYYRZceu8V9lTbepWYIRr3p7n2Ox3PYjObClOSoTXSUoySa0s
rMfcBRMcMcLEwGwknptfIKh+4/ee2M/vOjQyhhDA5V6T6al3OqxfnuY4luR4jESWgq4MdaLQy85Y
XP4ydxWy2BerN1J7JQLWQqnPP/JVxIfV+OjMWkZa8HKG6b41v59hIE798RMAr4ZtwegT/Wo6OMo/
MlH/RiXvPBvyt7yCgUimDuW04zP2dqykO2s9jUE7S5wCDT7el98j3NmnRDRDfSBJswBzpEOJ/Dsd
1TSYJvkZFgGYpK174Giu0hR1vHO+W2pPbZXJfGePVyBU4vq2L2g4az6vcxvdvsydz6KMJXL71YL3
QKz3RmYFlE80Z5xtIEzkXhzeb6jZfRxMRMsQi0JXwlC2CG+mv7WtzIgkWV3GwwIs3ABUPxGMTdEr
o6FyxjABwsQBMJqVn5A4s6qXHS1NtmzSjXNhzpNQY/RohJypn9Qqa90J/dgADqbs7/b+8rv4PtBG
rf/pCCAYRDlVNumWX9s2GbeEGXfRNl4F1VzzQugtIFkGElAcQuc1/aAVDqi/EMSwc7kPvarjYg7/
T8gmwrn2L2w0uLuuZG0+uWH1WMuI3PfpcqRYuWmAVvBoefwszDcPQGJPo4BoVACQLofuOAXYNbCW
Llg9BlnsXC6DmS0cLG7RjqYP0SAHRgiPIv58iWDFG7aj5LIMYv34JZUao3yZMFu41RAlgE9K3i/u
uJkaKZT9hWpCXQSLSlvhpdvMvdiXVJ0xBIsxST2U6jTLIA93e6wfoheMU9zY89wvH/XAVgI9zvcf
8nZCxhoUzQqrdG1xtF/8CtftYsaMB3VqN/OuClJc8t5ZA+DjfQEHw8S7sta/dPcL4c+FuPRafpVn
ii423X9r08ylVXyQ2fmg8Szz+9mNvfsUTylVmiHk0jjqzFU212MwX27a73rBlV/oqGGcyk1SVJ0m
b9eFC0yN0+2RNxqBU9lMtrQW7XYWymA0rsjqB2bKhCAf/abbx7QelA7awNel7/xuLF1zSq3adypD
cEJt/1MdXV83KdNZLQqcnoAdEjwEmbXgC2ODeUus6YptB7otLQKvASUiqZxvBuyV6K/40bfTAEkw
juHMf05egoUjtqg6qprPQu9g9rBxYCww47vCrU5saMcqYI6JwLNHyuxQ7WRTCjJq357FEP4rWXM0
A9hj+1ebAxV3nBdRqRRXu4IV/bfrJU1Iq4EVidAOrTWnGCW0jraw8HRqcMN9c3uhkC03llf5aSHu
gH9cyq4bVO65w1fUbJvF5PeSJ3us/B9upR+wN3eLzOBDX7r5t7h/xcDctFgUvEStTFgtxZ97sFms
DbV4tmSdC/QgxQpO9/6EGl4gX3BcoIhp3H5o3trUUpHIE2RosCvWWOLJYKM7p453towrJ9xut1rV
vHmXE/UGN7/k3929n55/FrPb+B0dnbAEdEJphk4Fjbm0KNDqcR/ppcmCxa3Qh9rMRMRZ013vT48z
zfLECmMA8YcYNCIp/+7OsGx2u1jvqP/Y+HUM6Kojv1UbZX3W4wS3aD9MBTBN2txwGOCuQBhVhQkY
showB1JMVbHt0LkKoTvppurtJ/WEM8RJUQq2y41qdUanatvEeyUSyEg2xDrOg14FHRdNHrjdsqnb
S6PL/77CnTfs+/+6as1DOw9FHU4/oYzSz/jPeODvuoPMiPMMtBP5DGng26TMx3xYj4GA16paOXHn
kWe9/ivaiw+1qMHbwZGMteTfqMuC+8KTHmM1j2uBVfIbzkHcMQ+Y3AeUej16SOhUm9ELzh+Z/HMD
6DzRhNnugQb1/SzLCj13r+I/+cWENYqYMlrXJPi40O01QUUlu/D6iFLzShzrCxbzMMmULfhvTozv
Ut77lmNkwao4mJSTm5qjSDbSnXABP594i36w34MzkRoQoBHsQGQv0RFr5kBr50y6iVix0BC7PqXJ
cz3Ivzp75RGixMcz3la9cj1M3/iF74mZ41H604bk7883wkmiBbHzqJplb+V+jf/7d2kUfIaNKoIb
/gfHhFF1iaQxdrvlUEEEeSZNfJP6JtLYXSO5LgooVkqW3/e71NllKaoC85lSwAyu+7jso1nDP+Ji
32NHFnbhFjbBHik2gfoYQBZ38TRr/ipQXodvxOamJ/SzTgEshsoUN6U+iwgT5gtr69L8AaP3/jw1
1eyxsET930Bi/yw6HxWg7a3Yqx8zPant1Sz2FcuKEJTWX+RYKSFRZxF3v6pIFcA0zkSUKYCkmu4+
XJUdGhHFYU5l99BhagRakIzvZoyuefu2UlmxNcxdj3HYMD+h04j79CBekvRKNC+M5N1ORTswxAj2
EvWIfYv1ZezYqr+X+O/pgE9Ei3MP3gvj8IKyPsyzKgJbq5I4umo0fQzpFaMg80oYbPVRO2UZ4pkq
Mr3RUN4a2sYjkb3wZGac0GoC2vsuB7jYDIFQGmcdmwujJhhEBeRTA56ykGXUymR3AU1vK1OS7tol
WocXtBtV3gvWEFpUtZR62C7NoVhJBMQHGCfUkeUxBPizUtQKqU6eX9frlWoCa1DPeMUKqXapxuLL
rlK93gWYBS+bXXqcQ8/BLAGpjwfugnSw9Atw4poC3nlaWSziWH+ZDfLYaGbUc3rll/Vz1td8FgPR
RZOlie9LvjqSv7KiIgf2RmHgXxIkGBVVsQyvn43S5nAQkwTqxAd7uqfFXOYvSnp4zagO7PO33fsY
Pk98N6JK4hmF55XIiqWdI7AjrEmA2MqzzwVUbZowdve5MVK+VTcKFkw0HEluvd0up05EPtxOF4Vf
hBzFTjP//svRKPGiFe3/DBq95uaDOVFxp2xQ7h19YjRZ6v0UEgZnvy0m0ucun64jI131Nevdfj20
XW4j7LKJEJjL+SIJoz4//yF0t7yHkTPSkR/cE/X1HnIS0hGBGLfz5fhcvSsw4jmaqIfs2cm/wIMv
zU7LlwvExhtLyJ+iDbn0varJRvrrrqZ48Uta47Jve6cdFkOcMLiz/CJE4MXMFXvPhI+j8K0wdDuw
+KNcW6xYrUK6FcaK8mdJPixdp52+lJ+c+ljYSC56MvDaqAmXNzOpyw/64UxG1cKYoD2qHUae5Gj2
7ueh1/j6NLLe7tCLCYEVxl3JAEB7d/9srprMpVHWqD0OSzBKrAI3ZX5QNIhu6Vv5HpjyTbRNwN5h
1Q2BRtNTQya6kZik+MMM+MBEt0RAx6A9AHgg6nCMS1vrUYOs63MgBn3cmuQNXO46askd+Xd6aTrX
n4uEfS7x4DKyjJOgqxyZFfwaKAtdIjZVu6Vy9NdsekW2Cdc9LBHKrm4Y5qU/sRiheZ4fr/+p/rwU
EFSHknJbBaajwYwhj98IDRHkfDVFaF5ExvwDqTze8D/jO1zq76SMsh7zSA2rXDMJymyRLTC9eJq0
dxEH0oEoea12l4M8ZLYPuh8bJi12bZdlTo0di+Rr+otkEPMrNRvA/mU0Q+d01MdYZwRdhcSnpd3p
6DSth/QO8ZXEGfPwTv6/6V9LDzb5xFHSJyRNdWUdtB40KjDOPwTBRkjZeGeVGp/0EWUtlnn2dmjR
6X8xxhyYaKi5M7zTaMcV3aTq0iqGPgGUGqlACHyXsSVUvrzladGL20D0mbTSTKdRVE4WLwjZH4oo
ylXwhK2CPz+dpwaxs1KPmWLtireR5YUgf7YmGeaymln6Ciu6z1Dply5Fiy7RFp6/xy4B7UmO8EkL
EEz94q1KknI5PbzwolHRg+iuxkmdut4JITZOQDjuoIJPhIgGf4dYES98sDXTKKRVo3QKA33RiU0g
4QRrod69TAIXHh+IO/0xQVqe31jRBdyjqcRRRbIEF92OfrXTx8AUIXGqUrwoUg/wucpFDKlsdjjT
oUM9MkJqU07uM4bIQByp8UmAS06By/U69aG4PAWxSsVRbLw+S+cgpmG6lI83L+eHp+MaymLSjuw+
S5t7UgSpUwbKxz0rVEbLkikCM+PiWPjZVv8QZRVeusrnoPd1WhlSQo14hGuFb7Tmb6fuqB6zrbBX
QizSWvOmvmgvztWNeG5mmx97H1qHj0gfm4q97JisQdhUmaq0mm8A+uY9XJj9+2UGyO+Ra3ZwlSnM
RuccV8+JdN6T85YK/C37x80FKwIWdUd94cphjQoUieWAyu0/EwA4v32Uhl+yR0riuvbLB1Y7L9Tx
7EzYMWcU0A6qaWq0FfnR6uTZP4zuXrjmXZISiGucdc6/ku0ah80a8ziIPXGeIhFkTRd8xkJeuF00
C0YFzYLJCOhNsrlS1c6UeO6mKl7CsiBc9NVhlTKtJFc3Bbxdu91YmxGTVSa/MN+UvF9i4s95tVGr
jS0DRYOzRsRWjpqfPOILfUBh6Qo2oSxVK3Yy+fnqujWF6nXbzZX8R5tlqaUuqzhc0VdHZE1xS/kC
GziQkF4CgiS2Pbtx2bp+mTDatloWzmQ3471/FzJE6Pa9PwjFwzCdT7t5LmEtegl69fsktkOc2p5h
+Y4StlxB/H4wq6FmB6EJlGBjAKgf7p+6VZdc5RDKIqlDtD7U+0EjeiGrNhLIBSdVPSrvlje49wDp
qDKuo7COU/X6DqBQyH6KmjzWtoM2QvFOR4zHPzg4Z8PPGlxq6/E+yjJyaevNmWhRcNC5ZkinvjL1
IKFBNDmsYBbj4OkU4NZHG1zG7p2nRTfk2GRFnJ4Js9NhW49kk17ZDMdoI9XdtmwqzhD2yGHfPMsr
Gy/56cR/LVxW3sPU2RPr2XGJDBRUvdWzM5VOojrSLWSP0wno7GyPvnQV+aeYR1XflzEIhmqxmwdT
B0EQ/tXsQyrh9/zvhWmegrzpxQDz8Ir/uQe9vq894Be9eCjpLDmxPKykVU4PRiqjh6SP+r/kTdBR
V+2euCi7l5tc5P9ygXPpMVivi0tI+XxbKPuUTzc7XClxN7ifR9d0jN3t574vtHdVCugOCBrn8yNx
WpLHfMic1vUL2zNu/tQMMHiPicHqx00PXjVRLB92xd8CR/YFUh95m2T1PMQLRXfemyBRybMpHsxc
2RcYL6s4vi6Y9/3kqscuyNTrIwPyjfCRizB8Kb9ApwsFoInRaWypCf5UgAwHRVz3YeYg3/eUfbyx
gIxbMjZdRNB+bDyqfeLrnG67Q5UbA5IDMkAmn+nJVZUjIVCsDhnVIKjxcx0lEX9VWBxeR4TUuzgJ
rPMQR2GukCqQSS3/tqrKfQkdYl7reSzyvoJiI1UuhkXMPXPNR6GoLAJCO6pWmLNSMkK6Kt89zsuq
aTEAI6dLbeVpqbU9Vhm8Glr68NIRfdXQnCz8ITWlhHLvuyrfvocfV+Q5l8QHUHdHbrP1MFd+DO8U
zjPkCBiX8z70bwmWAdqP78GS/wQZF/w94Tf4GSLXuI5W3j0J8Ftn1O4MfHe0GdYyEWmQ6kc3t65c
LzE0I+Pz4njEW7P+wtDmgQqhhcU7vIDfBEc21XLxkRZDxEkMSXB5qLCxv0PszeP35Tu+CYO82qoE
nDyTCkXAYS9Nbu13AwqA70fFCLB1q7CoZEsX4lDZblKVbOK7n4+diwemcjX1bAscYAo9Z8xPvtvO
JM5ar9EvJlBJiSlb3EOhyti7Fygk2E4TXfh8Hr2sxrVanayZyj7c7Vhq3GhQNyBPjNvoA+spd/bc
Mq2DeYlgmA7gQVDAP23nkOBz/si3WO0S3mCt0ftXnAXU8gX/C0Vxm8tk6iJnyGGT35RaB5goUOdK
qT9mOs/Bv++t6uTU3//zi6y47ajkQDVoGjz+88EgBjAI4DR8oZgvSpi+yPddiwib68wj+OvTqHEw
l8pDdHg3EYnop40Q5nn9ZIx0KXPLvtpTlqpiWJEiIqiKs1bH9j4+f5LvlK/D/U1AgrCzg+nG/zen
hxm9ib4+XsUzfwEBOu2EHIMO7W8/p3vzCWGvkDkIcFYy/nCfOpj01QiP21K8LgqT4A+gOKyFZXnM
TvyZ5V+bHjBmYmTeysJ2RlunqsXJcqE0dMzKC6+ud/9VfNCzmFJTlZSwVs+VJ2EVWz7I5p5OEVM8
xDnlib4CErIwqxANN4WxR13tIEBZ6/Ph+A9r44d7wgPrzoKThFUhkzIWX+Z03nTAsS94e+YmLezd
yM9XW8bg6GHHoi3VhZi9euM1ga0/MY6HjbjwmFnb4zn2C0otJQnXazJBxqzyzFmfTR1YLJ/u/lfH
ctWOtxom7BS0kizPr3ZdaMp6VGONgAzM9RD1htKrV0x02PgprPh2wyezbhAF2Ih2yJwllRcf5tEa
JxA5c4Zt4+lUe5SX7hkkaN6Iwa54yT09i2dQXPurXs144uQyrDI/+OJqL5pJmQTRzp4KREx/x8Ld
NqGk3pRRmTDhOW7TaM0IbbafofCYqIN0JxWIokEjSIwiSyji7f9LlUUtS2Te6Cju7MsHfW3vM19q
NYzcEU05SlCntvwbo1vOVmJHWOY+3p58wCitjDy1XyS1aTT0qn3+/0bsKJkTBiULVWAgUD8TjQEX
J9l+rQLJXXr3zx0Z+PKDlYLAEIseR2nkHKs+h9sTZIKr9mI0DwdkVR1os7XwUVq9Vse8lVhHzet7
UY1efERiBI7O/ExGc+vVDPUHPwj5w8i3ZS/W6qBX4DNBr1+udnGM8nTOsV+c+vvahUd9WY2iM/vV
YA0HshM6Fd2c9+J38IsI9AQxgp/yfvtA2ub3+5TjE5RFP0CESXWTIVa7ZsSLApoSEBx4+baRlBEy
UGaAL2IrhKdZqFjOowWqVXSZ1J0wc+096b1CL5yas9/u2+Eo5Ux7CkjhCHi/OW8P2wXZco/vJbSK
+d+KtPEBtFGyMi+E6ZgWJocmYWfnElzotvYAYOb+rlN6qN1Tao4+5vvKQGG11N8NxSY5YxCdx5xE
orDiS1n55oFVfE1Ow+6xhccfXa2rk51JYl1MmXQv/wsyDxZniIM1JapGFJ3YbxOwk8o/Z1a/jHCW
q9RaTJJZsXKfE+11iRsM0otpCGLGblySGyZfB6cmWJLBKD7hc+Kwr+ZOpBkMGf6iYwsGp4x/4keI
Y4fxQiet7oRHA0guv9GilYNZn/Q8fpZJssIBv3Hf7mXZgZtNdPglNPa8EaTeqcNYZYWZKLcQfzfb
oj6tCjVE6DrNnTapu5YfOJkZqBpi4KoD3AqqynAif5yd13KghCH3kX3Lxl72zCeDw6QFTemJrBIs
0ItpwvUmtzCWzQ31HkQCHHGxeH0FWvOCC1IL4IfujTL0dFhVDp8/lyoNx0W1CPkA71aWq2J2Gg7J
48D4S1e933yByEZE1z54egQubkC+t3kCEWkwl+gplJKBVD4UHfZzdIPrN1aApu4cyOjbdnNOuZNd
LiwfEnb9rOzB8/oZ5HyJhMnz4EDS/hQz4AGl+/Xah6/qnwHTS5Mchwr8t52FVVeurWRXV+5k+YsV
RsHvPjSZfY2yWndHlzlnS/93mkCxEyjfHYwGR+uGgQsqmOWQFWEdtlGp+tjuB20BmlDCEmacS90u
/NGt+NL/oew9tp7des5EE4+6UroEH6oQdp1qQiNDXnDGeY2fclMMTBDdVWDLec1C7x0nLUfxsm+c
Ndyk0vj2aPCvedRt+KQ+ngmKYwS3VGIA2UMxY/4VM6WdbFQuQwwQRfREkDnTKUY5zEIEasahcN0Q
6h+7p2eLgNfDlBnmBmOXnPes7Cq1VmSW1qx1rHZgDdpHfHbt6QQIyXOaurJEuJ4FfVdCUNDSuBE+
+petCinqfF9zT83/axhjc+1S0R7KO0FYUUXjZhXGuvZc32PHTKdgCEPAEQ2IC54/t8r4KFZxRRoq
BNlfKAzV3TyC2/vy2DLGZ+zLO91aYqdRkEeS5MWoII6DMTmV1O0R2X+Jeq5pZ2GBOOwY6guDj3Ro
w6qvM0kz+3WLw41ZJKS5DKjjkkhXoAel77F6qxGaWONExpLkxz34dq6r8gf3VGDes/UULFF4XEaz
eF/Q9MHbFBynPA/MJHA453XyoSmd8ozBT3ZHheWe1iDI3xKfg7cUXuP1P0ZccXQQBVBcvPvt1RuX
cpmVtdwfKJRaosmgqOszefL+Uuv/qXV/1BQU9J39fltKRSXIDwbg3fdhkpInj/GBlQZeXLRfFM5s
9XTnsUOZpdSTplBx8IdE89Bsw5d+TXWR8YvMeCTqN96VU97KBZyROtouNj66TfBpe/qdZ3gm4FT9
J7j9TtEGJb9RP3VitAbNt6cDxEQYWVZb27gQpQOmz52R7uVHHheRTfXtidOoVS/33PDDYSZH4nVT
FK2G6SkW8FinXENZ1G4t4jjW4RoS63eSoCvaZPJpaKrxpT84usuS8OBzFeTe0cdZNk2pdvrUvHQB
mKWRLtpEWJo0f7wU8RkAI7aoANuP88KKNaGYgQRgO1CFHl50UxzOT2ZvFg4REf2gyGT3+vlYpKxA
yXn9sd+VKEnzJ16U6sge3/7VUGIYyVL53nCwcaLpbvIPYGqwRUi9bU174YdQdmavga86uwCDZiu0
x/accbkTJNaIbgjQSiJPlfU522dC17Dw4xLdzztRCifLGeFCrN0RufnAVryxkGcw6wqDcR5nA+uM
n7vlGd10HLjqgSC6hOo/OBKeqRnNbf/BqmvB/qyzgONiTU806U+UQ6zhotkSr1FQlAy1ow9ocwdK
+Gw6hkk+jAocTxOZiP6G62skqkAJB44lJKFF0mohiGIRf5gWC94zkMQNQ/QmeHYscIknLVzsDiVp
VvaNQhBCHyqwxC2cWigEBM+SXUb3gFVMGjm4R5Goj6U4HXingWlln3Cd/V4shV4TWdZa1+scJv1W
bbL7BqZOzb6cuhELGzdKwJGcRLa0rcRqRIUog6fJLCrxeTJD73nQ9GF7QPahdnFMgRuT/06We+T0
m/2z0BIWAqKTgouk8VhjO84hp7Sz9BzAB8uHh3PC8aO+z0S/1FIYZKgs9U4+wu9gxGSw/0ycxyUg
4Uw3W5XcZgYnoXAxP7LdIGL8P0lrgf+HPk4Oha0cDh4LfuiZx/fMwARVipKh893nzN6c2VbczKJS
tRFhXXklgcHDC0Gj7z6lsWbOevXPeAJfceceoEahoB/bsFeXNc4UWMFibvgb3nKNpiFWbSGLtBMo
q7BFGHbACJ8/xDldDpowi9EydtE1ycoqkDc52Fc0mkv9p6CR0fVENMKwiquDR718Ovhz0iC3Ka0J
s8K1l8z226qdwhFQkwXiqilABExHuUljScnimWSwp+eA7oh1MvcKan9mWgL1DFhlck65AvFl4Wf9
TTUYF8kGMHbq0fb3lU3cYAsXEZL583UzpjQiyOyxeaVX9nrvkVlu0aV311UkvMc1BSNnv1lk90TB
TAMPcA6lwMPRryF8vv/liVGO281eZv5o7M66ZR4hj6Os5KHhKborjCCK9o/NKhJv9jq1sm5JXxdG
Y7lZ0FTp93X/lAw3naz0fi+DYiOsq/K6lajFFVewoiNoJmMEcLFtQkYrvmV+CaRZfx0YQWEGc9dF
GJyzJB9p/fSCgx/Qoa4AUD/7pEoqdBV6CMIilmXz9k8pjusTigOyvBeJNskMydo4NqwDOJFnLC7m
mtWllXyf7puiBKhQzeJq0628I/WFtOk5UQtwsjsRiephfqf+4jKeB85OBBi5mA7H1w1QjCWxlopH
BJqNA5GUJiiqw8UxEOMLNtc6z4hj276qpRu8FZIofx1RchKDC092aZoxhTca3dGtNYXWvyeKaHpR
q4UC8qRBY2IX1VwB9c2nRNnmqApGmJl9jv/QzmuIhTiFfbDiWM20AU63uKZdbIcAg1zlfcDJDL6i
ypoGzLY77ohsndfEOp1Lj3ReuLE7LOOA7Kf0pM4B4+xYCQBBr4fUYEQtchPC3p+PbodnVrcu9vle
+G9dFj2MUC1vPLFEY13N5mTHSohyjg7ZY72b1bWrX98bKD0Bnb0zJ4eKkIcwYFLYI/KFpX7nqM3H
ENCRnHFytIr/DBfgxm++kGZD6W5SBk9sSmUzbdPq8zfhbuCQZ9S8TbzhVufXg6OVo1g3H+8sZT6n
ERR3Y1ejzdDnX1Jg0VdgbOfX8VepbSk9fK+YekAoGu8pVDetWfVniY/bi6etNVP7L4q1Xz+j94X2
6kGoykvMEOYJQ1IHB/4kRL1eKAYLDGPcgUmPiNqxX9xG345SrrwILSFjjT4Eaa6Ph67WZ7ZLRPz2
1VV1WXwt7quQzlxzTK7d0LYXBAE/XfePuZyAfvxxRcxpCGu1ic2J+eXdGXTP2X7hitiWgnzJVGZa
5+25OzzymScARa5JxFb+pGCzLg6Dl60BrK5DxBK/LZrVFRyUNv1SBfqeMSriw6fDa69qvyiEx4PM
YsIoav0cyqO0cJzZQd/NyNOyYH+907T5glnbpSJKLfm5YNHl8BhWOMlEjn+EOZ31wtVMcDWEj29S
Qs6ab9bZJsTJe+7sPij8leFoMIyQaYK+jFGfxELAS6dIrB+j4fOsenAFm+EGX9oFiKpr/VcnMg8K
rabCyC8L6ZZViYOa8y0eRBlBV2VkBuecWBglQrWMerXFzTBQM3Nx6203+lcyZhqzJI4I5RKswLg2
95RhPVU4GRIteWAmOFg95Or7WbUeEtxAYVUOGxdIa7r7Ms9VBDYn8PRUCQmGZHtx0tQQEEq3Qcja
uu+rsOTAtzr5ULZmiCQg18rxzl7AV1MSON77S0bORDOz7bbwQ6E+H3hd7FJdthnW1auup6ptflPV
/Uvv8UvvJ2L+pax2vqH7Ljq6+FwV/1acKJIU831ipLlcGUIOmnoaCek2fXiQv9pUHe0ey5C4hPTm
yTnH4woqEGF+f7QuqWkO818oEf7lyCIKvWqZ878Ik39F1ektapcADzrhz6VMnwj04B/odKpjfPLS
Pj9kUB2hP9gfIil6/6alr5ExKAxiWimzG/Gr/qAKequLAk9EcVGLlnL+kMFrPW4LLAx0d2E6A6YS
iLscb5P6VIaf0JkiAKxm2whd7cn7z972h0Ie12Diok1+f2K6F8QtvO8d5OYVBfi4fH+rld+/0B3v
rFQ2OOP0PwnEwFXzomu6JMaH9CnNv23JaTtYozzq3sRYRnyrB5g/LNSE6Qer78GipkzLg3afyS6/
oDOmPjEL7tbsp/YcISKWLTWWehRJW8XtouIeLk5UNkho8KTsKEN1iP6BI+qYkGgsjQeU5S8dFCZc
mKiFOJkK2ksgfW1ECQ8pIFHc9/TSZjtrLyR63IqoOEqAToDYU6QEvcMrIeE/NkvGn1+s8y/JbPTl
mrv+cEMxVW+aYJXh8oq2W63HhzpuNPYWC0x3Od0XHrK0ouPXtTk33su/MXvF6qz3lrx/jmh1qmHw
SWQHaUAsw0fIHPMrOJ+PP0QfoFf5rNjOuQELWgdZedRfO7wCwtK1fJ1gw0LN1YISyhu48w0UEKCa
3OES+TFfMAzDvgQmX7REOVOo4MsIrfHnDQVkwBhvWijNjzKRus+x6CPIZ6g4GVzzCIvZ8QAwGBv6
H5tGi/GaAcjrMd+jgBoJMvslFKmqbJW0W4mBOa9XFJAVZyc2L6p5PogHpKXCvY5iqKqW+b228u8R
7q54osCF2YvAbwC3/JZ4q0MTU6apj0n9tjG9yqmYR0D1QvmDDqPYw3yT5W/GcOBH+A8Mf1dgqqZU
aeRX8wZsbnuLX0894kWcQ1b/AHz0OcVu9OZg0YQ5XlMVpAte4s+oXcxK7gj5shpziUprnKRDUJSm
x1IW99jwa4ZNwhhcOJr9mgB89mc6ewv+nl8uhhRnEdBjYIGjwwt/sQ5iYaVU9fTT60aYGSzEw9WA
cO31gRwl+bwn+jBbTsdbnJzqFrRpnwIL3VVjwbTVGg2pxGoqWZb2jOhOTktf0sw1/pBjJtBM60dE
dKG94hwBfixLoSsrDrYcsReW1WLMEFrdqxFnQIy25FoyKZ97Zi3clr72EtbsjqKajZPkc0cSiwhG
iN/GavxyP/iKZCS9KbJ1eXaueu6kSiKG1OiidPCwO2xqybxVqlut9YS+q7Fv/SWZbMpRFAdYpGuZ
qxDBrRJhsyOK6MstRBpz06aK6vICoB31SPDilwY7+mmprmzlZeY/mhqbnoq7hp6D2V/vEAwzLmv7
8E1RlqFWo/0oKQj8dgstK7sw19mJ2VN0TnPNV+1Rhxn+iTMDzultWFzLFyQlHpXVTjHFK5ffMJxf
hr5TAT7cuJDHb3UAAQTOfdy6/xGJ3rhXxn04AJ8NP+pMCm9A4caQYrY2LZzoLh+dWQIozfrOLaLa
2HPzfATvkVYMFBUPmyUcixro/ZDTdZG0nJs+buKcdgzkmgeaXEKCyI0lSObCRR1PyJ1lSU1mWOtV
0Vi8Zn8cqUD1e0/gxFOs65m51RzcRAwAA+WXpjMQbfUIbUZq/Wk6rfrc07VGUgKNmkZjFe3D+qsq
BXR4LBYR02mL4ttGRwOGkd90K8Ki51AndRUfKwiBCgpCgokj4Aln8zgWIUkZ/yUCJQUQ0g42AgXE
kJww7pd0khCCAPBOohkXqrywwoqcoDqG0NZ+zDKprFcwL9NdzyAwMSmwsADgUo9DkeERtQVzV516
J0YxwbuSBcJGkrrBQjO1PBvk0/ryKuuG4vSWBdQue4vqu36jPM5SOilBluBnrOekbJA3MzLtMPHc
bvRPif39Nqtbtd17/8EhT00WM/g75xr3BIu3xZLycPX5F4b6aFGsH1jH8Hk4p5Y7PvVL+T7ZPnFO
0kxfRZ4D2+LvG7npNjTZwCHlbmWkQhKNbkCfbyBKubYrqelyCl+EldvKyVSRS1aVfIo3M4r6VHWT
QcmQiodQ0IL9zUIVuRc1+C/J5NhNo6fdZeFqQ84c9pJgkKRLLDbudFgy76sg3Wi9tbsuuI87AHoL
x48rFYF79esgJGizZ3wt62kaTKW1bH0FxFUfnp0NCmTZbDfq7ufodI4z5w1kOJR+BQviS4umCCw9
pMkXJZviRQZeXKJv8IgSGv7Ls8n3whkBGVXEHurqOYDnkmc3gW0+YqhlVjN3R+6ZYlWuvEIh+c2r
BkNFDvPIF3Ljxjb7H03Vt9TXIcgudSAc/QwkKTVkV/7HHpMlsHZjIE2vmZk8RuYdKvXbxPMFhMCF
XPXwP6jkpNtf7lJcIHALI2iBvTaJNguhws0VEqawxYaU5ZYXX95YK2af994ChPCjl1zCmj6mEdLL
C8yZpB7VtwxvWSMsV29G1Yw8YrvdY8hdJNyQgV96oq8SPqv29mznDgqg0J1Ply4zvDc43+J4yPu2
SXqs6s+GymIPQXRZydjECvvJvoeIQt8Usj451ix9V6SIDvdQvP/sCc1kK+Pi4trCnvSLbKyRY5tX
0FPJ4dclPFyJ86V8llNC7uZmIcYnwFR/UnpAdAmYtf5665Ptr94iBbv5kwL62wwWEU0HdDDRhOEW
jvmSlg18ngi2D8V+2n6Dv8ksqm4sPmhF01J3DKrLf4WlUcG3d+tnuMNP/x+lpMb8o1Nj5Ua5BUJp
bWqg0K7Ijj0qT4lbg24KpNgfC8V7nvctzKQlRCJhEU4Ht31YATJikjYnBVXi8Lk+38AAeH5fZe0J
RuCcV2PQ+Z0ojZ/tTzbxILfNfUwwnQRTl02sHLlA6iwdUbWuGMouDN+oENbanJSUuGU/YQKbFJR4
8BHmuGLDRa3hqQJvFVWq1LuFjZW5SzRLuuRRhCsbfn9ltGshk222GxZV31TeOUQCEbDpXNNbaaX5
xKg+PtynLB3uNnrvAFAaNyg72pF3vM1XjiFgEYY5mA9XM184B87TGI8SZmVFCEzDOUkWDTKlYUEi
mEGDF9nn7qee8s4/R1kAfUXM6QRI7zqH4WuEm9OhDh/MbxH1eQu8UdQ6dFQVjuIJHJreczWyh9rM
DmjGlIu9/jsdhiejbE76YkvVaJjWo3CdEcdkQGVRhCmqnxk4Qsscn+QJhd823V0QBIfkD1J/HlU9
3e7NwgRQKHV0ynEna4pNYvGZIiLzrsu6sq1yZ41KkYN6XCDzEwyYRx9uRz2wT97MDDT8mecg2o8o
mFzWdQa/SihEFlPEthMIZdjT5pUsg3HEzF5GXANgxCldgIfHbE9643HLgFNwwiemslXrv3f+m+CF
U5Bmzumuk94FrW5aTaBfDaTG4HDtx9rsVGBDscunaztRBjWYTwv9niEE5QsYmnhcIR8PUMdp5Oav
cmN8mbLxZ9tOH/l//p2OF0RiN1rs6frxrRtvQTV1QVWfRrh+D3SeXHNBIJf/4XzmTOt2NiAqjohA
szBQ0ySrLIivNCk3KwgC0y8Ckjh0cyeufU9gDvaeaBo7jTHnqKwV0hrfT+KSOGPCUZDqWpQ0w5bX
N0cihRecDpInB9rWReE3HQYnra5pLcTMWetDEPmxCk6gEhVvuV4WB0dZUgxCY7V1KBY5lCWw6LzS
epU1PLsBSCVoBgUh4UGsUT+k5AuFcnuAd5nxWutcQjjjNtaCiIzBtIAlQEO81SMwMBUYPrkWoj0Q
3P2uoJw4Y8cVsb+Zfp/w+9W/MytQmWw1ObD2jTJCWmSDwkrdjr+Pp00X48ZyMxLqpVj0oT4dnLZE
PSxYECArjVkaMwY4qOEfQroBTFzO6g+Wneja/zrqbTYTTTxmAQB7gYaA7e6o7wpfubKVVpjH8SHd
R33jW64didhjnwYXLnoglexwYxo4ttol43/1h8hFOnag0IBGOLSSxz24VDQqXj1YYkVHyZ99nYnE
hT3ezDa6y+QLZ24N4kyL0oc8YzTi0kRqr8exX8iL9MmgALr/+lWDQRTSNHr46kkL/5KFVAnwlomE
S1GjX6n74vTkC+a8VrxuLXuMNsUbZ6iCj84ygvbySvW7lNxrgsBnwkJPl9v9mkHcPZGdMrflvH8u
T7F32ympkjeZgQ7ewhqSC+jjsQ04Q9AKh8gbfuyI8NAtJnP/1uQNAvjYPJMVefkpqDHcFAvnhbcC
bdk4KF4kzw7iYD0OUmQa9o7tb+sEqA/qHRBtqbQlR/6vH6TpeXGZXMrqgoXVndXyxNu/G1nDPTVB
r1iJ/a7me5g/oD7hZFS8lesD1hl19O39DfUgpnGr4dEHacsT2HB23nHA3NAFtsyi6kVy+oiQajyr
PR44VNyN8xMu4I0haJArVzHVRHbUxxU9V+WRbkBPgjDd4ceaGCpLJc/cwYUVJbSXL+EzwqhKK7n+
E5iSyPaEiAUjCjYTPSUOoWNbLafgLMDBpw4aQKAZwks1dRbVzOef3mnp3TEm7T0CrTxpjUq2Wmyt
hsqkNXJBwJ4EfpODEbsDAv7FplRYsRJGr+cfhfgrCFiolvNXXcduSz8whj+CbDQFhzOcApbR39MB
zKOGf/AWljy3io7HThXCkABF4cctkXbSn3uVZBreF2r2bOXPSpCWDhEV3A8pypqKTkwdq2vrX2Fr
iBw/VXiNMjKOHSofLqW1Xk21CAl8niLmhDgCDTCRMFpCIMmjjUUQuDnN7qRaAbDRP77SY21bgRLq
U8w43DRixyWLq8fxPYwhq+X5Eu2c1uX8cItPQ1HVLJBzBvu8hpbSh412cv6mJXNvKp2b0S/eIE3w
n61QhjTT82i+5Qm/o3dqHkEZr1zQu9WWBjn8+uz0Rs0VZ3iTSjoJzxr9LzBQ6UTgcCvRKNxE35ot
iGB59ksGObwJMBWsM8EG5JQqtTG+W6pxggDl2m09euLj37Ugef/xLjS8SRxMA/tJwKBh8TIY/JRl
C45XdFTiXVqzMHQPZRkPKQ91J8t3nb/EZNyhVgigNA+XPBps5jKFqjWEMXsnqepCdi9ImPxeJY0y
e0JX/mKsgIkyYwhJjvdzXn4gfxA0Zf/Z0rWD0HElbWksFiAku6EZBNkt0Za4V/uYOO1lYiw0TsTz
2Ta5HXu2UDzL2kiYaJh53V49U3OpuYeKc5B/NaPChk61U5fUnjfBM1Xo73DNMJEws2Cu71LtOwnb
1Catkp5Y5RogLkK3i6WgSGafIlsB+oMAKc3dUdFOCkl1oKmThg3CCZd+KdzdWnU5PJ8dhDlH3mK1
1zDPXjjqHVI58GVKJ1JWESSZSWTOXs6vxnGduoHkeg7VFJcQRWW+i/vRzE4lR7QG16F0Lca1sGJe
iC7UEj2xp+V4IrPSC9ESMm0hqMhspGwWmnidjDN2kT1sD8208RNJ45YgPV/yXly7/8N0saO8CD8G
gF5wtsH2szB3SlzsZvcXM/7O8uOEzXzAf3EhEjYXc4KD3ZKGMpcaKVKiAR7XxhSR+e1otidFBXai
yeTiWrn/L+gCfXLz+NokbTcVkwbJZFKWX7nbqPbV0PSY7sdHxG6NmgW5Y2g2cak4As3051pjJ1gz
7E96dGcVXGYzkaiu9HS2g2G2YvPAPHxCxrgRElqe5Z9wgyk5J/1PGbIfsapmVDYxywczK7iP4eWJ
C7NuqBYmPWbSToEC4dimF155tLDzwuAkGKuDrExqsKifZ8EufBTgHKqqLofXBJ/ee8IjTfX3Nx4i
IgVNM5XW9o0LW61mWaMOA8M2ydGknmbAPCAbMfhGk3SfIA+olm8TcQ52SAlAkOAr96wJf4sUzV3E
g+zCMEgIi61OT52iFBA+wo6TADe/vWfVKpkZJm6nZaTNXBl8lvTwhKhN0otYyEm23cYV26Rq4M5y
G8EQZ1Qx4e55I9b5wye+MQgyFuXNcBpu1x+6OODZwzCXlxumwhpRKj73V7ZjruIP3Jjykp6SIeml
EpCE3a1oIJIJgeVkg0JVTMkL9xd81kgOUKlYCDLiountC0CZ5CnepsLDkfiIcNY0b5RZQPt92SS3
y0ItnVtbDhbOFsDNMEq8eWhr0pwhw9qu65FJdvrDYxBVNuf8Sbmz9gYf2jQ+TQQ/rsqloLZdlAS1
61r2Sbi7wcUEeJzl7xOJJlcDD5klAvBEoIE4So/5BXtzseB1uL164VUwxonE9UAzl5z1OoYgxwUq
Js8EDbjJb19AX1D4bDtmKD/Y+JrZkp0PJGngvHZKXFwGjtf4XtU5GntvAmNjDW1f7lKG6GH/X2yt
G3x4/UF2usFl9vB6/IDVKwCYmezuG9+O2+ANO3245NUZ7/D9tvSn+pCjFvSYZDy+T83GHmzuH19a
xu/AGlIYdpsqY9fRYNauJtriBzolTtXHUY0zem+nq3GwkTelHn1sfnlxJuyVsLxECMjecNxqbDVv
SrvgQlW+KH1/wbbvCBsHt8vF3hlbDXEzWXGQqctM6k4iT9xzMIJKORUOH2SrACI0k0SVYmpUY38X
+HA9SmbqbAKvYn7SyT31802uHlUc6Y1T0xtScemfnqQzjLg/gf27/mishjBKWDXd40YAyNRsw1ng
UL3FpBHVvxS8hsSGUYcOAYf1CIYhdTbpIkhkC7dUWeY3f9yupXP6ReAYqhUj7Dn8AUH/cORo/sRV
ePGyEmFL0j2ylJ7j5ADagtRfCPB7f4PCjN4rWQzwXawegBSJAMeghI9LSh36C+F3m4iYjwFTqlhM
B+8Sx8eqQn7oQpsmRxU0DI5NcC169Psbd+XYwulfSyZe1h9ekGlnL9EXay4fPGVMWcHNjcrqLReP
IGf7pSIGSEKo9SdWc0DVHHJSj/Jrv7HjKsIIrOAKlntCTkbHsTcGOrUChK+oYROE3o26g4oj+7U/
jNQbYGy+R1Rjl+1bq0NjUXj+4RiFf4qFQukn4EH1gZT9qYXrXz1Fvn2VrDTGGg0Sm98rT0NoXR9e
XO0MGCzokK66equ8GZcuNIZoUw7Ju1rVzks04ca5qVbjFM95ZYxVzDB9MCZX0wro03ZrEY0Zjc9T
bNlibZIeAmBIrr7HPlTz/hv07kW0DskFTFzaENd5lvTFq+2W6DUoGuWXjAi7O8almlE8RijYqnyS
QOIjfJw49zlfA5ghp5lmjsUEH+dC9c3G6iHYhi4wXwoDt8TYt5ZkSffT/fma4DyUogtVVBo6sCzS
i9Np5PETH+UxSwJH+L93u66LU58CRs2Zf3l3eIgII/F8AzisdVBawpyx8Obd4dGCqulRLfA3ng/b
STvFMy8L7cW2gMKhyyqhZJD6IgBLxS14sbh/LUhHpqiTyVOMwKzTZB7fYK8FAiCz0FX9VQhUmhMb
IGr1YSr1JzLurB4bfQf5JIrBQF8Z0u4xiTprcjSiiTtQ7lLxTKIKK9pzt9eOTuhPkcmS5OCTFVF7
1W0qvqSm7DMZE8iYtuBcb+9zDw9Uz5eOyNxvXD6tAOP1pHHSV5VyCOsvG69rNtB7OC15ZM46fNLV
Su9uGS3fZyArQVMqgiGh3FzJAW3BmXwSfVYhn3RQwelZSjcgAGeY7kF5ZhakiF0aFiVhhC3Q8NFd
f20UgHawu3rBUIXtSQ5AYTDLS3xBuM33JCJCRl270d9nKSdp6z3lGULnRA6pytOzHRXAj4Qerfjb
/R8F8+wYXJfsW4CWL4C/DwcAjsfkw1+TMDmhhwZLpx6HBO2jszyEEV/+ShCVfm03i9vy3NQ4htQC
q1XenKN5YBngYoK11Jty0vtdSpQIcL17XhaAPUNQpJG9WT7ibffnECQgVjmRS01BafW8S5/d0TNj
mt2bbuMa6TFuAVwdgvGmqubwYF2YLb4rkwqocsjR5TQug4N/RY9pq6QBcHzQ7i+LmTTcY6iZqwU6
pYd4j6RmonWCjr2f4JICejPmcmByySfFi5sCn/mwkeiCZF4av6bOGYNhEfL8bbiv/SI5+a8ncMBY
5NK/QprDCfOWCKQeTkTjHJ0q6QBpJbomCUABs7G8XUyQEC3XlQvSdIK88vpO9yaoKFU1+7VkRJJG
v2B5fCgfZS9cC59SWSWcb9YjesDninSHMniL8XkQkqOPyW9FL6FvwYOP9sAuwdNspmqz0PzCrFjD
xhX7wti9VBIUgITjgyQK6r4K6AdluJA3wMURUqokoSDb9F70iD5ACsW9WCitUytGjaPLVefpWMv0
vlXX7DSVArdy+2Rl0eO78yPi3ITnq7DQjm4jLLEWYaoj1O7nldR+XoogBZGJ4VJiB2iJ0Qc1S4rH
O8cSmpjCFRVHt5KzrVaWTWsn1RPRYymdjH8du8cgOtbBXORjHd+nd5YtvGerenW+fHx46abFMcLb
WPOQLdVqaVXZYHzgH/m9CVlLMcl1Fgec3Zk6+GAUABDWzPMdyj2tj0N4J+n8GoMT0LxyCgZWW2hE
Bqn/VVZx3e3m0zJejE5CnCi802vGzt/gZqSiJzqxkWJotOgifS5VSyGExISneZcmiPlhJ/UxiDe3
8Y8zYsmFa3k1No+AOU7neRvZVNF5H9Bc7O7dF1wsFhTj1drz4syNM55IB/aOR2ZyTLpPGseIz/Ob
pdXJt2ra2kbdws6pkmcvkjYKvfmMcjfyaw5y0AD1mgfTvmmgm4M8PwR/74ea8+XtOMdV+Om/R3bI
CAwtwyCLomxkLoqWCwoaSpPZVcXYQAO/iwjUlCI4hdow77W1wdgYQePAAESY2SkiwBnMOdGPgRFM
qd/bhsgn7Z1twq+nXfyyGYB8x+mquXKBLfd9xOxKkPN5JjHid4KsTpcKg/gnTozUplXl0Kctp2kS
iU9iqyGv+P3M0wND/tuPwC1zgv7eBqszS+yfMj98/BN0uV4x17CZ6gKLF/8vkzjv0xrIBqZt5U+5
GaE7Mm2jngMZiQcha7y0y29ifu06bcE1ftZpBxIEOn2FDZ3rx7WLNBvROQIldGoi7mv1Ds1PHvy2
deE1l8nXiHB2KtelMsF/esobQ57yTM7KSNf56xyy134E1pEPg0SRYOQzxbafP7wgKc5Iu2yRrCjY
RrmYVd3Z3Q0ZHvnE5Hdx7IA/7cC4NMkrCgbMj2OO6dbJE+7XiQ42e4rt6VyhAhDThLy2qZ36y9TB
h3FeiTeYVieh6SSKZ4HDhyewkiZOyzxMRMs792HIDcQno8VsxR/6sxGVE5YZlz6cUTOdD+224MX1
e+m0UiANorkhh56ca7KpcXV2aO2H4785i8lP3ZafIWxk63gEmKt1uk0fXU02qpphyof9yK0GqhfF
w6Tp2EkkMVcoW23+8HT8mXjLfZmvI/ARO4mrAoPtSWtJ7yYqnjY/UZfRg+YY8Hsf+HEZ23LST/Mx
RKoDQHpHBXU7ZyQP07qV+P+dlUZn3zLxGXWhxypbtIaZ1f9iHNz3UQXCG3wGqftDUSxqgDeye+SI
z8NHT+GK62c1jvBPwYYIqpUPPpc4vJ6Lzi20uZ2dM1oLuL3TF9zMVdbfkQnEw2bHxy4LgiCMCAqR
GmiIaFTTqbfb2QzfbwBtAH9zkL9ABugJUcldMCj/1kQodORZG2KTn6Ne8FHTrcepSsfWSi5lqyxV
KfReN/tWJ+xz1jIsJkIAhyUejyaM2WAUWmjiFS5cTYMwvnCDnQUtbMLJzDXoWkB6VEzIi11lWhaZ
CPX8H0+cDUCMUBnN1xUHCgff/6eNE7/Ky336o3TRcUUCsQO0+l7umtFj+Jb7hhxRG6gjLIO2aTXf
jYvJi+yyM6qbm8No4/S5SUbo9n2/4gotTtVA1F8Fzk2uuZO1RnTdbWlbvRW92xqTvhyjtIMPExfJ
45lIT/uax6O+6JE1Ws5b5BJxHYO8195HbjiMKoUmiDxf7S1sODhWCAu4U0HSqmkAqEDj5IhDT3BU
qkSni8mYSGU/OOCkgE9/9fkyjpKxHaR3YxL4nZhcz57cK/88LOhmpGud7KxhAat2HGryewrggqEn
JXnVg61Q0F02ihqiW0t8JSs0ZRGkUUoCoWev7LbxQUAXqEIsQaCeeSxh7/GEE4UjZAaQONxctxyk
fq1fbIbBo5+QN17uVuEhEZp+oc8WT/i04U8sh1HiDJLI0PzsxYccN43GpuWCdDn6OZeQoq5A1GG3
w33Nns0e+Qx9sJmMtIwKs/DUZTq6vZLvCzLifC4dkRsw6XhIGKSUBYmlZrOlBIqnvjAXTnnuXNEE
QcP8k+JKY42LwlOXgI2Q4vAbAQ2DSqCORxU5j1rKIE9jfdBnNGQY4tVromg64RaDSeXjNHzSVCrc
juCpGSlSA5A/bHa5e3HfzdgSYXPLBn5ouPJs8Zon53uy9kJjJa25rwcvM7L6xAIfbCXz9xNwOHCX
+VBO5YjD+o9zZZ3GvulzP45ko46kXw+jLiI43vfsgmFxaCExqwsYNs+JHotHOu0y1AjbRghzwXNB
WFbyafY632YX6VWDCVrasu6hVJUEQVSjsIzY2F68uL2Jpgajcw0kTAjhK007thsV/TkVV/8OzBrA
HHn1dD13vOan4taKUEQ8GGIadrYI0eXcS6NEjI9RJ1F6Ty6PR7NNeyl6KytLSerVaimRzrbo+enZ
8vmII04StCBSzMYsAmLdBtdgeLf+nPq55uvJu+yQlpHu/Jzshya+FcimhphFtTf5IAlVXd5EEhB7
IjYakBfR1lQCQ1EiTAaANiq6ZSPSAIoe+lUE1cEKgKNoRMx4Ge3fwZ7Rnf1gFg6QaRVDp4EPYEDa
lz2Hy4Dx1SSfpgDmAJqu/Ugu7/MQqYvC6gWQaqZOkCEa4wZq6PFQVNo+KIhsX0xIwDwIA/J3Xp62
CTe5XLnQtyYTabQCR5UID/Mou+H1hYXnceeDNEbMSBJQ1TxFaUUR9n6ztHCEyAgSBBmgFQ6Pibjk
5ShpPMUzw7WBt3zbbFvjfH9WDEW7ajq2NKxAZlh3+PVgaHrZ3I7ywYDQTC7cbzBx2FneuzpMlMym
LVHrRhAYwvRkI4oFGZgGCQGfyh5/3fqpVWQzqG88HDBZvYvkR2i0xlp4Qgdr2ymThULb5JUrlWq+
+6I/PWBM0cfFk+2PKRd0McOaTHUi30owKkQ/6eYwjp/zBIGWrLznMzpQ5tpP83XLJ49qgUhPdAPg
iNlnJAWbYH4mCD/auqNrehqRaSERvonnUjLGzWepQvTOcfb2gIQ04p38jIjd3nmaq5LjwKaM35po
3/vE8tEl3lClotimWIGf7WKVwXlsG+NLit3LyoflupGys+4wj+4iDK7sKeeK5oMKrh8/rVw37zHC
QzmgqojrvMe6SwkUO+MUjQjeGv5WPMtS/JacbMXgJXmnydgdpXGhwaxZVckl7mfbAXzt5fwZYf/U
+YGV65MMhPAibkpP6ao7JuRxLwXwLKKzG2nd7jFog7s35UgbsDiSzF/I0KdtM5wmwAYbO3f+1I35
++U/z0MdAcWy1aOqW60FGydSsZWoEm85YE34aLIrsToMW12DdnON9B4bSt/KT2HHqXBHyArIYNhH
xlZGe0/P5t6y1D8rTHZxrvv05OwYexE2b1wo76ssIZjr3DDrsc8bf4mBn1SiDlOlXKzp0XaVCGfl
Mlj/WBShf48RXLcDhKimYgGhCZErg70jBP+ZJTrKtbP+vH14hNxMAThQJMbbH7PgxYhNpzLFBX4n
HbPfC/lO5InyLjcILkzPPTSZ2HVzsRdRXSZSUUm/9IHFM653AV/YlSu5eGLF1Uo8E3JmVvcOLzL+
HhWvhQ/u28ZBzWHha+syFv2hreZCBwgaT9o+3XiHWyw1rVddouEssu2PeIliq07TQ9UCtK8G26pL
QQlAsDAwRa8S8hJYJpK4PP8wT8rfHoCufDC1RgN5wDVL8zy2p+jnyuDZV19PraGvya+oYAGQkwIU
S0dj1G9muVtbFCa5P5FfzTgmDFrF7Xwcodb0R+HbHY49//IROqH1l9KZVVae/uESGLyFlaTlzZOH
a0z10zl8J/fImEG3veRIMOS/hy8Abpk4P0r+2IdmPxW7Q19EVFzOBgvvlHfHBr/OaTS5r9Taz8Uj
RdTnJQM8QbCy85rfqf3AR9vMBqt8rY5DZ9hQy9FLJZrrgxlZDCyZlkSIRMz7sMLKIfIc30WbYFIw
hjNUWCrElv4Qd+MhkA4+VAbM2avL3o6vGZbNlVXEYHv6CGbwO/5W2C2fadvn/hsIKe2KdGRG7dnS
GoV0EPgmPJ7NbM9dH/UVekzWQ5/6fIMQvD0uys80melihw8HddWuD0u2k26/f8fOviLxcc15/Vt4
MOAVbJg04DC0DI68q/kz/1h00tVcFYz4yuWYkSB1zHpTg0a+raypQKog80D2GXTAx38PnkPR75+j
EQO79EtA/2TAujWyAUK7EJADz4kMpDYoyHvLFa6VVbjwTzdquAY0Rk9lNevl5Cnpfr98siF/VAq4
9sGwzWMpXlmiXrrA9JxKIP9VdHslE2XfZ41Cc5Vn0utDzHHqfrgvaJBcVPbbiYfPvp3aZh4WUC3I
sK/FI32eFS22NBN961qgvxiGJG6Ix2OpGfx9PbWdY9SgsBJv9ytGxcuWk74jsPKIXjHuTj6tqYFU
NvLAynnW2PP4AugHEr4c+B197OXBfcGo5ZrXOapmWcysn+S1kNSYqIGY5TuvIcTIR7nENrIdeoDy
IOaHQ4wvp+vji/YQ4TgOebWERNfGO8LMHFQyum0UtNXUnBRUTPCwYh275ksJahuN00HIPxrWLqpx
VottfoSnWzC4v0tDi2jvDXsxtJ8x9LF2AT4tg4Fzsd2/vB/k6NdJZiFlo2tDvkYP9mVbF17sBVcl
zmH9v18E8VVm7rcl6i0FsEaULhHRgboQS6HFU0RPak1MGxYytEAAHuYYY7q6tc9Fd+MKaxYNT57C
fpfIUYNO4vWkM+Zhjg+WxOrJqdHgWtuL0YTD9nR2D7LsphILU59e9EkVnltXnQ3WbUjNSyaF30gE
jcCUUO8k7id6Xd8t2SW7vsPWbS2I5nL00o7qCJjqdki8rZMQqO/7VWxlZJ/0wSyhY7HDW76L6rdw
q9fAYjjv+jBmkQ3BHetwGeknzhwJzjqN/M7eUGdCBD2zGir9xN2AbuC/vRuA5/RcN7NPqx1Z+ED2
UDrT8BMuqU2hkqlq9jLNzx7wYURUaRaNFZ1dUHCCsO6v3sXYaYr8oHZnHkZh1zPYQyhnLN6+E42e
//GuV8Am3wcnoGX02ust0JAY4VzxzXPAkU6SJiJf8DK4emhY8Kjw+vEht6ro5utfpnGvp2NHp0Lt
PmlHWXLbfOqfrrNlpwNW9sgLkJAeT336E/1Qf++uhsBjscIAH4L6fGW75/qXY+absXTdqtU0XPRq
AgEYbBqjlNweJAurdVBS28nuxDgb8nmj+v0Q5EKvWn5AkERnGM6VPYHaovTgWtTvyptbQgs/qXNr
0g3jbEukRq1sO/IVAi3FsMLf7FsjCum4u0q4yd15U/RkXTNar1y9YxIZdLJtFPc3tzl9/Ys7D6c3
pEk1v4b8VBsbw/PxqaCegziWminmmc7BQ9gZtzit9V70TpR/+O1IzRegfHPWTjsmqKHys4B8kypa
7jMRASWVWL6BnnDy6SXNJ8IVIgCyaxkS3DFIY1i2B5IgPQgibe4RPkZPzIqrcqUnYHidNGFIfveo
gm6pX0YqkvXrNzi4McufJ4eU0ffsnuy5NazItEhSIR43Ila1rd6ZsVqKjwFdHgt4m4+pZgeM2FkI
d9F4hM8p75rXnoPNM5DHvddRnSmN5fJDj4NUlw8urYcP3q29g7oX9XGBoJrz76iUnzKKj4olZho2
7KS1L2V5lmB8W1jNRddiJ+cavx+jqdV4LCyaehIf581JWMxMM1nhEtG/rK7g9nAKQAbbwhm50Lq0
c/vUGX7Q1mQJNBXCSd+Z/CyDuHj4KXHC8i5Kw3BNvONKDvLbQThVmoYwP+9tYDOkja4ZHiS+IOc7
cZhQM/ZQds+mlvmh+qwHHwsqVguUoQY4pfMRAQrxNpbASiio4Z4aUPso72VapBO7tFJ+lIf3RUQB
PWg7K3Xl0fCTS7WxOx4altxf4Zw3z2VM4rtM+JVZIATzsFCy07QVha/XtX26mnAD7/yH4PwoPlXh
2iVuPtbWJQGLLHv6PnTEdN8X3zfsDd5DzANzQ5ebGkfszqzO2e7XTOCmhx1MG928zNo044iCrW5Z
GxQwvErSYoPMmmqAsGpDeoA/yS529xFFrsL9t0YEHQnnRk09j1o4rCuIX0KxduEojSB+vRFN4w/T
Q7ymeHZA9WTnxwl81isOrTfTKj3dAW4wer3UyC01AIFSi1tN9AM3hycAxcv5JCYVHn2lJNG5mRDX
iGr2yX0h//eqlPLk2cPVtqUbnLVbaQEVfeP6xHDM7Kju64k3Zn2ATleTK7nZtkvWFdsZs4jvarjL
ZnI7yilxulpbUhYC6C0h840/bLR/0xop60OiAzhxhx7ZKeVlyymX/FP+xQMleCbgNmC3QyDTDNV7
YDZpOjppaCGXMbUjlEU/hNkQ/pNYstET5n2C9Xn8eFoYZP0fgaVZ84rIfzR3YjEIBS+f/RxHtgYk
vhM2mHotGv0/YvlFSNbHqaI3CHbL3YjU9KuDmeAXGGV/G6pGWbiSoMiGCSsCaF0shctSVDL4BwI3
IAFr4swXXeG1OyKOCWdrbZS5MCmBSglEeOVYnjogxGbvbovV93BRhL1ihjKY2jsqjvnEJhj8mk0u
4jXeBAgneVzslh38Fz3FFgneiO5Kn1YHbqyz87xkUl4QKxkAVSmXrl3nLCIyb+7eam6KzTj7NoI7
LddufWkjtHT7xm3O/y47pzCnKeA5mT/U7U0BRimkvvV0UQmXWDC3tpTV2hbAh2Ro/VXb9nwv2C3H
56kf51Gf8WnvXaw9L9Mx8uo3cLAt+Pb4xDBzXaol6AZoA0bUfd0jOP3I95hQHtSGgNbp5N4F+Zza
vP0MsKgtx96zl6R5qOFAwSevJhSqkgMpWOuEDxfC+yjj8cK7/h2WYKHfmQHauE3fKp1+UVtUYphL
r+1S16u0CH2sMrzHJ35ltWsjb9aVxERfPGwXCo4K+7zUP7fHbi73Wl7BAT4hYdAxtTKi19BRzFeb
GTKGwzSDnxOXXSo6dwCM48XQJxldeKPGkcDaUf2dcB1TWaTZWzQCfWyQICbZ8/9Gxpe8N2lnnp3u
weSnqQ8mDQ90HBHK7OeYK2sIpAxSYt7QVOjoCWKwx0h3PfK6D/kQP2wAF3tXg0IisdVeSxjimGBy
p73YtUIn66yCykJXbwZYxmehnL006KvRFZCQwvyusZKWMn0TwgTZjZk4zcOw6DsYwdGQyoAMpKi4
V+mB37Gy6LdMNMt4A1pecOIxEA8tC6ANcZNXkeFxf3OZ/jmL0fPoFPM3yuzvobD70VbICrxXrNsE
dQkkqj1iqjZZlM5QDzdqdw7ewFDy38OqEy0DYCjgsS+Y7AVUQJqo6RMavd9ziRwaR1j+0Oq2T+Nx
GRLMox2U7mGVE5+HckusC5rlH7CdjbNXXJtti4hUkC9UDqN6zsYVkvqXq+pbOznot0xLbu3Bhgh+
SVral7kEGHSjAD1OU6zpPCleTovLouw/O2eBG0Io3gr17qBC1AbGV9y+UalWKlWJEmaP7XQ7Kscg
tMBpU+ccwwWANQ20o9fa6JmYc60Py4x8IS3ZR4G0gKIRGfwQe/+XzODaKjzVsEjLv4EDMnER5a+Y
Pd4ng5JYndfd04c74dClv53EjlXvi/4tiSOINeTGja2VIpkMvSgQRnV4UBLEMJIyV7S5dohMWI+O
mYJoWDM+eIe+5ESZpHOQCN1j0HA3K5rOj02MyV9aAx7BN0sH1YVd/WbLrBQT92Wsg/1KMnScLsFI
fP8gbLZsI/8dmVFGtSlmBv52NeajdxQcaYavzbdgc5DIGCLWnA5A4gADHNcmy5+uGK6TaTe8lFFF
1hid149l8nvFKpB00H583raA5+bRRqOl74FqcEmJS4ZweAHoTCzlmH2hYP5aZtnTVGirYpNObSIY
GnPPBwG7S3XQ4W92hFQsfoCBQt254dMVLJ0DSX1ShRKfqYm5xAS+XBS5hOUcZL6QzQfdPliW3bDs
gCrkGYNEvM32aNOVi6kaQ202mKd0NywOsaGJQ9SRsOXTltqAzhg5q4XZMUy7DR1i6Lx5oUqu1DFa
9DaWpolxV+yJtOORwpUCbaRjWteNZtVArFQBpvsb9FGgAYtsaR04NW7BGkjPLNkH3xx2IBXjZNGt
6aNFIbuOiwLj3Sx1i29OpFKja9SpMTZ+j+ulkiRjgXxAsOm85ONiWY2Z/nU8qk9Rga6xmdnx24QK
HMfRlDVDCU5x75eH0Qqt99QeT14zivB/0jYE8OFAWHFpMH+nMLdwBn4eVSGxeKUZCAUKwxlSGs0S
4hU5AKqi+45s/u4TvFmoqZZObPoO5upNewcBqmSGIrtVB8VAcyEMRK0qGMovbVhJCSk0MFcudohQ
/XnMB1/uZDwZH1VnH+JK9Ps0VSluNXiCRExnnepNRBYRxsnq1DtOTVtRaTQwbpWoAJlv06vxta/G
ABwf7j0QD3lCq2o9K5HKPemzcrVJ5Tm9TKZz+rwQzEAb3jhOilex754HIM9gzPR1wHWqx+XfYJAW
EM8Uspwrr6tMuh5+LtQCmGfzigP7gtmSawOwc7rJbuik83xh0/fhQeFNBPcLgX7873cnmJh9iOzR
lMpzNVKC9AtLTkiLvREG40ZlJ6hIEMMhwA1V96ccvm7dw4ZpdCYkL68dY3JRuEHGfQBDSaKEJ/xA
kV8xAyjr+cAR7rh+7RrWIWk0IQu+miBkhekh7lYTsmZ5Zw5LAzUuZIv2k9zAqktj/MkGK/EmO3s7
a+QZQ8XfIqnoJzFrwkNAcGtAqTRAu0t/6SAjybVW2p+GSxl4xpqX78JAxCIsloXWiycl71RNRNcM
4eh3Kcpavdcvaofcx06cEDeQmAGbGsM5ZhN6xxi/I0AOrMyP8Fp31Lcvh1ktde9vaEJhMg87cDkj
ibg54y0AWabls80WBeqiZlM+Z3CCQfsSyeHugm6RXpy3IQcLGv81yQSREwJLrUG3pmYhi1BcSDYs
gyfPHZbXGyoOtv6ees++bRgr4Bo2ddVHsfhuUWJJMLfltuXFh0tyv2oKzNE9mUSCCxZdkjJM8Pi8
xYuj63TlcivJD942sXdP3rgsnYMblzhW7/vrx9kGjVgb8q3aaSv7v9vTf3OWb0LGAfPOQgGFr9yd
/gbuYhYmU2Mc3CUOnOvkl0by7tYFac2JLwTjEENS8eS+Bfs1I6OSWxX4Irt/oMPQvKCEs5fs2pT+
z9V1UocBniVpHEoItmp9oU3sw4VjHAd8ri8Ridf4Y4rwgy/eK0/8IRX636n3fcZXOnWql3fSeYqy
XzY0mMLr8jQi8lTUFNn4VFMKXIIhkQzZGGxU87AzrSASpEp5wG6gTf8BxK5NpT3DXE/fTv/RtqQH
2BNVmsRvEcfTywxTltQVbf0KhNMCAIsHxoqv+Vg9bwhP7P4joRdIv2VGjBDLCxbfmmS63YLEDdBu
ONgGmolJlDgxhXxtipJovMaZ3738VMEC6clBbMZVOhDv7dUGjNnzj/rgX9gNvcdXOC4+bx9LdW9Z
JgX1PCAbUwZvyji0bYbRvvTElNo82a8rMt7KhoKlDKRO07i2sb9LNcb2FgP+EYFtGwIeTMk1MO40
UCatQ6TDPPWW0wZs3rnEQnMNJv6NEJNWEuT/9lWSVSnH3N2Af/sN0uouabalUL/w7SCj9EoYieXD
g7zAfV3gwxd87iPRwt2OCCi7H/MuEHUfJvH9zkI+QnY5v8VJjgmTFOd6JDpAZ8YtM4OSzrw71IIA
xrJMNOH9RsfQWZkuMk6pRI6KATmsAiNIJeOm5Ey0kGf5rgZPMkVWukxDCUkHe+YVhsUBvxoT4wXn
eb6YjmbYt9TzWBuLS9MhYrjeq9T3NyJ+YlJqIeHglAI8zBWdA9lu1jm/mfF0rCSc9v9VEy7UWh7E
5SV8LB9gZySJS85FFmgQQJJeFNRGh4u+6+WyZ3TCzko8ozxgPhetq4cc1Mc54LOJE4VFWFpzvNII
UMvPr6kEABDmxUOUlEpo/kooTd1N3k37uU+U8HJJWI3f6wFE9+x37vLITlMkEiJFmWAE7xnCm99W
ylscu4X6aPLg3QGAW6xmL/oHtojdLua/qIGj53v4lMl+yyTlGlIYwPNxUebVmyy9xI595j0Orpb7
K/neAinxWZTYIXZZrNMYXTX1qoSYXtFiNorcvf/Tu07TUeEvfLQVv3tXPOFWt4e2br3uuz9moMK4
b4nbLJRVfEn1qf2lDac0dO59qrGHZhvV3crn5RDfgXeh6khm0X7/KoLEeGdOdnSHB4//P/Er6e1s
z+SggLHsuSAKsR6NzEnwmu3aD9zRkcWZ2YMyRohOFTI6gbFPS+jZXW4NLr3h0+0lZm6d6WutcRne
D3HGJmiJ3qwGsaOl1+moL3Sztb7Sn9lu+gj41XY6EkELFi19gCNSgExZn1ZiwCXl3LU56lsLSgbS
/18CBO6DtGL+hg+5MgPZYs9PLPuBYFA6ZpCPZHEG6vJAYlpOlGzKREeZOwml4POD2fisqQQIv99B
ZWHCgC7weLYC50ClKB1IHoXlpIpp9iJXxKJbXMRLkNQL35qxFSj2Oqg9goSD2xAakdRpLckxOTqL
djXlLM+mHqLkE83Nnn/ljL+YnRkc6GtW8/3U9asV4Kqs6zSLo+bDrmpPu7QGWKxcxawRTRdaLFCj
WOK1qMcCAex0qrXPa4l9p5Idtsfa1xc0BUOK0CaUBhy6sR4r/Im/MM+8Xn5Y54D9O5s/6q5NGOqR
IQe5DLEgV0V68azcX3uJ1tFYbm/62H2xtx0Gs9NODUw8Xx/26Zo0VhO8Gq1wAB1gmXZKmz9X2E5D
4L2f2ZHDOO297h+kbQJLqNUPJI9x6O2E9ElqlxzINAhENmQrSRmtestQ6hR1LrShJ+kVSYtlnb//
VczQNS0i9UGPLwyidDZQFQhGgsBCVUqbCT0NS08wrNlFcd1FLjisVUPmTyUX/3TPrsq93sJk2z8R
AV1AFgaChSHh0aoE+ifqZ5J4NG8daN7OmbnnbBqrspCNty/A7TIm+GA9vl27DYflQQr4D953/Xss
3Sg3tYVzvbPJF2mDF46E0SvudeisFvMsh4A3LMmk8WzZPEjHqmm1rn5PudTQXSh7xlnNvDz2rIyV
z85RhllKHXeL3+qdiWgElhwc3Gxss4ztUgundjO9wwVhVzuRBJb/ksK09akhaouMiT85QsDn+gC8
CNm5wuQDgN/phwZLVx7GsTjHI3HOZJvbHXLZo/ZcsAo+E8OaNiJt0AQF3D2xiH25He0m/8/o1ne6
Z1W/x26heQlch/oin0tyMLZd9Om+pC0k7w/evdREE2Qdqw4AZlf39WM0ehCrb7rpKd269PZHH664
ALeciuKiJURQRZXCoSho5ehqEfWVcLoCD//gLgcSP/ZTXhwcbPCVJNolH2TuheXuLUOM4IXRmYcA
E+PefPBtgvoaNAN0fdO1QsnZa0xsNpPhzZghM8m45K+APTfGQOlBJDCbwGoi/d5D0/MGXUqg9sBy
+7/5UwAaFiWKicyLPQAeF6pQqiUVMxtm1A78exklrak6qZ1XIvAF5UnCt4s7MB04MY05NzP+H0qB
mwihKAdy8L1ke/H7r+FypJrxzqOs5ETl6m79bVCdtHYgQkMRJW4I9seRdmrr3OCvjpdTS688sGqg
VssCr5JxMP4/ay6K8+kudHOJRqZd1EEMSiMBw76Zee7zh+UKNO8tO6MqpO9shg6BPmGg7ZfwkiSZ
a03DRVJnBTqDaOE89moRMF4nsRed7E6PvCeaQb7fn4LK6BPBGv06J3lI+gSYk+aZ8IdmM9huFgHx
HxiJDZVHFxjHQkhp4snIzRDOhwywx1x2a7r/+KY77CWSnTiazzeFe010Wkk0QSwZrQKumbnqpIiq
fRA5Ti2Ruf1vT51irpUiOXgIHRW3D6dq/MNzB64RF1EIm9086M1DT8V5nqW5CKfRAHP7qIaefkVx
YY2hkVumm2VroB2oV3Z/vKLncRzrhijQwPAPUnvp0Z/0SkSFbLPnjW1RxKpGRzs/HxFi+Kh/1zRP
639CtViRduN3F98su4rRun/qg6QCPjZM2IGydECT8KzVG7anGA7IAm/gxlqQo5WWJsWt5lm7XIU0
Koz8Pq/wkeVcdoqst7ptRENLebbjQ2dX9n+HUyfVBh4uFPjJaE9MQxjMG6G6fxwHzPYK4ZBxfKBX
02JTpB3i963ACSgEzr5NcpR+NrF6SkgWx4ST/xoKwVu4jfHpAx8PxLp7p0gJG3fsoB2ohk303Nv6
n052FhfVTzUcapsF/wLo5saRXQyJIZ7epWs8xleDpatbWe1D266aq8rq6UuJX4NBeUJRW93MNtDU
47ZaGOonljnRTiJP8oBnjVEUKOpIlvZcChKBiHLDLNzUtqEEv9ZAIlRs1vku8YYES3MxPDW23yrv
wNCyZ9xeIAT93CwGCLq5NcNNDv5bcdGok8kFS7v2QjF0ZrJnlpzltRs7rhudUjPikTC2Spefzf/M
ELdYRULm7GJZQdwf7dzzSIKgdWZKYpfxUBr2JgZOwuZdJLGz1vaFwRDCRC2hNtm8EIh3JdZ+jBIk
lg1ZXUK5KS8GwcjBJKb0mO2dciVaFDn6xoB0rgxFd3Nit1PNSC2C6GDGMBywsgUa3EEPRhzuVjq0
1gHzvQXxby386AMzblBZL+0hPUT+4kg8TJs7DVlfxAvLMvw2PynnPdQ2rQzxapXL46lUhLSElch2
mBurfN5LVY2AfpHo+gcPsCUR/b28h6F5jU54HZxC/zZ9Ai+dMYA/HF4NaGMqdkppsocNDKsw35K+
DTBGn9jio+RK0W/OZ2hvtWIzZuJqzLrvwwUk65zGYNI9tUPG6xu+nyio6Npg9BfaVPwKDvQ3eAW4
VOEiMXDGxR5yOmZz9X4zz1GQls6fHI2HbVW4DZqhQExDQ+1/HXSoskAQKMu5/MZ/NA1vTBLbPaAd
73hTS+hsAQcpZWmN+apase/bKbGSTIryaiKnHnTmBaCOMoyHMAq2M8GQoTM7kLrVjymLLmWz2M6k
STq+2frF5TUBMrzAeyfQzkdd+AkyFAOJB1oTrhZihykKFGoNh0EVmeCn96u2NQc20G/ROuwZc+TQ
KAmHkkQHrJ+vgkEQlyKbs9m9N8stiiGRXJCVfi8T+uA4/IuMxxyj7u0PnGKa1IMcWen6RmTVM7RJ
hQVtHr5ujCv/4GchiuBMkVPYAlTkCtEK9pzQyz+N+6xIyFQEkAHqE1MbZkEDkQO4c4rYVXp682Wv
fxrWG2mhDFeqMpbefvIt9L5pIemGav276wlP/ZxgpZJ24LLPqrtJ/I/MjbJGZwU0kqfxN7VuEveB
OipeeWvu/0x+D/NPzn1TjKt+2QZWVgmx8SX6QDxdQcGHW2SxWhOMJiQg87s5g9UR7FANifvTpXQS
d2Og123SVztlYJQbbQ1DJ9ab0f9d6EoJFlPz+7rgvBzNjPIygC/UkPkp8oBdWhd4ku7osJbiaKuJ
+uSAeHWekjwAzdKBX2Z78bL2JwZkYz7JitW22c6v0NpE9IGO37AwI2FJT/wZ/Pb+RpIULKfK300D
eF5pEkLNp2wVOowBXwZYbveWQA5YliOLej4VF/yYweXcKtFfu83r0e3CUVIdoVK7eLBrLnuZa6CT
sd0f89/s0YvypWsJPzUQDQ0yuxobqLhhezKGj1nZcTDKwdAVplgVhH8Q/p5enty3Udj3ZmY0W/D8
gI9Bp1uMf11sXu3Jor1uyqLU2AnI6YVC4ipH5mW3lCJaRiBqhdWaSpjTkpMoKH5R0foVEXjfNQ6X
IogxVOLAmF79SHJFr0Fs+Atm1R15Pmq5Qf+qDWQQrsdgX8DxWmt4GZx67emRcXD31A8RONLXpWE2
36Vd4wUaf4r2SIumPHxLNkE9pElaB635OOFCeixmx8JOH2aYqMRNQslcLUET6Vb6C6VabdzL08By
nfNiT2F6vBdLWeA99O+vw1qp7Ive18EXPz5t87xq2lC5GeZTFiSDOHjwGYMazqBOD1tF6XnpwOym
CAw47RHLYdsHpH5N5hTEK7R+/3GxYxIi+vHrFtNJeG9ysXl74MKir6GqOz1awS0FBMGT7yJEvfdp
7EgOcrl24+eXcYPsbQ1yo01IS2NrytnzCoerA8BDZdF5YCPMFYfVrSyTL/kETugJEBYVfHt7sKn+
Fo/Bz6EyveC8BViqusYrZ7CkeRtD24v8b6p65rG+WaHISVWTChNMLR/KXC+qX5w9LpawygnPc5jZ
isGU+JNb0XUab66EpQmfK01YsJVyE9uuUiTu1Wnc3MUi3Dp48z53xaNr+Z8AB6ZTVdb3nx+abJQC
uCnsYCv0j22P9JTbxK9zRk9mR231XzT3MU5+4GDRcdv3kwNjxZV2UAMntjfHT5v9DuDeQL5qbNXO
E6q9EI1XF66LhDshdRiW4PrI2nmsaWqLEiLg7EOe2H2LkXsh3G/dFnS/UwH78E7yYX66Jp6R/26N
LpaXhuymNYdqC4tAzbTGZ4Xrpd0NMWCW1M+QN58c5dXSBGSDTQGUyBZTHsJZ2U2xeWDbOI+Z8Mq/
i79U9rYXMBmz2LOD1/7M0NgawAaJ/z1CG9l0BoBnYvEFgHzQThyLsAMrFYYPCKFtwrnApmegx1N2
zQOOkEkDhgD7K7Edbl2Zqmrf9cGpo020aZHG8RnS66gmclqSp2MXaxwdX3XVIxUS9CZ1aAMbTBx5
+9/bcpkFKUwah8g+BH67qfSAIrk4L9tXUgdniHpv1VvP35gxMfA7KC3CJAeOvJmCPCrTuq5t4BqT
pFu1hnMheprXXfR7SQYaIyQEvoO5r5hs/XvdRV32vI/BbsexxfxGO3a6/1aZX4qcGUGZ3cqq6uzK
SF46Gp+kVd/3BPp4enQCeuaIlij3qySCrDR1j1vEaG+wecpa58P+LsVL0GFUc3wleePvJQJGbcd/
ihT3A2yLOh7sc+NdZWUtqNZ6FYGtpeCURD16SdvFX+B5ndYRXeR5LN1MBnEiGgIHFth2n0P3yYeX
0qVL5d1/oHu6dHCvh9otNfw3c/ZWVSior+ci5LFY+KVvB39DLjo0OD74fSzL7FLmx0StuDFe/xRJ
iK2Dy2EGbtGTY1UIkhjP9PZASmtYUkBL6vYS7qW6uE7nQhZrFfbPlzdOZ1P5lRKmsvlBmsJUSByA
PX0NZL65ENS+vHa04v1+yU+hamG4vb/ApsW4OzKpE3qP678gleqV86XAV1gHI8Me7yzT9eWyk9/K
HblE4NLgiWB3Hr19lHV4k1giDhahoWu/IOOS4aoiCa2d2IyuGHQ3v0owyX12kl/EHtnRxSw7gjQ0
ZX5aUGZsPLt66zIYhn86uUv+o0j5NW4Mmd7jwHNBG4VEG0u7t4nzqCUZ7xOve24BA9AeMAMfCMax
1iHZBzYFikSJ9pKgHJvZCDdj7IwucHlMVY1Ryg9mwFMgRCJubeb7hmGM02/MWmJi6B5twzSu7a+4
4uWs8XVgBFHbpXl/voyXKUje2XR8nlK/b1dZbMoq8m2fLCIUhMbLH4KK+kJPrRNgnhHS++i79xm5
Wbgz0Y7KulUAJ9fRJPb8lxZmb3/NSuSrLNXao+EMGBObXILE0IbQZbaScZ8hlMVrqg6KdkxyvbRr
XfODCEjb1jaC/Gz3PC8UBZfPxRSn61iazNXOuTRQ9ONTWaNrjTE66VI7jpgIDqgueWaNwHkf8KeL
FfzxfRm37jgRDCCgwO4SlpCt26IHvq6XpaegydckrkGkpLvSFBGNx+vpDbPP9lPrE46an9JFAoE9
SHS/GBv0K9+MEF7oNV9+kzJHPludPMnxwmyOSWR9NXHddj78lPoKgRln9/lOxZjUXOEyw+Z9dAQb
Bu7YJBrvj6U2aezJR94jXyr2G3VjtC41CJ8YZYGO4potpSUz5TBLTs+aYMMtSU5wcmkwwAH/TW/L
yiXKYM6Kity1B2Bvp/4ZXXBFZxqsARq2nyza77cXi+6DZrxw3FRwG8oE8RkikomqAql6VExFkGb5
3yzjZ7ngoaAO2lgz2qFhVFnFSpq/8qiRzAmo8V7BakpiTBo9ubFCe5PTWza6IQyte8Da8jV+VWi7
CVIOoz8KdiwRkwMw+OuGrBhuC0BVk8c9bp6Rctapm7cAd1JO2qxFtI3UA+3k2WzauH1aCkGb2Eqa
TrRgjeyIMiYs0ZzhWyraO8+2JmDamHVyTC8MdtyB5J7GS/ypONYtZu4QAeA8dDsGtftP+jceZIH6
/AOjDjnSqZ7/N8qNhTnzJuavXExCAjkqrzrEX7k1LmNR5kCsfYcY6F1VcGo3yE1SfCsHs3VkUSXo
hH61puqi14C0JleAmc7z194Pt4+v1zgWjgikm1XCgA8AjChmrlMYMP0ppVGHzCIDZJfm9WWMBtYs
iz9KEUnGMRHGsok5EyzFx8MgZipePHHpFCQAoKC6YSl5QMYux7HAFlAGBaR2fTBGwH0O4XOh5ruH
sNjMDmSpb8B9QCQGlxvwik3W+0pfhTl5y3heRqZ7dwnLGiX7+jh7AC5VEJBSrOzr+5qGyeuIZCnh
2PaIYaIfqeSr9Rl2/4abF7swvkG+mq/8zPxs6xvIsoa+lAOJ2BBV2YYVuEFKUKc5q+kygrAEYLHa
ZuKy6Ba9SYiR/xv4GRL7iSFruOXH29NaYWQgFl2WOpuUNEhpGaASgyhKVbK4bC7Z48Uw4V2MCQ7B
5u5i473yvMFgc71PN38JdyzHMaR1wjS2230kyHydDw9lCpUAZ+4GksIaMPfen0MzpaqjRO0hdmRs
fIWuqWrlZnOHFmO3kg4/MqSmhTuVsfsWOxdba7VFtTDwGt6tMfUFzbBo90qoCoUeq/FrfngM1e9A
h+7zh14PNDifkSZlAW5JE48MVmAe3QhOfeIhi6GqwiEFPE2sqVUjfejacfCBOdwxrxzNJX8daLTt
mA13PwFahYq7zvgRgCPNdKgPFH0+vHPqaXxiMxUFojSEU3iPCW155nmwzVswUjDSpDWa23xQU4d9
7oJrMt5PZ+L43PP83jFdzZD9ACUDRBU49HFmxPwRMrcdQr5jhBamMv67rIGENRGuCqAK79pep10u
gYgXpEwvlBFfRsyFUKphJ6hmN40ea1BVxtlbxBGjnfB0l69UgUGc14B+sZboyOc7ha/WZApYYsOR
mx0/nD3pObgid2deDGtRB1IBHWqDKd4M/HTiWZP7441BFSvVbiB0WsrVzksgokrsW2gmSMtFzGTJ
jEmBCRFIn9DylRuJzIGUPKRqZfp1X9Flojmigpq/nj6F2ZwSOgJg6rEHrLYt8zR4GbkhB9n2cJaJ
aZ6QNVwZZiAejumMmpQX6jy6JEW6HCngGez9myLOQUofAPHNE9uUcjzGhd3ediIh+QyQaZroil2k
0FFjez1kZYTtvWHTmJ0j6kAaTmapzC7i6sDZ+dmiW+DXP7rG3R+BnDl+HI2m8pqBG4xWbYd//q3Z
9vo7Xg5jzjqKKxPJEATAhSQMhaJZZKl7s5y2PqOMs8kcT0QWs0TKh9xZl6z9vsgYYDUPG0OUHxCY
gfQj2LxE1uVmEtPwyqknyD90f5AmFsNvUFBTjEe9vId91w0f2vvHGfdNnyMDGKuIvtEzQ+PtrkVm
vQaSINW5VlGDKJqHkyraff5r/Q3tVY0oDKjOl+tV4ZzsUoBum2dAFbGulNcHHxD1R8qlxOWn1aGn
8PdKg5YOlDpuYiHDvc/wRspHIz46QNV9GL0us1S8wtukAXIkkez8BRhHTm6BXKv45W+SAB0HtVDm
tBApZRaefGumoIbCMxN0rTp+Cl8kxqHWDPukjGBnYVVJ0XRNLVIfQUgL4WSK8ekYZ+jQdIWLcQlN
j+0woLx2GqmhyQ/M6RCSVtcGUSNdxRg5n8JaWMXX4mZJ3A8NV5PAl/+coEYnJy7E9BJV5uHN2Ig+
z3XgiPH4iaAbhU+zSr86thuo3Ohj4+wutEXpJof11RZ3sWCPyYtHNj0VxWKm+MOUw/jYJsykA0UE
v2fxOtsNt4SxX1T8kLo43pNuknDRrFO3b4JZr1Q5Uv193m7i4yLih5tqvkSy7VE6mve7ST0wIKWl
hKNVl0/zbjdSrNYwP9rLdVoQ7taaTbcLAuy8aVXZk+ZSd1/eWgoT+Vv3Lzdoyd6btZsMU1l3dGtK
DaPcePsooWyXdN8dnaSQJoEXWQTv1/sy+hsbUE0ED6VlZfx0AbTB9HG2eEn5DF7EJVauco0Rnod4
JXhnBZpvvZObf/Ma6Ikry9xMnfs3rT038ORYRwxh13xYS+doDmAdcd0yho1a6uDmrckVSxay3eYR
V3AGie5XoX/1SZBgHanZUZhJa8QA8ztZ2Y+SZttDXMgqMI+GRqdvBf+6IsqV5sP5gwuP5Dn+YFxE
u8uVSqTH4oW/Sz3cyfcRBaAXVB3D7+fIjPpfa7oCrIxuZuwQqqgCtHJgQ8ZCMbJ3DrOn8Yk5Jk/Z
1jjZ/iDw1pVIhKOoHyFcUBwmLI0Y6byULQWIaUsZ6m6MdSSP+GZoiOj2aurxVdvzDuNUZi3x1qER
8EMsYDOKCebs90ZUAjZRaOQ6ydmCTvDTNNaqYqyMmSAEH0tavDkcoGeZ61QIt4mLwsquoikAV22g
JMzufNZ66lpp/K4qQQNhDnmcbtGQtULZgSgl3LcWm2AdNl88ppTlbU0A2F5mANdQhEpBzqlStiSu
Q0bK+jowsv6LLe1+SYj+CXOoMzosRU3ffwPNFd9twCzGIlvRDbUhLNH6A1YcbfXB8pXq0x5iXIzR
RrZgjQiOYV8PH0yU1KcgkcQEnhZcNzi3IUXZw+vF+bs1d3nipFUD+2VGKf8SJAftNvltlaO4IGJG
TlOOCgz5UF56FBFNWzEWJDbmchLVvxesLdY3ey20qTetz5WLMSGaBjPsNHn0B44CBJ8SHg4nYZRN
9C2RwfBfqBzr0NpGjf7GuYe8JyzX9x8kKnzga7ExmftzEmgtuGABh6e+m38StnWkBmH5dkgP07PF
MsKtqYVv2AllynIh5+zx7dIMjnHmHHjs6ROAyAo28AbeDvRGTP7JuIclAMjHFDvUDW14tCv4XS0D
vGSH+6MlQ73CuSnh+zWafz3lc5Z4bb2gIuTMsz1vv5ysLKAcj3LhlCxHYYkObxyIPyPefMcpIdin
7horsjonQZKDwaueBbUyyGMalFBCkQDi54r/6ij2iY3APkA9Wc353/CR5Rag6W9zKaIF6dDuWWqL
MvrByPgTPuKkMlGA2o9//M72Ezk6xxey0HsROdlxeZ3ENZ7jhu7wP4dlbJsV2/sz9eUhVs6B3cmh
GMQT3ZdlyIPVVHRIx3Z2WCTFOr+YwxOy0Jb2h3u5W/BzpmyS6p2sV6wtBFwmFfkoXYHaxHKXdGm7
72b6VbFe+7nnuWJTf7hs4wn/9sPdYU8RPGXAFn5mbG/W/m/9f0yLJjSLo+4W8YjhEMUb+BRC+3Od
diEMBYfUxDPm7/DVc66L4t4TQP6udY483Gg12QvRiFiwA/du3dKxeOfGZ/QQU9lCl3m6S1AE336V
QjcpPx5tjuY5zOAcekYEIZAh8+P8xshclGWfZBMoxLytawVvFcr7Z6hIqXZFVutJkcNTPsveVYwU
56yeFnpCXEwwg61RNboEoD48QejgmaIfj/mDgVmNrn+lWyJfDiUT96b6gQvpgO3xNCnCxeVIlPH/
MDqBrAujs7Qc1nO1FE78cGckXwcS7F8ysn2e+G/zf1cnQE4GfAT3KkZRMxoUZHWB6NfKH3xDCQ9i
u+aLY5ktZ4sGADxeygMRxUzVfbM5cycEM8VY9FifoyXTPQm14tMOrpHTETIsG8OEObZGoKTiBvUC
HAbyladRjnTjSNMX1Fql4mZ4gtkQBQ9Z73JmAV2q36PnFx9Gp+hZ6jKCwTxZVSRYdbkTIOzM68CM
mw/IcIRk2yu5N7dnWlOywFN5I/5QP9n3ZyZA9IhfL9wiLk7fLiLX2BWJWLz+3SeGjJdjyYoHT6p1
0xKqEGhap5ff76Sm5Rz/di/fFISdHqBBw6vdqGMV01aJq85M1NoPjmR6RokCIJXyWo3CEQPjaYV7
fpXzP6tf46ND4HmdKwbX8ilMkRS6oyQ02LdpZc9MwXUfpq/367/31Ov0XWIJMxfo9MafrZztA8Jd
CQZyP8b8BRAmQNJRNN8MOvwjfyV0c7hG2BytniKEWsf3Sbr2SPr2xFkTJDN3jsA2W6EiIC3soRA7
hodJ4Ptrwls1Bsucs+DlHpwKbbB34Zpc8kRQkLkEtAd67VoHQ/95gRfXMh3n3/4aOurVeAJ5MFJ/
4r9HpvR+OT+Xa66dS9ZGUH4MSLxh6LnNDhumOnRdv3FQUHBcVt5hOA9IIlhFbTg8kCX4N7H52fGD
OLrPKyGFiSBk14obWOTZnCPf9I4knDgC678K+z5GcXc9M/Nmkzt7E6e8jdSGjAEUTxkOKcFeMHBr
Fb7VzByO7vTVod97nmXURSlgHpitSlAWb/vmqziLFx6h5wdKyukpPTcwVKO6bUmrnXcVI13FENDf
nu6SRT0SD1uL1rrsBNDxCYU6yex40uMONo+83YWNa7JbxsZMni4kxR6e6s5zXeQENogreYcjDBhr
h+ZnaCI0VsK0KLtcLdqj/1V6VcGtl+JGRfvcdK1GuTRVrHhEHMLo8cO9D6HHnLWoGaLudq5wC7Od
Qhgt/f574r1zBnDvwgMru2/C76zmSWD4F5fHMiCvvrpmh+JNVC3jdUzk2e3MDrPhjrpJJMiR1AgZ
nGlwELOeStWlRI1JurCEnW8du5zFjV+tdXL0+S0ey6vT+zdYH0Rjm35zUVhrJVMjOhmdPlSwks7h
+2eSJZFvpZa26GFPdgmsjLeBnhPebOdL8x8VJUvJgSSsICtHCoFgv60A6Rt6UFC0QOKmf02TIvnb
NGZ2lVUKVZgo6DZwk0eYda1WvBRe1jvuv3/QYyi6Mn1mRZLyfcvw4sRA94Uw1G6Alo8AyNoNMT/P
2+QxWdAPS1nyE4Onk4K/QB9LYmh++jY9fKKUe5V0lh6VAsmlCll4vIU5QyLwhiwI7DrOBcQ9NBHB
as3Nrd7SGbL7/qr6bEJ5hYR+wCMdjx8FMdp4q1hhVu8i//dhebhRvD5OMD0RcaKpyh+up3Ak4Tnd
J9kJ+YqucSOv5DYUwJ+543ezqzv/vCDC+APAiyJPot/zsIIjZ6L04gTERP3r8ifA75c/T5vspArX
MH4qZaao8VuX68PaK7EwgZmqNE+Nm/lvMFXHlt3OKJhHkaekxbWqxhBHlYLtFy39h6K19/qXP3jd
OhUGOz/kItIY4101w5B8gByOY46eJ9gmHcpSUjgE+Z2c8u5/ESmnJN7E4QhwNUgezIqRCCwAsur/
39HqkxqPcqqqItvcly5zW52j/2nHhBWWrMQjm4mWzTZps+DGcOh0JxNb/zaCjdZj1WgjkoylJr4E
JBdwsUnaiuCb4PMhSDqwRpm+LrdLxGJoxtgsNPPfX41Ycu1EPfxn2rBjegX4e7/4d/hRMADGoDOn
dTCx/pXVRM415lDXpuBHeGWdPADMXNe2KzkrhwtJCXCOVyoelHWNfevfeUfx97GnisEgeHvGC5SO
6Gs72OLDUQG6pL7BAvKSMhTFMzuIUAGifwGnZiCoZ1cTTs0v9r9wAoqMu0musVKqnyjmVVEuhhxn
PzlMqScq/e6pczFRsGdCIRIw1Feunpje0TBP7W/FgLl8BbjtvF1BL93e1TD10gXDPzSO8+2EJhaz
BUW/1hdJj58Vwf3gf0rA6WySAvyKANAv74lV9XAJhZHtEcKKi5MMVN3EsDojJG9kZDmAcXlVZO09
hAlo7WAdpKlLrP041Iq4XE8RibbzgJVXixvXfdI/oPduOqZbuBltsORBtUvCP5OF9YJBNbHZTvZ6
3wMQ/rzTkeyUZbJ9haOE889h2KwrTRFWKt1244dGtKZ2ThTwbAGETx9ttMuRSn1pokS/ZwbcqF5b
cQ2egYFZ/5sUnJE3jubBJQ85WImZT0VrxQyhCW6CMARpAmvRBcP/56XNqQYSt9ygeFOVlzlYdJ3a
0HasCOmDh84mvv7/pLm7FqrNhn2EO07/Fbv3JZnFXLTgrliFievrWFDHvv6D0vuhOMX6hgukVZWb
j0cTNgk0BeIWTODwBMDBvJjNjeh7MKzlKH/ITRiyOv6TjBQDc5myjoeaQCqbTdkGNKbKaHisqII8
kRS/kBdZ+wWjz8kOGpQpFe8eoS2L6ILfj0NtdAJTYX286VWRUKdt/Pb1wSDiExXSt9iCKw5t7qmJ
To7pL9L0GnwaLW16MNLFctkzNa6Im0bwYBkF9oU15Iwt7UJ5Zkp5zR436HKznjKBkbc/v0TySW6+
zDgveJFZARsb7rdp3iXNP4hWgYz69aTmEvElHr2E6FbQtYEpPIC/g17vXP1WEFbsAxlx9HKSgWO1
ROjpl0QmmvNIFHbU+cNslAZMObvpLP7H+4EjodLX50isXF1hLu25ZY/ZohTWrUyro1U2ZADsYxce
pLWKb95v56cB2aCgZ8lskuEaPGNelRMWHyaKUZmst+GZQqGzj0LYFGv5Y8DU/C5UmSIQ3aYZaqvc
1gqIu2CjPrdoa7hy24oObvPcpwMzpvgVzXZYZyiCM9HLGfoJkG+10tWU71b1ZyvObU8uemVmtTVO
qfL0P0qr1IG29b+123eXAJPI3hHC+glRBxUv+/Yf3p7fq1dLE+BW9QJS4WTzdgGJ465wa96fBLfj
ePYDk4pRTIpiMS0tfBSjpslIPpTNfBeNPWsLrO3PGEDhmNZjfCiy7HcCu7VV1E3EwGlUFEZlEatg
lCdSPGCd9seKBxUULf5OvManZEEL5Sg/PjJ0EA9dXVBUrHNVlszd7uCEG9k5vQn6ekFN4S02lco8
8nEaXjD+4qvAJXlXNqGia4SFMndp96oqs740ZdkjBZaJkCiNXH8ud/AvY/46zrcwWMMSVq5m+aS5
zpYmEHlpoLNvG5SiA30d9FenjhY6C5shyuLA5REhEDIUgq6E2Ak+gmbPlCKQ4WpAb745A1OQHkb4
wglm7tMfhry9fW4NUS70GBdMGlE3+YwFkEdhD1Ir2PnJy57RWkieQ4GlCaMUSrn+2TNKT28sXmfi
IEEVLxyDynIwairud6+KoDL+QRdBrIclnB2Oc8fvsO4sDAmoLYrTxUgsSGZ+pp01DzTBBZPl7xuy
HLpkgijlIAwvo3rC9j6H1cir/NyWuRd7Oo+aIZCfVoKOm3szCK3GDbBhgqR/ZD6hHmn/67krYy8E
dySEueRriZyiFoFiLZQAjOveozOBrCjyHhVOYu322NkOVxKGXQ0gG8in+KOzgpHvRG/sN3S3RQ7V
VCtaKEd6BH2PRBDjB1z8JaX16f6scrfJQ/xrPcK4nUv1R/jMtKooLvVO0anBw+plIG6udIcDQKRQ
5Q33qjvb0nIxa7AQ7TFyjqbWu4yvmXByqgmAGy/E1B2SRULmennc18GNznxEwkhti+NIe2LvFIM4
9syEQ8kd/Wuyz6itUxc3fA32lr14Uae8DXBdZhu8DUC7OZrLk+wVDJa2wzw9QOU+zFlGRW5+yoj6
vhsIXrdXUGJaw2ZBDPU0VQh0WU01N5As9IOOr7ODPMoQzA3K0H9aECkVFZmia9u7scYiU005JuQ6
1AvXb/Hw/nIPUW0D79Qm1ZoL8I27eN3tc6HqPmd/xjla5DHK7YGnA9LSKGBhxtYgVvWNaheFVFdv
ax4dZORs5Pfkl/gCVgZaI0MyKT1Nr1f1V4oEfgtMT3o0jh3dtucc+GCpg1wI7Up4NR1o2sRHtcxL
zssCZ7DGIG4PMQxiV2T0oxiAO17FKaBI8BM1OAWIknAsNhfOTcrk48FcObEAirov2TCmgq5xog+W
o4ht6vyRL0s9IkEs1N1euZ8x8g/Rql2hwWQErRL9w0pGSzRngWBC2OMwP1vvLOtWSHO0oUsQsirT
Ymqfa31RvPLsUR22rwzDQWMsAzbV9plyZjlsYyzECKcRVBaK5Ehju8W3ktAproWprbbLX4aD94oq
mie+3WUrr1j8kmicLstzLO5Rt3yi6hmFs5KFEQcq/TNdy4L7HmuRDLUN4/lnez8Bx70ZbzK96Q/O
XVWWtUhCw+Khz6r9Y8vfQHn6H4loZR+Xvu2RJRYdBOhRKCqIBUUzLdM+ILcG+XvHjYGNq67bRfvD
00Tmc/jqH/Cu+eIZcn4VuIC1SJuT6Ys0Pgb3icg5J7qbwK+0PN6o9SCKWkJpGg+93JBU+kDrj+8H
ukAqVbxZ47aqkuLPa0g14z6c17XJd5XvIzfhIlcL5TD+HDt3aREoAUhfsi8B0eNCQuVRHctkruI1
fIDYH9cJzhQz19jM5EeI0qWWerr9Y6uQF+7Tz0qGIKxQ+t7KZO+5DQ6jo4Fkxs7VeXfNpitLSCjT
GJP/J8FDVbQGn/MATu3izuemIs/y3dpACgMBiZYk1xFlLEB+RupQhCKSuQthqVIDNFzxlo4v+idZ
Tnrt4NZfbThvPxqcjcNJMWhWZNZbrA4rc/8X/zoir7LuV9Uim3BHc0nCBtZlaxjnsT9ZzbEJiiSj
G6FQ/rwI1Ctyx/8l4RgqT2rJKUhur//myI75O5u1moMNx8G9GofCaQW0NqBY80WbLZ2agjC+ZpXm
WIOs1EisP/EespbOP5AbYVsl7gXCIKFa/8lPcAUp5aZguxxPILeY1N7iUVrYPjEcRBmt7L8q0h2R
LZzlksGlZyp94QuIuNwgqB+Odi0jh7g6jGAEP+yAj7hF37J8UTpSABxcI0tYp/wkS3z61ks6m4/M
VZhRFLnysXcCPZe0bA6GeD+cWHqrYjAuNTYGIbiqMucM2BWFHIMLcthaG20jDwdqE1SjP0xzOml6
S7BE5SgnEjr0L1iZS/zBWNxAfJ5INSWnceg9T6hGkZBHxY+cQUYU8FintNbQIgNdkqIq4Gf6skSa
8/W8PC0Yaey64WGUqPV7woCTKUdlJKBoroJQ2aw7vrs+aP0MK8EIuVwgVEaXXSIJpnDwiY1N7YbA
L0+g5TYX8ioQZeqOt5YTU/9eel6h0IeIl23jdtyrWaSSWxuszYfxR1ScOE5XC+s1+wm5XefMs1nv
pXewp6qJEiHfHDDxPpCSeYocp0JiXwhOTmljpCIlDuLA30+WM/R7o2bgoi1m94FtBp8AXE2PLYWS
aOgmhtRogAdNaT+c8zpzJwXRoMiYtvUxjg4/Zx2dbvckYyDarSCk2jKA3X+iqRcaqOez8OwDX17M
RaNYtKMvTkZWrwg0nBhADSAsdp5mqWeTuQRlF6sqxpK5Z0EYcwsWVWEz8zhGEW3ovb8UCudloDPQ
z526nohyG529NQx/yRMAiATug9llc3rrppOAOqTdAFwW0s8vNUuj2/qYcUuphOcPyOKAEDoGo2UL
AScG/3mJ2wG3nEjDpP/gE/YPME7an4dTlnilJ1oBjFUeX/5WxNDn1gjrTADkUvN3v4lN1aS2xyjM
pzzSUXON9xoCeYOuxc49xL/hLSbUZ4rzD7NfRLVl86OWkVH/ELcO4BV+rrRiIPs0mLmSDpC3cSLp
XjcYINBhG9E7EOEl67S4t1MQUDeRLUBE0+L7CM6R/qSV4oSy9EgdxTy9iY0L2LX8vQp5aNnM+WMF
MNncBq739nRYNhRisYfqVBW/+tYnNs4a2u7LSQz56OXa2QMLgsg5LEgwS2F+EAMWrjpEc0zCkYnx
uKwDIbJ8/n4R9ltZviYBn22nZA7bTPV16anmq0lOwbJtUrvHn9of+lY4MNNwg4xjt/0qoBeHXthj
uOLkuw/V6xr0LYI8AMreqypyrrlRDNrDaKQ1JQ+puYLtSA+Nq1u5/o8cK4r4IOyRXRh34+ZQvnSO
TLQ3tfRKfWv9HfTeZIqdk7tH4dCEOXGZmfvCCsDUY77lyRo/4VX0JYRzh72KMu6EQDNnSN8f4aQw
qw53DDsvGA23waGSmxiqzsy19AzMocGFzic564fg54oKP/QOx9XxAvvdebvXM4RFRaCxuGU1SM9d
azw7pJRRDaOR99gKpC3A1OpxFDljwKdi2FTy33jAIiybegUHnjd+71JWGhEyv0fx4XWVUdYqp8o4
7s5V8AQca/4JR1+0rqOmjC4JexxssVVRmBeWJ58F0JfqtoGnlNX4lxvs+Z3joYc/MUoiWCsAm3CY
Ymih6ukE+jr6IwUFEwj3R3VPtEaYFE9uxAmLMpu3xY7xpROCSfKLDuP2V1LCgORln6VM0aeXHTN3
MmNohx0YlHvU8MwxiEb2fFEyQm9BruyGzIUBgPlPEJ2Lkt24b6ZIx+qD3KTRDWqTJd5DKHFzfF+M
8s9XeGeVtsZLuSSmz4Vqyl2j5iM39+0xsTxGf6zeZ8VcvkA/Ss03ABEa4Mcotp4EPsNAioUeI4Cb
EBJ5ygbuYUB4yqfFa7PzOU6hG1QTOixuZH/VE1KMKkgoPWs6Hgt9WTxeHZDvtP+3T9AR6nJRGslt
T+98hhColpTC1R0yDzp8GNT7lPKiw4o+Vv4BrDkMAKRxFBdAV3oOQXjaPXHE7FznP9dHjubbZ5H5
cB2DfZOrc/MNSM1Ej24d9TAinDmcrEsL+V31QxccStBZmB7ckWSLu7ZKIAXQM7HGJ4R4/ZVDLwsK
+UPx8nt6oshh7WhJ8M6lotXUGKfwYLYcB7XyIVMONe6D1CveW5l9ekwfdSrUMf1JRA1Htmv3baKg
HLzt1aSGnlL5U7hBEPpaGPSoNPwFhLNoT8iMMgrqpoKUDE9VGUl13LY8ew4mut+5/WxMKZ/M4NZY
sBfKDp6enxYMTsKT/rKNUd/LKW1SmtB7nMUmMUA8PGGS2wKZux+1cgiHLYua77iEqpZCxGxrKZ3C
3TXavAP6GGsVyS0cb7YOxXMBlgXHVhvMaCw37CwnJhMMBdnZ3C+WhVdPGfwU9VqMQd5v9zLbIyAS
yFxukZ3Ir4FkWAK6S1+X2AlZdMmN5XSFfmslOGy3kpMG5TSGZzXO6WUH2myyTi61ZktIKB7RxoDa
niNpLAab2V8Sdm0t1d+Mxj4udl/h02Z/r/9+yrm42WABcjxuvbCoHHqMTteJFohKTNYx+WGV2kbY
PpN36QBU4vno+mkA0bFvEawv1kvcm0qj0OUwKFh+yklYuu5sM3xsWH2yxdrlNm+QVGlDKZypw0tz
p57bH+j6He+b0SY/jn3BXMSkB5VYsN9njSRIDIH2tofjKHVrxONvKoSpay0LpYK+PZSVnAY4IzuA
BfRbEk/RJYCl2TKbHFyJL6oiz8qj60vZD9AoC/OLHiVGDssdfzVJe9ycchObSpIFguKtKaX1jlXc
7fBohdkoIHhIM/c8q3MBI7pgK8Bd1XAxoru3dJ37gZ/tKzVAQn4TfeVpr14FnVpqul7m2Mr9jiVj
oYcVi6tSJqzQ//B7Q6enlG9OYbTu5lzNx92Rkyv+j8OpPqFqif5T30ksX7OR3SlEQ8eIcVnLDBkK
aTg1oTpqBliwfbj0kIozR1/ItkwHpnTQDddvEashhRk3Ca73tYTFfx1qMXUdx6tsAhsny3XTQlS8
t4Nd/JJI6CgDfo5gumo4Wz+v1TG5I0INpO4waj3nUnhlQs7/sDXa7v7AIFixy/it/yrKkajgev9F
IVrmZyBc8QBStlEdc97ASEvFByc+jhF587r10ooDaogkvDfeHVeildtrql9jqpUFtgZ/asgj+4ON
uqgW/SSMSYYJp3nz+w2cX+mOMFB2dN5d3w9EBaq9V4Kurqcyiir0TKbDG4pkU7sWfny93R8fEyyR
8N/D/mv6g2FQ3CmM1pTmdJ0iuwsSdNovxdeviXI6G1nXHP3UTt2yllXE/1W5VOvUxWrSsQt2m5am
XCHgdpNfY22+7QlvJSnEOa5Wpym7EFU2YVxPvxk8IrpBg2sbiUj7eIXZ8BDOoGKVLFuAbwzOLIP9
doxnwYsUtUD95J4AI3aMMrkWZTTgmaK/uUjtcv6BfyF/VPjkEubuyc5tkB1oQDB9g/JK59qIEZBq
p2SrbBhMlYerQOteD3c/Mb/yV30ZqkQ5OpparOQTqLpRbN8+GmQSxdQWu6fmFTxp8BGnRqMEcJ+e
Tea1uESyaKkmF5kE2cDgBJhy0TCsvzAHp6QoZTodlCEynAja9xaixpfh3fCE71LqXs0JMOyIpOxS
QrGnjltw8EnhRSEc1tK5KPZJDYwaXjRKLcc4BCxPRREJskFSElf2N1MfZlo/g55nRYygtWbnQkpJ
Bzjp3wehHzRM21L78Fs/jCK7146OiAic0A0JTFV7tXjv37NrK+Y7BuOk4bKs4ZP+2JvExGL8Eu1S
hua9pr2ao201fJE7P0wBBv+2fBJRVrleZxhu5AUaGbm3smHgYQAwPGFfQpjtF602Dl1+BAVy5l4O
1zxwYCAi8MVRsLWaxrw+RttEOqVokPG2lCIlvGcte4ZdKHlhQYwzIMxt3mCkph7HyP6yY3ZXhrl9
q22GFhe6MPNS95nY9YzdL7i/cdxPfuAOqAou/wSVGa7Ja5/9dq4JH5lJC8D6oXh90NFYJxWpo78j
M3i7qd5BBaAKSLpvBADY/WJkX++NVBcdrDeqiYG1ZaDA/mKvcPrlJOMFeFYZSu9dZkmCTlDUn+di
EuGJOhGoGIGiyDJjNJ6yXr6RGzBtcpz/EBR4xwugC9Ie2x3CpGrqR3aNXjPQNtqM+igMpDYVRn0h
+A4GR4QtI7xNr3yFLmVb7YwhcRLDkN0yU/J2w/ECnkOGuRXtoeMI7ELixIWO7+/Y57YOjecwH9SL
RNIIWAaoLqLGP6oYSxxCTOYUhnFe1NT/qbuP46XuMzgojQpHQCCdBIsQ5JeaPhMmojjutasgkp7j
MELvyNNF1TntV5GWasNfRfAmmDB2RQpZf/wMBqjHNsVhvCIxXxS0GnbdNfb7v1VA9pEKtJB1m/rK
GjLeDuH5AdlDjqKxsXET/8oDI6TKCGisqExY2kgVDVjYJYjZx/qfAwdgjADFIqR1hqLP4BYUeq9P
dnOoV1FsrdGMeehZ3gUQYNF2DceXLgk+lDilZGgFiUOuWQy82L/AF+V4vbUbZc2E7r8H82E0qn2p
ikVUZGk5YOofPFVGqhGGarCJ3q1KQFPsPtIYSSeuM/GqJLlnTpRneoa7Yz2u6PxKJMgrqRGiXpUx
Owog4wm7RE9vbgWKnaCmuFOmRHH0q6ljJOcIr8/JBUwbzV7wIsaAtNLCPAvP/4fEH654bkGQxbjv
PqYkW/UM+cp9hWUkOnYMTAwckF/8TBhpBv2RlRkCCfCtdErx+CltSWkjZRMfPJS4gM1DZInLOZEa
vHMkl7AtoqxsQ+ryPnuUHsLSqvG9qp5OwfYDozLrmjrqMbg0Wx/VnaoLvPBeMTTd3PFNmfLUbcj2
a8vRg/38sCaTpNIiYwTLrJZ3dQx0iebLRJmSH8rmElMxlp6ARdCZul4ofs0PukLDsbLZDAdMqeNh
3jE12Sot2wF7/RToG9wQ/QQwWSaOBKuDhgK/JaWET/w1BsVqXH1tbYfO4Jctq6iy1mS0fzEI02aR
EX/ZH/rWKecF0hrWdz5EDddX67UzdtQReixO+3Ey6KbebYLBnOU7MbAcHy4X7O1fpV2khlQN7mrL
1W9c+8mYxofJ3c0c30zmhqrU9T2gcC9oJy2IR0cUPhDc8TEb7JAJdy0viS4NUZ9dndDYKF67q360
ADNRk2mCanRHHM+dYo67tDBUUbDX9qbxHYlKEhKSBRO4GK/2hc6kM7evRLMu+7id3NkZwRoiE1+c
aZonoDhKUenbwIqsL/vzxOEWwp+g/sLR/3Id8yLg24TCvqu93VeBzQ9UpZJz1QLVixX+16FVmGs8
aOcjfjvmeMdPFLkdNaYZB1wtwXTxedMwJMUTbKeZqBgu6jg6Yki/l9P+0NK6gO2JXrnxVQhDuf6t
Z2d7C5LvnIlF+gnypzYnv/YxNpes3xRSxEMUPerMSvuE857UCE3KJmGRlPyBGCz5nSY0M5wg+lU3
0pB1UBmbQZ8yPDJKInHNhz+PLJyAgKehhKcMvU0uVEvyTOzvoydVWYS3Y9wGojR/E0nGH8vIlDDi
Nye7nzc9USOAN17Kbxpd1M2TgRoEYBRfPJDP6HQqGRhXlFy8QW76w3nuFyqpvaodMfcio/iXHokq
abzFJ/YALGinn6NDEN1xDTSYcJD2Q5Q1XOmWZosChqQ0VFfp6U1ZdkzFPI8PlRArTcUPFT8Y4HbW
rq51VrDmWzHIUJ7B11KcyQvsAPvLJSBbEg3O4jHOS/ltgHs2kYzKCNYWg3Jn+C80HT3LYRhsycxi
HeZd3PFwsF0vr8sgO6I4myD441cUxAapeA6Kf7nKiY1Dz5JXQmCLW2aoLdNexI/NKy0ECBPbGCAU
1yaGoFYniM0Is6ce/qU6hkelBn8YGe2OB+1CcPjvU9HciA1Xb69k7BPPHnw4Jw4m/UAVPV3bezA0
+WhnQGHoHEot7hShQ0UjBHdPaEcBP3CJCKkG/d7PgZfOi5Qu4lXCNXm9k5rHs/+lNBvzJQEb1Qpa
SfyTV7OexWFgIt8HEcTLkg/YQxs9HK67ibuYGfuVgPOq6tfiCmADyepavlbBig0Ms7nRee2cOv43
1VFI2jfi/MkU3Kp98fGMK7Qqb22AqbVE8v+HSLC2VpMrSB9io59VEJRBqyRmBEQJx5kcMmJwEtNc
wEPPcAryw4p36/MmcYnjfkMhLdcGP7l2ypM8yGaFJv2+d4Oby57bohfL5NdvTwlHIzvOQAoKBwD0
eLC8jZek8wn04Y4CuhoM4UkeMgirzmchKRFe/1rHtDzqtofMtyKpRTz/WUHWOotYL+5PKcDBCRb7
NjJduxpZaVJV3TDrLLZi2BYuqQVRfLUirYGlzNnno/6j7hlr5YdylMn244hANmkDzOvgf7L2j6TS
zwrSAyKiWUrKpA/ikmbx/6TUYu+CRhZY7Y5fwWM55Lg0rRRxHWaJK4vL20qAdXp6FEqpCDrg8ke6
OBCsWa0H7bsqeY8ZXv0R2ZJwLfSOO8xwErweqS9kX1xKKnNK+WBeonXyRNr+0CJra4SaJ+3Vub/N
hWLwprLrX4Kut8Jof9x+BD0QfjlOhx0KwpYFZSws9NTmUEhLes7GkNoHrq7gM6FC5BXWVCIr30h3
s4cmWzZwUDxOLGxDMeHUkA6MgcqeJZALGrflbSIvmdgiVoNUJLOB/AwSs5AoJYiLptNJxq4aijop
sKVZZmmuQQadz+SuD9YtVLyava6JDdibX2x8q6ecRdwgUtmrLWsm6bgE3pLIdi6ikHy/fqhpg4GY
z3Ni5xpKmZ56faDbchnX5YjTjp6i/YrohSZ4ww8JEoHQoMu/m/AvizB/mRAhSnwMGZCkadUObwba
itxIuGIYPS8ewpMvgQDTUC433ePcQ9X6+i+5dJw6nIjL/mpI0dN6FK8ElGcz+wfTiKLuoVYsLJtn
WUxfnfCiWACHimwukHguPJydG1nF3PB/SN+1fzQrsrUjT88vFIKRLGwbqUQVnexVx9aIbSOMM1FS
yebiLuEmNkQeWn8tHQKvtzFjOWsvFqV83PWWFZbkS54yjF0Ilcw6SoXyuKo1ZAiHNr8lkeVgw2RU
n9kblVbtE/9TbM/yaL4nCajvNI8YTxCVSCLgaY/5RjLLn+dHZOar2dOeb07YNxQCB1WQ52mQzSOv
O+158Dw2vkzMiPCFC33PWQ2oufiUtFwdFvlNZrIrbSv50AN+RZz+J3fDT3wARLzUBEqSKpvJ7lpn
L1FJEjD/30eo9aKpfvcFretRlORcZAecfWPuW3mws/wMmRZICKQHYOgSXY6xFSzSo0AjqPJ6LhBV
DejZVikoIsa9Gh8ROGsauEWeIHLUglZdR28Ri8QmXGCzpfYG9sHHI1dJXFHUkNETUNP2ISvXsD5s
lIdUq3GZfe9/aqtW3W6GfMCKDAY8UeM9Anu2+YxmHWJ9Z4gGWnFJZt/f+/Uzwwfda5asljtAZcW5
5TW0nEeyC9JS+RBovA+8cplEHakjXs8kRIBR6vfqrTmNV5TMUkPbqfa6zm/7i0+F6/dTyUFZoBoR
cc2INtqF1GRgyCYaokWRihK/iKT92Dunq/sj144dOyVVHeqDtF8NXyGKOAA/q/rFic3LenHnDWzL
VRfdT4kfypeSLNzWHKWy5aIHiTnf8FTQsDNAGvcgtKut5vq5C6OG+543313QqQvaVR+5e3v8ztcV
++AM0IATvPMZG91y743gE81+rzdxINapEsCD9AxE/rSZDXxteL2JFdIL/UzdqcpItCMET8B0QqXX
wtmJSMyM96Esoyynxw+Od0r0ocRWegXpT3Fxylk5vsIGM29JePAJZB+x64sG1yxwvsXtVP0B32Ff
fcVNu5MDUqyrhivhTvXVvIzvmal4JHjaoY4VhPOqqpQNqllO61km25Bd6eNl8+DlEBbphG/0jGw8
JRvHB7ti7l43lMPPVY7VpmouP2xd3IAetMAAntAnfRApTHhijR4GdVryJg3N/J+cZrvjZuATWNqw
mS+EdihKcA30qO3jdnFtQKGLEG2bX6/Yu0w+AjlEY5jG4ybOYeulvNxngWZyiSu21zgStqp7TI9a
TnIc+GXMyGuOnA08Lu9vwv72+TCc5ut93FyOj1ImmNIuK9Wgvq0XdyFb8hxMxbS3YP6vvlf9xLlJ
wCtI4jfk4xZfCVPot2ojroQMZakzZifrciiDaUHlq/lNNNE9uypDTrOwA6xd2BOs/2gz4Bf+MBqw
0U4SBIWdTrwWvHOrZRMgyt8x7s3JN+Hals1fv70Ivc2owCM+VEKON3aft7rkMjjMlXSFROmWQMjf
JgxfYKAaWerWpYqyubd5SFoLxtqZQ2enIjX6GPxaJ+RrIvf3DulS4CD5Sn7JDapPMDui909Ha33e
TQR/uiZKyYbvZ16zFkJ1dox3sqEpv0H0EGaWDhiauV//K/x6yPDFeMODp4iqUb2AxXZJ18ra18Nx
izc8Yv2RTp1C1b/2JABodE+jXzFw7pOaPGqjIfrExcwdBEEyIHkgy1uu2vK24h9ssZZ4l4NYPQrx
nGubcfBEE9f0BVdmbof03H8GkNlAjoE3imaXn9S/i1hGJeYveHSGWHRQzQwPidxE1bXFfVO1dbBB
3t9yYys1mhBy00WMn6yVpNqyDqj7tzQ6utJe/YPAHAvG9PaSzrqkL5UKOWHzXP+e5IR9X6ZdgX4D
WN/TQh9CZ5T0ZlMAgSKTIcSuBVlreXtzP5QsoHfpMrCgV6gpJN8uMHv2CVvIT/3awxsq1nqhnrQS
JynUsekdsMqTXWROY7gZ3Sn4u4T3GmSsi8EmrH/TY9rKKOit5mJhZqwTGVIVLBbEhFXrp/YIVTDO
L9Lb+Swr5bzAFT/j7YJiSY53M6aQmxafPP531u7n1fXh3no9CQGhWCfLdzPO3GntyuNQNSTRsKwR
NRYU7gdt0Ioj5ioYH2DIbVapQBTjCnHv5NDfjA+2HQiWVLAoCfSVjO3f6JQfrGWzSrbJ+XfIu6u0
YQOyRxVnlXuaKjHLycQXJItFa1c16vxj5soWo4YIUloZukCCBMqFyzCGHjDmJeQ1RU6PAyTY3JLk
DUftrHeCVZECDh7jarGLKsGo/6DIcfJWxlHAxJ6iwvzEIr0Kp6DoJ/ZHih7dWGUdNzse6Qa0ILvT
/k0Sf5Nq8oa8TlbL1I52NZUEdxBcwJlITl4EertvjdjcP0V0PFfn+dsoYjggmXAYosshMHFP+1ex
rj4MOzxwJbJhAva0n6Lqm6dzD/5bPuv8Sp7YHMPj5IUGLLmkuF6fkPvwLZU4iL/VMrt0q/gmYQ0E
1O9wdbytnvjNr29HeKaRn3icpKJe+Cdu6nB5HFR1Zm8UmVuJtVeaPaVOTgRWjK2hUkC3rjjPcW9d
A4rlTxVFYTQcnwwI1fV25lfwA1VqaNsKKFsn07umJpI9IzhtrvciggeOITxTbkDR77xWfPRYyADG
PDyTWylRwpQtpfOiOGQv1NHNEOJfEeam2Pg/TGXFcfMFVYRnOR1++nE8JonluW12lhuoZFzQEUww
5dNqDDTYgZL076WkLKUhQJMDuTDbr1DbGNHNA1HdFHLFywitvCJr9mgwxXzKQZZFnd2CzE/YIh2g
7xGS86FB2KQGaorr/r0t+bIiw8X+u/eB5ytlL2S5NyGQX+8fMnbGk5SgULWPcmgKRmM3KVyvaBFi
80u2e0Zp9tUNjyRa917LPkvkdQ3BjaCQai8nBByGBHHy83X+jAc2IaXGF3n9Gs2BWzhAhPOoobjG
yYYioAYLkGvqFe//84eb4d8FgVa9NSyaJnflfa6vLzoElBJK5zz5rWmaHlqWKJESD4dt8PmY64b/
Bsohgu7nj/tnDSJ12rDJo6T9Vg6xu1aMbeCjAwTo4twUiqT6I4wTDoWffxYvu/03HHrCMwshahrM
Al3fsx6L7mfe7V1MmAzUnuoOOyafQ9j04O6KZvkTMNJ9dcteJnMGfFF2xjVQuU/n0p1h3XpDVsoX
oJ0kT+8TjTCu1tjZQh8V5iRcuzoRTikt30QbiAmTqtcAtPnGS2NXn18qU7MXAMvyaXs9xB0cySgK
3k64MhHwqf3S2ko+oCcF9pRFctTISKuUtDVqC3myxz37YfdtMda0FteSAlViIe34k6bp7+aQPaqH
Nw6HVfpVfm6Gi4dW2Lbj/JCIu/xAdu1VVn/MVBbpda3NWSsDgQGjwGUKMd/h4fDU35+nvORlmfcP
1I1tNKK78xJ3uTbuGDguNC9OM8VuExRdAwNweRcOzF0zpiJ1YHn/yP33LlJKV6Fp85635l/1MSKG
QPOv5OVffgxCZcF/cFDrhXGAal4Ibba9FRvSqhmWX2SwLUz/y0d64wd3V2FB0gACtZOWPu1CWs//
L2jtUOjY2LsiwxTlF70ctEnUtRcz8MkZzKgt65j6SnpBHJxHgjaC31KwOLdGlTeSEIuX2lPleuEy
2AcFhkqXfzqRWBmE6kPq3NC0Fk/1OVOB1lklzAPBbRtW8dSkf3FgIeJo0FC1d0BksRVc7x2tcRcZ
IJw4zbC07IAcrZSo0RX+holCbXuEvatqbbgoDesO00HuRmGlEBQP/mp3twUwr0kh8hvrTR++CaKP
dsI4cAwe1uEQJNKPhLVclF3EyRNdV9Vf9kGmc1UYXhUBPuo45QLIIG4m66lHjpNbtY1198QG3jRY
Ug2OJvWzsN8d+S0OwjWHVrtXhJKPrTtvjXfH31L/wrfh5wSSZESwQgJdKLDituxwkcYgCOEQBN4f
ftaYH2irCjj+pDHZAWTEjZKHvqG3ah8spXuhxVMTSaG78VHwWVz2OYBmz3zTJyHgF7wW/jISFs8c
7lx3NREDXJ/usmHp9gYvr1Bd3NBehZhwgxP7mZcnINL4G4OjedcduK+qz92ioVIywHn64q4J6hMm
vIGdITwJ9AeUnyuC1RsJfXz4WoWG7QdZ2xm3eBXY9zSKjYh7kHI/9Iy7sEaVpKwt/vKcPPZNSgYw
Y9hCTcUjJs9ReSsKxWPDLOMmZ0TnZMAhYl5leLng4aVnBijUab6SHHrFMa2xPnpLtmJ3ayzZUiA4
vW67bMN9oDq1CeE32Sles8mgfBQ7jdwXogNV8T0h+14Kj5YtBzauVK6Z7L46j+WT9RKOdWk0NjrZ
rNz8ILXn03Y/KL5OcLyYHyfyWtTwzU/5tIIJMxyJFOogahwceAZP2JTk1kOFTHpLiJiW4kTYTtYZ
HgQfRuuyRNW2uE85wnd74jObriKO+Rx2zv1+uIrFJSzsxvweuLIopZ6i9pfZiecZMD7GgBP0E2LY
blXXYO8zhCZSA0AmYfgSaYb8jv8ht8RLAs0rxWh6t4n0TqP1H7Vr9Q3kJ+Z093ji4jb+K7xV3sWT
tpSEdgY3zg37Q08Cj1f/nqzyNM4nRYtJTHlLD42cCWu1LvAcK+KD5yw43+85a8Y5HnwF3E1/Apiu
b2TGu+5oKQA7aqSUkFAm74ZPF8BMHLHfvOwiIsLtdt8PMb+W7F7YO0uZKUnDSWcw6xKzn9/bQgzK
/Jhp7P+j0xSy7sDz+BaHDg24XWSjyVQmaYnIYiHzuX6nTexFIwRUvFcgDZE+FcuMXsmnmuGa+9o8
7J4SQl2nvXtMyHJTadfhlhUNrNg82od8WteOIu19BdtNoqhhDCBztjaQpgAPDd/ARuZJwhEYvmWg
XFOqTmLl4sWl/4pbkiY3NOodjTvN82uh3tKijRrIlbSB2kTdRb/YgXxbmJfDPKNk1PwOnXyJL+Ri
7/p+DPJ9/JEpBBjdlu1YuykznBMbyg7XXd6rI9lCRp4MXf1AYUIqAv93+ECY0mp2NK1yb27+1KRp
95LabHJJt4M9pI5FSCaPTo3A1H2CKwISS0lAUHHeQEGFmAlhuc6upewb67qevlHzTBlcjKGmwr75
bKINy1F9PYwx1mLqOVcrSoENjE5m3J9qVQwOyjDFEa3NUJF5cCh3rUSVSrUXN1NoD8/xn7NG3MPe
ehcJ2wXPEt+lC82mR+X9DIPHFUAMgCkuC2/40K4xFcBcbozrBcH0yhFFE62iRoFtWQNs1DmcF7Qm
KUD3CuGztQ7Z6YF/iUcJubqhWLDVwrwkRLQVQmN6U9rfzjg32y29k6cx1YINqL2HRR7tQcTQArNt
3O5Nj4ZmIn67KJzHNwGGRA90/6pQtt5gQ9iawd5QF638kZbRKKHqaHtx9njsuDua32m1hQVmI1y1
4WLUs3xKiIwcs7/frnMzc7L7d8xQ3QkuNeZSM31fSX9BBH6CnHfUmK+yA6g938Sj/rtFEYMVxnz8
sXQ7y26vOcvZBoHV7iSXDyVpYF1TObgGCxcqbgodV6e0jrOJqAd5RW+RcEgo/B/nlUC3YsKIbDZa
W8wOUbq6cco3ZeFkYMn8oubb/gaZBMc6Q5nejlc1IGBmOpa6WaBP79BQ4U6gjJyJDngfrOTUoJ0P
UfBUWtyWAIdZpBz2KPr82X3R7VQk6Q90dl7h7mW7N8QjfQv1C5kKBxpFuDDcQIoX61+rDlp6K14T
MEv17P3+ffCtfhVFnmAzYhVhDh+m71o1oUejN4h3FBzEGebI41Di8dLJl2W15iDbOiENE+Vf1HJl
9YquLQKQ4/mU/ZjuDyZjZOLZebNsiQRCw6qmq2eWobWcUbog6GVpBTQ9lJ6lAMEhj8QV+uDs6cac
w1PehZo76T1XfH4P1UVNftjcnPRU5XiXbAOq5db9qBkzNzYpe0psneJJyQPNfrAzp9FjzFJelbtG
4ARNdXmLfCx7IUsAOvedp3bE4Vgr5XMugPDeXk0+qn7z28yaDCJSTuWRqFZfWi/uHaUpmaGRPG/U
DdoqJ5DDCEXWKr+V38R7xubjb5RvZI7Iij/n+N3RhKCesTqzRnDqxd8k7/ppddK18r1BZ+/KJuQe
5+3+jGiGv2FpnQJSajI4KzI3XLbBKF6VrA9bKhte6jJTpBNo+SnFDfG+6zQNr5muaJ6hGQueDPgZ
6T0t7AkmKZULtAM2NR2puueHpcA4lXzJcxU4FFVPKzhclZnaIx7Vs9UpACPL9PYtT7xamXaaKMKt
maNhXc1D6Fx+c/Z1zMVq1sxCzt3M+lPiY2rbubJpP4CAmaoWWl2xsDiwqKrQYlJgPCvMjxiqn3D/
yKYL61rahtX2pacS5oYjyiEZVFSJD6DV0ViRwz2njwvEul113imevo/JOiXiuIPqKGbsLm6L4ja9
T9p15JgvK/2xMFmHsDxmd3taTMZu+QhhB931+B797Nisr/V3+AA9s6t/pXXWqfBSzN6NIAvtizV5
tmvmpGMCSGfXskiWkv+/V2N9sKQtDRfa4cAov83ujjeTNDiOWZrDly15koD377pedmJX3eoOiwho
62IpD9wfKDvJF6tJQ8DxWATg2h5dghmVY9Ujei9iM4l5KoosljSaNpo2PMd36R6LMT65cEUJT6b6
YP8pcU4sfjZc1R1iqiujZx9rfcz/k2WjTE9fud7WgnHe4cX4bPtYp/5OwBlH4+a1CHBS66rlkPDF
Hoz6yeqsbg09eRzp+7XswcpwonF6ddM5snUR20do9ez31olQfA3g8c7xXSEAX2TSPLqcYyJHSOyU
Vz1QQVUqtxpnBC46brnyzCQejQMmOA5E0oTybpP7ALDz7FxuoihiNlbm1AftlfxUCcLZrcPbuaDq
eD/Vb8qONSllW5v7xZh09E5+GQbMIelkFnLUGcAM0NxCwBAnB2CMj6rm9qLSh418djbwt+cV0KI3
Im4nyqROW1g9yS8qvma7WaC9nOwz/zMHR4u6nFk952sR/sj29aHhtiK1ybbZ9QXtha+JxNtu6YTk
F5w72stLhZOlXNetjd3i8znExShl/wbSjqkqTQlJKwxpSxxeHc19j5asfNyZiswuGUrMFJfPAKWb
/KuTxNZCHcL/7qAE/fYExtoEzlK92O+GmbexsGpgQBi5BhblfSpIdNgxE2uxL+ohBM1Yfi1Iv/4Z
u8xibi5nWH1nZoQyJ7AqGRC/mZeft3arCwv9Fv2UcbdS2VU9Mibx+g4Sg9M8QZ4N+tfkzTWXvK7u
lImRY9vo+d6GTkmcIOll+ZdnEjwOL37yy9lD1GYMDzwJWhyJVBXw9pSWS5aE1OhY96J6pYvnLdgO
0ahvx3Ljqrk+VSrLcrQkJeJH+0BnO6CyoRw9772KBSTp4PL6aGsXDumUk7pY1mIv1WFNqUwddnyv
z6yb/Tmnmf8zctHhTNonZtXo1F18xhKAAYoqydw/Vw0z+tlcqja6JkW0/ve0zH3sAQF3jiz2WgWf
kxfl3LKm5g297EPYt+r8RnBOJcCwWbPyNE/OHO/s5UZ49bxo1BwHaf2utOQGza/U2C66285PE4Zk
Rc/hdNbFyqp4QtWRkjCxQdmNJGD467D3ESrrZp5ip7vEqKl4boMTQKeOFD5jOAiYBX4wvR7XanWG
CuXplEtjdq9nXzZduGw7WzexuuJlpEAeXlpD1fK/2p06w5q75jpRDNzlioXApgipN1oq1Xt5zTq9
EuE+TR+e2zIpFSXlaqoAOOr3qX7LlywuHZbBU7ZTnUHbB+3/arfBQUeHrdhzyjLhCKGIJjleyYW9
5M31Rq8SszjWZeRvVxSF262YDWqcoDAJZBxtDVcKFMPs2y/UWEmeuPHrag1Cs+F5yib1B42mcTgj
p6Muo9x8J9mW40T7cJ0PmcQAAq8sroS7ppZBJPa7lC4dKkIj1/Mskn3U7PJcuhrLcYNL1xlly9w7
qKUfPcjfOn5J+CqjDLSsZ+a+okx4lQ2QeaNYwHhn9Vz+Muurs0VXwITRRw3Znzob+J24oTh8jZyT
XvnlueHGVd69hd5UjDjot9UqSmX680AYFMQoDtiu4H3AwQsRQr6w5O2ZMO5n+tcH3OQxBRlZ8NTu
Akl+r04IQo42KUjo/ZuWunlBrh2SDpBUGdoxpk2YTm9bqTVNfj0akVYX5RxcH1ogDKPETqB7g9Bh
37ZwXXsHhmXaTdd6uJwjlgxEGgpQuABNrMTngYHrhKwqLGy7fbU5U7b02cUQVCJ+VJMw9GDF1w34
90nDnKRymOudIA4hhxpYqg47BKlkNtWBbn10ShkoXwAElPYHH3AozuofXZjvDsWd7Til0JiclSFx
XNK32TkrGUoYqcdcu1Cvpq47OLXGvNu0i49FgtZh/Ii9izHv6Ona8HS85LXrZnpItyGOUAAeNgfs
Cwl5dv0kILxJlKViuT4NDKAA2glK3dZfH2yPhgL3Sf6zZcPUAiNjcbqb1+yttGKRnT5I4VGTFrqm
9/qImVaMDS5Zb8CiywKxZ+P1KYL1+Q8IQvUKmoGBcIEeZEM8iTnWq/6KlPsYfe/luS+GeCepA0Q2
/VgxL08lcwgUis+G6r0/SZMrVoNXa/SViTTRJ9F4OKYaj7sXF0CBfi+k0IdPnaC4crvz8jP1Goxn
0g8tvBFHeLgThvAgcjOksnFzK98kUGC4ZtNdfVsY82WSWBMPOKRznkTxK3/LexaX/6pNge+J2Jms
a2UPob1J0fJiOcgVuCXfpqnUM2EtfCH1sDV30ku59kbqZO0dlNkBPY0QJXFwuBei8Lu43ZeUFX3L
O4ZD2kpN3BehBsr4aXxk9faspbS2V1BhsImGnnpxMNgS+PyvwhcEp/hVoOjSZBnLolilWyxPYnyZ
lj/pTVRctbzsNJ5jViydqmUWDWg1aG9UCfpXgrxndBHU1mw0dkFJateE8XgRGXpKqu7MLiX0SJV3
WmidG2kkpA+B3w8hq6YabcTvNDFje8MzBodunsBSoQb083NPE/wJXnvd4br/Ozi2223uYmw1Eb8h
4tP7PDigyulzepKXykK+t7cEHdeaMbv+ouB1CXvdaH5+fd3orvX9b98AKtgwYO/2ZqEKWJOTWpbL
4tlet15KENN6PZoTRcbmdxaflNX93hjLauLkjZZyAGSjx2RryIEap/Jfx7bwdcPzU5zfyUD9dKkn
DKq3I18Ncv/ySLwjs48GwlNtnGfSolFI90Q8nORfG6EXQEXr0/Fjjf814GlLDGgUVMMyJ8ivaFO+
N1uoDzuJSxlOH5HgyZlCEsATNnmfMNOPCvifUzDZi9HOh2zl32oq8vtpCpKQcjMPIRxobsmrJuSH
yY0n6WmFmrB1OBZZ+6Y58bDC20sLFF5YFfzpmOj90xkKjiY1e9aJj6bfN6LVQQmdrATMgezCNLH9
Il1++691us25To1AkX60ha4v8juVW+ZcCDiR2mjoktRODK/2jxMQt+aGdJ+kXxM07pjoScRc5vAG
WuWgRPzU5ZX0XwbMzHVgJLX9q4POnBx2jiHcSGbqD+F15R4/AUBYa+N8wOprv9l4L36PWB5BizBP
QYax65ncyHmaRpWSCUsHig1K2DEXbi3kefljX1TNwdfn8C2xGn4pAM3urYFBHsoC6jZOXa3wzQG0
4NjRuiN/eXehZnmNKSMpxq68AvVu2J5hBKoQ7XEQ8APWsCwU/j+ZGaYJ58s1Zlv9lCaPS0zIFHVF
UxI+tvCcdfiK1RsFOImd/4X63MhF/zv88k947OARRTGLMC/SmQSkxuq+64DFwQHevYUaA/9fuwzj
/TM1vghhW73oIkFeU6v8K+iAk6R7apYIsDltN7soMWZHuEBjgU1/1x4C/BgmrCkPQCCuqJg2gLpD
s/Y9HUx/N9PfWjVJPWGFAq0IA4sHFoSauvavnsyhGh7HUa2LYPt6V3K/7slkgUxz3lEzn6EAjEND
N0wswtvU8d1FEF9YeAJfRq2NmY7HeuRgqvo33fYbEctnMHpQ5qEjjJvA4/mBpGwkeHIE1nZ6eEYE
hcuLOwv742aKdOCCUTsOoYn175dcYfcpuj0m41PX+ctc+rqsaQCJA5cv+0hyZ7Bq7N3RLq7rRtaa
SyK4SpWkGDNnpWCWwQ8XyHsNEY+R8zZbyQMIWMTOYaXlyjU2ZTFT3I8HIEXB72Z4LVP/g4Uau2Cr
ZsBwn8hMXKrOdI7+lF+vmtsNOd+Uy/sn3jY+T0GSkaWqCrqgrmlqG8ITxQOXgWXQsCed0eyJiby9
Xdd0A5JKU2V6sqt/bvDeTBrPW2kB4crMtIgsBqUG99gqcasnVeXJgTWaVDxFpNQabIG+jY29yo3E
CSWaDsLY1hyCTv6Qmh6D09tqCLy+UNMl26z9YHOf6aneEzimV1wMnWBlT+JcpF7P+LYB5P6nPmuI
0GpJn61sKS5Y7Xixtfl3d+i6R30Ob+eRgpMAJtaHww1i2uul/U7DXw84ayDGF/frGfTuqgjwpiMB
AqMjj3ZQW5SGpv+yUpvCgn21IgU87VAbyKBjwQH2Un7yp7ASeIq/wGORNzIYma+esFFPT0DVfs1U
8ZWWyea/O0+3FvmzezWvaFWp4gfijE9/mqR3ybXKgsJV5lor1Hx8PL7EeKAZ0SJz5HDdws2dHo+M
cho+C13o1yljb/Oc8SOjDV1zTBAiiIUU+f/DBatb4+o5VYBbTObB86mgWKSd1lA+XreiSZDjf99C
goLXQRy/XLzbUfBdgT8EU65ALfTKZE4JXqpmbslCg4b4vbqNBAPvI9YzxxV7Q9ZcWLGWNon7yzji
0sNnPB53nmHX1k0tng2EHf5MYBpGfwzXyEhY+Ys2z/Q165jwfcINwfqkp4cB6TpWZ7twgc9M+01I
tJ6u+/5BZwObMSzSu+IlTaqZOg9g6lEJdVpP3GP1ByvrzYVlYaE290s6PCqEAtGBNk9+Rp/ERJd2
WjulioxquBGt7d3oTKYU/aW7d1Ib067rCQcQjhThFQCrzh29Kaat7puPomJDhiQ+ugpZx+8HVb+i
4wIsVG5RA8/yGEIm9ltgQPeRb1T567A6jrIHqv5HSyYRKSnfnvbyCs/A0V5HtmZ25RWrqiXBQ2XA
aLbjc5xiOFEKDxI4W0kQQQL5+5TTz1cq0kRPc78HjM4tzJ3z4DtSMfUUQCNxJ+1hv61WB5WVgRFC
sM9QiMZrUMwLUPevgrhOFzI4FWraqNUXkVLOzpM7g6NHtYWIjIfaqC9l0YEmAC7hKqj7lR/iZG19
iPixLB2VuH89GzWUBTMlDxNHua9z3p2JXoXeKqfnBGBVXN0MXIwBVT9pZNXnt+ByU4I2/xzG52ED
lDQeJIn+Ee1h40Ym41N5QrWQi7g3Xm/uoMkMMaEbH1cmbsq64LXJE60Fxrfy91AR/BDA7pqS9T3H
0DM2NAKyHpfdbUtXB+on/N05cktGeY8Tq8MuQ2twBIPW+dBCuwK+QJu481jRJgylafM5ZZVzrhvW
X8zYWQs3Ic+G1WExAnPgmdPTmFxbV8SZeuVM7k/iF5v1mBYMHhTgT/5cu5lIXkz4gVYgbifziXRF
7IEv3TDG2qRrbZCcETJjPmGr98Bb2VuRg508t6vbTqdnI/QzW2tGqZNl2MFEyIAjkMsP1qCRlE12
emTo1vUfdu8x26TqSYQL7XLrBSAYK/6wD9faZ12QD9XpT6WUBNo+AcwQVL0rljnNZwP7jpz+zkNa
B0kg1sGgzlCNRp4UebZnEQNQtENbUjl4jFEWCVFjH2mOXDI5+ejSxkEbnL4fHVhzD2ga8tOwsNav
Yse+zeHtZ0UE5gCHs4hyNSY7AYTOrJC1G5n+TgtEJ2bc20aeysCIutpf985s+bkvVh7eDZ4izIug
67/Lc/YckvMqiB7o7GSvHcsHMV/s6VSxYqiYc2Kdy7OkGVgCvVorF+aUaq8rLG41cHUQvQRPpjPE
JZP/Y6RouIV+f0UFxu6cXNteHkYQb3Y9l9J2K2KxI5/OKV94ytdttBTfw0JlZTcBB7shS80pgwTH
q2/frO5GRXbNV5m1ElyI2PeGepw+Bfjg1a2UCQymfgqR4eImv8XoyPVyMiHdQrqcFg80ioEK61Aw
EGzVbQ3Zdw7JV0jfKxFlLsEmCMwB/8gSQ0QxaLSu6G+UZ17YgP2InuKREYAcX0pUxIIGR6PDqQOl
4ss3pAHdL+AXK1c6xRB/5LdS1PE1PDyTOU+RnROGJBkF5vyhPki15beV7EB/eul7LSa+oVYBLCDO
al1SuM7vOkPTMFBauewDDIHigM2PSA7HnzWbMZZrb8gMk+P9shSZJxQSuXY2c1SoEQ9LzjQdBVo4
hodbHYCA8nEQRbW1WIzu047uPW6p5eo1+nSvhgt7yJWjUAPVR7JSCllB9TkGk3c6KNcRUhuhbr70
eJMuwiRIEFCoMiLGcC5/4tPpaxUB9rZWsRGPFnEJ/yYZc7mgAjpj7jTtNL5w+MTQF3PMKpnuMaBt
H2/tNbumDweStxiElPVvINZGMHy6gPUXkjvRNTgerXCjmlw4QRqZt1FdVuWIn41OPGSOP1dhT8Yj
Dln85ROJ7BVELJTCc0550ZfPmyhogUhiod2sAFJFINYrdFzc08gdI1XEc5vpUjd8ofFbNerJhOuv
2adgjFiXSq8wNf1f5WAxpVKI2eVeLeP7KrOWNPERUmiHPmORuZ+xbxEWJ/5o+wvzFH4sKNqhJ+7s
29RPkKi6tmQycFc1Eg/HsqQDy62iV9nyl7yKVf2NsdvrarVaxsj/wCBsUuPXZlIfglucgvP/k4gS
cT58hKUZn9yLF9+GByfm/eqyIttYCAjLH1HRARgJ2XZ9FJwpOKCZ6WnNQ5w/7lffGlbW5xR0Ke2z
S9246VlPr/XflgcAwro/MU5sjTgEoSEtKiXc3m1izJ93+BABuBgakkJmCQFp64P89IUwNjcInjsZ
0rQqkgiQw0mowHO3WgqaotvJp90RYloWlcgkr5Qo27WB57Rs4KBpuImZYFptJS5fw8u3h2IkKDfj
KQ6x3eBmu6PmIxaKt0u0MZJs27L44PFG4hhzxiMKgql8efFxRjoAbltj9ddSWsPbYV//3JZ6JCq9
jsaXlXr4lXnGRqdzFSjBALAqbPgm5WnoEJdGCLVGlXGRwJVmCOhje5nSa0l5LuvStlqKBZ5FfNuB
086UgBLHdro0Y16Toqan4QDnrLP4SHKBMaH8OAkD/DLPVCIE1CPeU7WEUih7kwwX4rldVUBytqF4
5quXfjs2VSv13yzZTL2re5+9FpXY3CFXe8AMR2vC7vKT4NS44wM3Z24e58luI80YgVPin3hYyu9P
NW3/+UC58J5KsyK04KKVnIfGD0QcugDMOnQYwIiOLhnz6JRTf/LX2w4aXJdCWXy5GKmSWkPTcORw
yX4dI5gxQCE/uIHgYPHME4ISq011FFvXxPFoQ2k8NLDXR5hzDesiuBvhav5DNP7ckM+u3I1lbeN/
hW2uBoWZaNyjhq2oVms2LmOfnuXaKvRK63V5kl5APppGqRO7NBQc0/PhBsYvBLUrYh6iWlNNu4AY
yNE3UuC5E7l5xR7D57FSY3ZsKcldsQDePGV5kAFpKUmyXq1LOm+SYtqiujsval8pV3TeNYnp/dXm
RJpsEkDNnRWFCIi6PjSAvIxKvshhLmdHQYMAFTDcz++Rb/pe70zGDHK+8YQQJUtR3GewChRYPM+A
SHtGAkvB/Tn8d9U9vmys+jgwZM34iVhebEh5DdnfUD6tj6FhzB0M3uQEg5OLfOAz7iuYfvr4Jenc
nX1ME+fwcyyiVImBZOXWyGQ8ZrhnAp/AU15dzF7KFHZWqbNT7Rk4rm5/nirQbMNR3xGi5JUAQj+y
+QfS9he52jpiaNP/ld0fOEBCFvYc6wCivayDoIPSM0hc53Zi+jfanmAzZwPqcwgQogkeeX8nKlqs
j9CSXQ8h1jSIBBBmvB0TOIKyfGVjYrfR1MoDQLduf0x3P0VpyWrPpFnPCpUJa2f1eV6yucujiiWE
dAXOnwKyVrblLGLv6FZ31aOey0FsLl5EOGYi3BySihSbOQNWcBbfEQtKaCLyrMLj+oirTrv1/Xv0
h2RPQTcQqxQ/we/5ZAgTODYjEc+Plmz5OtxZHzAsaR0XW6TJnNyDyM9MawnUE4bJb4yuyt0fapZK
3EUxyt2Ch0/PyIQSd5mqzx6Ll6RD9DHgh3MU8jnKXKD2IJsr9LfZ2DRQmrlHic2subyHQidx/Q7L
jygWzdm4qeB3bt3me/g/CWWYoCzGXJsxAVLsLqtxFEElt15Ma0mWf3+H4jsBxJm8gXT4J3dUETyX
HzwsC7/uU+S1thS0wd/7ca5dz+Ev+BrdLHDXCpocS/f6A8XXBffNt8ikT0Dw35nqz+a4En8gvi++
+7Q2HnRjdSsB0JhsQnc12iXf7sN9vzAfTuVTaKpNOxZ20oD34oZFLvX9WXUKDk3yq9kGBWpW/Oc7
TXMq3TkFxW+iJ7P10k/X0z3WqgM6CH/iQb3Ffx0IRNuK8+pC8qDONz9J0YywNL8fKiP9VDyyz9s6
tvmtQRrjnAibNzL8RkQ5n/DEXuF5F20cse1KGjj6QKtushYibMaiTkB6qmd/3Ga/cs0siwzh7dzV
ZepW5+fkxYmcWSZeWpG96OAbLCQrB/ky01a9ro69HtucBMyD3ErSE0YPHSuN5ra2XiD2HtWzr+Lb
EKXkd6spkGLQFn+ikzKnC8+AuOl7PjGokMqHUWjYsd8jgleN8VC6Cm7RfRInyw8PdiSJ8wnzzIYN
vzNeplkPW8QVC6JWSDcP7zhY6RXMyUbByRUGxsZeXuF7q7d+XpzqHe/mwSIRk1+l5Msj9LNOoBjJ
SCvTqH67XMRTm7C0PXysVFNempc/9Aw59f5YAapphpBqN0JsxvPO5Y31eKVinmYSEPHf+j91ZS17
m4i112lI++jxr5GULMCihIJD9Mw5I+EXyJ9t+2ybcEmgHwJUPcyGm+Pc1pQyr8pjO6s4rcKEO5wg
BXM6feMco5wtRz0DdQUQg3oOgbj3v0F6YcUvyYbnCCHOl3kTAwBJvZ5HV4UByr6C2JXZb15vga5H
okIfBmAG8cDb5WpMP6I3RUsKOCl85GO6jiCM/s6Eb58AaF8152/yYl2AEIOmMLNK2qkSvevDFGA0
eAv1mnBlik89J4b2ODLUyFminaU+uFsGdHRn27Omwt2fsDGkz44rw2LWKKZ/O4yfLhY6rkm30WJW
DlmFU49BPYd7BRVyM8qyzTXV7XHG8GAXHLUpB6ptpqGCswnWmCn39khW/FkkhgsHoU5VP8Kwttj9
kBlMgvzGSkfLRvkyf0VB4DRAho1oao1VLcYh8LVKHVpQmTXCabmIKZ4MejAhqXjMwK5sEuPR3ovG
gnU+8wtZmkcR0hWcSKWoAgYNylr0APaw+nTk1238Dyz9zvbWrk7zUdeDiCg983pEaL7pnvGt815N
e1xZnpsl5boGjOXa/XHBMe310XITO711Xwx2kAwS5jgWr7ZELGTC0iwr0F17zoYMIMcOYWouO0wD
Tib22CR3LL/GqpNA32OktHrKJrPccAGyejnXmzmGaT28KnmJ19edsd+o1SEbf07cEshS3RIMB2AS
XR3iq3P+wZyAQkAQyfXitSJvypuiPTTjOw8cUCCpaLZLgUAPoS9JGW1JwWj1yep6K6eAnxzt53br
16DaANaUPof+87vfo+tk3b5vVdhxEvhsoU0VrPHfdcpgG2HftRcoSD8JlxPz21dwEFySj2tEibl0
LERE+37j87AZycdCTRnLmNx1GbVa6Jpma0QI0iYlniFobdfdRkoKo4Z6SRouLvLzLA4QfJwyoeKD
ZcNhuFWNksEQfmgqiS29jQWSF0Xt7vraRPToW4ep5pPgmVxHYMdmn+f6X1Oy6sI/ghXfaWMIoasy
aS0Ersw8Ch5LKlP8s8sPWjkYB7WA4I0tlyBefS/pYddVCkj3HVHGJQ+z6oUjC8vY4WGU3JAsh+2Z
v4EHSJXnFhozUpRKulp0MypF5pWBJ6ZTpOhOOq/YCCZDV5IZXa3R+mDlhlnj/ADlwPbxN/Nmdh9p
Y2wYrl9rSFt9zpzEmKpW3rUmVZxMicCxx0MrhLwUgGX3J27pPg0czKm7Q98v141BzrBUCUjTBlSC
tadUegifVBSRGZgq+DuIFHCnfhUrfhoC+gA3doQFp9bhXu81Of16K6CjGUGw3/uHEupj3yP1hZq1
S5f/9Z05BPdW3Dt9wP0Nf91BXFhFKNLeQSw0CFpfS2q0Ef09SeUJKIRN2UbQwPfYFUhVpkNNTtgh
MmNAKeYnb/7WqYsqOgAsrLJGBIXlWzjjOHyh7vgz7RjLptrkmYTtgBSTJ89i3YSwasEoM9feTHW4
503QxO8PgI8RcKTJaW375z3Jonq1H8d8HVkz3HaVTwKwPcNVbrjzGRZsgIHgNX9x0IBKkNXlevr8
ccB7H3h377I5hRxBk0Qp3i5kf0s4gnsluthac/+upzk3loLMl1heYLgrAmMZjeM1EV+TN9oY8v9N
KnfwiazXdxf710A98AoUIfIMHG167UyrczWL/Z/smYjg/OjX99AsIzwq9lOoPjXWzOM7axoO7Avc
zTkbrnYlISWp+o2uBrbjlQQXkQKj8RsfX4ALSvCPVZml9CAKqiM6HqH7XSmcLcBwHTaKCRWELcm3
0odx5P3rSDRnebWWiHqs+nXqflu6WBU4GtNPoUHM4UMvEKlylKC0ksJmA0Tlmn/caOV9VGj/fBxJ
D+/NUZ11l7yYaRWYXLFzZDLwqJEbmDnc/BbU3pyN6S+IXVe21NWsDFbaYFFvEM0ggsk2mNMpdgDw
/Kam7USgVnEyltya8sSfpJYl81G9B4KK3VpCT9V6HURbY0Zlwt/ro1rningBOU8fTthIa7Dlz9Hn
0h/TWb3UhF5FsbKCuDXlrV6o5PhGC3Hv7rxrfx4JOyitlSC9tu8FZr3+vS1ZDwwCbJWEakmm1qa/
+tHOCR6C2YosjJLbmNcMIWI6PAmUTy22PyharpwOy1SZqAnyybmIWzI29LBljP80HQqaN4IUxNRz
znFktxYdG/CUINNYQeA+1VJ0lRxSgf2NwtLU4LUSCpQFv1KHzBRvvanGYAB3sYjCns4y9f9yGv6W
oQPPh/8hcNlkwyPY7a2aCGPsFf4ik5r3FhaEbCkfrON0mmCquciWxkqRzRqh36KGX/52W+cMQ/Cp
2rnq0sQp6CTDVQSDIPftYPGFkB4PVrlf+gXTaIOgYdOVlc7CqbQN8O4qXViD+dT6c5Ew8+7dhne/
xGIswfJwFtSw3jsmFCd7QndTjqAKmxuWcOkVdJusXCs0KP99NqcyKC/4UXu0Kh0pKGlX/O8w5mzu
HcdmHE77ULKChe6FF3Bko3mL/qv+/ekDILMi3Ppqvi7XHtUhEr42Fbehf3I39ygjcLiPtouEBX1I
kpWxpezpPBF8VNA+s+w6M8hFSrGRiFVN+lu7Tq6CjwGROnrqlDfX26eNbJQpMBWHG5uMQAYAHxQT
1F+GQhWtakBAWghFuWKYlkyDIyFkOCdp33UNz7NI+qmQlNbXDhJVs8vc9jFzdJZDqSP36pLctVx3
HlNWIlvev76cJO0sCQcTio9TWJFj9scHB8mkJwT57hwCyJnSzxI9d6pd0fMJML2a+x0BkLK/K+A3
v66kzMPVu9LuxNjCBl1tT3mBQRdkrWcvaxj+fhEu9nkyfOlpLPuEqkuXU1kDOm0VPsnNm70d1kK1
IBqNl2vsDaVS05ITQnExrxymW58wKNmt4DsMzX3cLlWBvLjkuIHbrIJ/jgJOM2kFVjcwGrnyalQm
xoC6koNW14654jZ2OXIvX3EsZ1GuemBKAGZ7ACH1CFp2CEiR/HA7+yw+UONrh1Jiih/8RiFoxRHp
KXa4KtZiTkv3MFdzr4qoROgHF79EqrlgHq7sWDduOTupXkZ2PDiRnJyoGGtQRveDzffKV0LkBcHU
P4FPfuEoxpwrZQqDhsL5h56P4uv/9NWBJZ7bq3ZOa/9hKIup00MhHfkJOqWDyVN4YqneZku6SfFk
D0IQxOidFFIs3Kz1dXjVm57rD7nepdiPvKdVcq3280JOfWEKoD4Jqca8ZEPZEmZ1c3E35hEX4rHA
3c4J0Ml6mA/w6wTjy44NMBPuScPZ/nH6FqtCJ5lvqqyPjLiBo1941X8G3qPYvZo4lYd+FdKKqxyE
pBjLlnHu+2MTfuKUS7QN/9vxCHGhmHX1o1oG0qXQrPh0J5hNp8Vd/tWiT9xWNMI3MSeeTmKbyzaQ
BuBBGfWdI6k7nT9SehBUIXw2MlchPTtK3+mEnF/A4k6czKG8bcm0lx02lslaIp22WLbC1rLe4N8e
YFzg3O/D+kn0/DYv0AZ61acedbWO4+/kg4jdHWYbZDJkO8Ka8sQULcTrhY5sKo1QNJybn22BvKtk
/rUYJB2OauEKYGnfFoyumBzhAX4Wmyt+2ZmsEwbnnhTxHUVA6qkPUOs3TqeKN4pD0dMmEyh5cfIY
q26r2yAlh3plMhz3AVx2F6ZyVl3rL4uEQJmfgbf9CX/Qt/FlmnF6/j+7/yAieHgTHV0QV1KdDenT
80Jx2pgPMC+mW+sxZXMeJkVePk49QmDrlTTZ1DXbpqTs6DE5gnHYLj4FovDFXOBTiQv6wFfPGKFu
DFHYavnhKFyNPu9PuqYTOCz8jGZGDSoV88h3qxTdlLN+yV5XP8jlyBz5f4bZXUq61VM50VhfIK6p
ht8QYchBabi1I9KrFREJ7UaIqgAkPZ1cSK41yEGfZL8U1za6yofopoL+5Xq/9x2XaWI3FAaJe/7l
AEhCjRlhABSu0PyRzH1Uz7LU7cdmUqMEwGhjmQXq3jCOUMIUtFf3VUnxd1oS87ypegmYIqlXaKiV
35OXtGWTZPAQMGMllSTlOhb5mQEUU8lAPTBXiJNL/YJXdzDM4jKujS2fVGczSDmW+9phYQF9zOiU
KmGusX4r/qWm12GgAMzwWxqHm+POh+B0gOrTQK3zATvpWOTgDYThcJt1FWCnfleXIs3LsuByKBHq
rQSWE1VOsRZkFAt4B5a8gqcdv1wH+bAh5s6wnzZfA8r5CY8Ndqj59HTKIgToieyjSAt4J3le5YJK
JpcgSArKYpXAewDlDuQAGuRNiJztSYpn6uhRHi+xMIYz3GLsbFHqwMr/v0xYWXe2TLUUc3FTV+It
rJo7JdokWZgWNMgOvNr+D7e0K0v9TvJrMsNgUYZJTnyEMmnUjYzYiJ2r7Nz4cUaPUw5kj6qOM2m3
sd9lKM2wwXgNa7wsJCSJodYL6cebofZIXbmacFAb2RC79jq0Sv7GDtUHrVBQqD1jttxbrxuISS3K
3NPtFfgxhQFi+BqIQUEhOEs47VR/7UNxQAIzS696z0msi9SLhVdrCi66Zgzrk4+gPPPwVm3GRFJc
kNh5HE7b0Dmbw8DPV/5i0hxmMHW4CwZcS8sf3ldivdk0OpUOeram7Tlqny8oBNWEt+e0/AFFwmDQ
oHDfCGBPhFUw0GIS1XoLtS1pGX1mEdPKPyhscdJwIlo+Tog/3OaAjYMxqbaLWyJERlUdMfIHZMAb
4MkVnQ8SprLSUznUPRbkHSfPMxnjF+V/ZyOn5ZDaoDeDZtsiRt0nhafIezOJWPtJcj9ysJlAf6X7
boyZKeJ+6hor9De/QaZjrztTGwuaaEefFZW1t+OScz9TzYo14FkKkL5YJ74VQRg3re49lylHEPGb
yCDaBBJZGj39ZWtglpxbIWb9IXBs/w7lr1ewK1sTrYLWVWj7lqi3WhZYmF5thPZHddEoQBc8LGf2
FYYaE6qz1t1tgH5YKP8bliTvVXigXur5vTYtaAdvUUMUJ9bXqc/B3hnSm/QUzC3l+1q/xSYmyZqQ
QwuPDkchT4FkkuKYUlIMdrnLfI+6X3jSeZDKu4gKDPF2It9B+dlbdByEz7z/y8zk726TCjqbJAfs
2XTUUEc1Sg8N8MoR3xpPH/7DoCC8iwMZA2V4EPgVM3/kwmzDw9b+9MxUxbvMLz7rvFPEuxjg7Og/
ibfpBqKyW0sPJTUx4jUWxlf4VaGTS5U0UwxtTZE3X5cNvh7B8NyaACYNyJ8CCWXvlwZ8GWYypi+k
OlJuxR6IAPpIcUgRng/48/FWZnOCqC3g+VgOkOP8bpctx3rDU9CpZtLDurH9dFfA89p9WlNOz6jU
g2qvsH7oCArn00D3bZQ1kKeYrVvbM603HJqP0/6qiMbq+rIMhQM6q+Io9/Uhyk4S+tyX6vdPOaQT
u42ThAyhyy13XvVcF863vtSLDAFq71BxHgfkfoIZlCWZdAhH+4Jgt0JFRWKNQ/uKFJMf5MlTB3eM
37XsQ8DKLyxlHH2UL2vJcVY7MY0NvJBtHCegZiWSeCAC1Kh8BzJ4EHUViXyBU5gi72wt8HKx3rfE
VEDic1DhRPdMNv4fOQ9dcsYB19yhdTcn6ycGB2lQY917gPn+5oUc52XVulC+gX7NL8wBzntoPP2K
zAUTPiVJCN9lQxgC/YTUXq9BVbuwOLk9qG34lB2I1zUXzfbb/Ynu+eR7HCqyeJJM9C9shkOe+AS2
lkYkb+ADV2IWQxcseH0cbQ2lFau5JHUqGj4nXhzGkcZzTb1mybeV6FkkzA9AP0Ndifgj+HKA6jr8
vm4255lVV/T4PGFzKVRM7LYOUOK6BVXxg/Vtl98Kn32amv79n0KC1vRnHbRAzUF+IpMPvS0qSfyt
e3C/jCAxHQWcwaH+vTRbfHz8g3evQ2reQ+JE3Lj8Dk1Ri5JyGdkWjNT42YXnv9KGshVlTh5ijEBU
1F6C/QOHk9QPrNTeXRC+P75sPIRCTUGsVhvLH9l5yvamAZvOe7S6rGXnTiK05x4Mrii23s3Q6Ajl
EH6oy2sivO30YiUlEJmkJruvGnHsnB+NnW4CVw2anxs+SWGSYB13+BxKxzdtztz+KY2dhaOqyg5E
aEg2yAQQMUhNuT5GmzhbOKszaPrhhbhEKDvN/WaLzjPpad8GLXHJwSMEBpmCm9aCjlBqt+b0xUbH
8Resz4rgo9oVZTvmxheWMT+haeKoooRVT+uclXpjV4O+JeBzHdT5nJgsppH3UFPA04NyWpOb0+CS
t21R9sSf44Pg1tikyi3VP2NwWswZhocwh/ByGjXAb/b03+mFgcYaJgH5dExU0Y3PXD5R0WxLDQ7i
kzaCbz9GqPIyUzuIlb8XJ8hhPne5bnou4WclWxy+kvyXUs31a2JZVOq4uNPzefETZKbOusWBGr2Z
mUrfhviAR4R1Crl+TW9Q+DHmaUCkMjiT0vCIOjTgD8I4NRcixw7qD1P0iIpaXstLyrYG9dTMIAuq
0/Q/McOMPPVYIuhNpZxOHSHfXTLhQaa2twOTT4y9HKpA3fojziGk7qOJtwvDjTo9eQ06mdLAE086
3q84zf8rgvxlXaMImPpoYJc27E08VUpV3DML8cDq864BZ1VnAziMj8FzT7IzO4Z7HSZIMn9n5uuP
euVaI7k0gPH0pCoZaY7UNqMkt/I+BrYEBDUT2xtkIQ+jPl3lvTQl4mW9oQnkZNgx8lmZfTyMdFwF
pdlQW0oYSpQWxjddSNUb+wzG9oXq76RqxJsPIGdPIfLBg8GbE2sNwbCs54k5a0Z/B4uHQhuDYQGT
VQ9Bifa+Go36HpzJWl1flFYZoW9hWBK61dZ1fkj/Z0YGocxYKCa9uLFjh0PykCC1+vzgs7PUNZHO
7q5hWWjPzoXUCvoEqdZt7nCxDbQ7xgv51cq8sR/bHJ9n5rKX032nMlF9ONq4kCww+ROdGCIl8XTr
iHRjArStF5qdhF1txWYmAzsP7iz1FbwdZWRod86rH8PmNX/iPOcbG984UtHAzFoihR42RuI6DJfA
F1avrNdWvCl4RbTD5uiR431xlb8jyhI+hKcEkaga0PPA3f6oOhp62EKQu7jUxzZyXpNaUaogzP3i
pIdEZtUxR1eqIBs87SQfiD9N+fdF1byXR26cVcp89AQkBZzeBHzaz+yv+Gm2YL8wroh3Jm57UPyT
9HQO507I359gLy2GaAJvC4oU817OStgkswJxzCInZ05aGnOOnqV0rV/+4qb53hnyG7NAODWrDwX+
XNc08qdLPLg6KXulllqVrXqj4iWVy5YM9ovfsJTjbIk++/6OW9RNLJpAYeG83bMZSXXNgGBLuxT/
G8fYw92mmG2GXUepGcpewPTyHx7IdQcKhu0FrbEmXZ6LckuNzw4QYEKmwVRYBHceYyJGH5i2vHH9
zxcxXIvWEeNQHGn+PGb+NhLQOBmhW2ZAM8vASr3uqV2Ct5X1oELRPawKx2Ey1KqSpS0HWVhPNXt/
asvwU7xybMBXwnB7ghURQ9QALzCuMpeKF3JcVXhDJgFtOYVW8c8mIz57WRXD/ktw5ww3azQHqR5c
GJRyl9Yi9BWlOmp8oqN6DBPFzPmk7tOWXMeuaxxeB2gOKTDd7qVGJ/2GcbmNx63jx28Qmrycnx38
u4/t9ApGYYPj6sLCq9UtcqL093Mb0AcLmVatscQmINQbIHp+F0Od33mQNjYfpXN+x5wxME386QtY
arpjfWVcI+x9+OUv7UVvGjOlgF1tfZO3RRTilIwX2qzqBs5dvuUKPE1ISJCFCctggIy0GZM9neKF
ec92+Clqs6hck6ElbWUyjFbGyfuZzih3KxfTGxYtfgUQmemy4cvts2aoJaoq1zwBA2kWPnaR1agQ
oSzBwufoaWxjYZMkiQ5pAlTbN0UFlaVerSNihs0rO2T10FVVA2FufPeVQyQ2Jkd3Xm9COyXCJLWE
T4qcClLmU7vfDxEwnK/3OjKjy3QPvATrFvyl+qFrLhHtCVjusx68oEDTDb3Dq/V1IHwloHkm4GFH
/VY2USb47iQ6CXdjIGT2yOG+Uq6/oIKS2VL6IZehvHZpbhLJauKL1mJGa6T/Wjn1SwJknHgt26Vm
iFbNWR9t5i8LaL6KDxXpsovpHHrh6Fa68u7K4nWNS6pHz/uSCzU3h2sV4TqhKQh2D3irpgBcAKYx
gK1kC9JevnK4KxV3JlqEar1UCtV/4rECHyLSvCBy2PKycC4/GhB9KlzO/P+P1lbKF5FB+1dcRUJm
Xxeex1YgKcGFhVTYEIMC6Kv3S/n1Q/w4il+1e5xyiCeCeWAomhdgiJvzHRIPnFZQsBWCwgXhnjHx
SrSE47VHIU4lJAhlCpAB8fb3UGvQRhM6T+sd1B1o3ELj0vV7L5U9MN0UPhvMmZgyyvzwaerl+zPe
nodgBubzysOlsMYDQnhESBCyckJR7SHrlAxnwyP4RDK3wwetBMrN8DrD1kgwGeMBMkC5NCT2kah2
AgAGvinNUtqRk4NcfaFQeN0+DzoAdhrYGnM4adcsuNzZE7v97HWmMkU+jOp4GLAWqOBlbiXR2xRy
dVe4DuqozvOVtP86FGhVZtDRWoZCtSSH6gT4X5oL2urqgyi04p9WhAN+KnikNQSqwMonNrz2mlp4
yY4qZUyP/SO+sIn0aj5jzF08J8u/+KhFzbvlPujSJ2cj63XVYRKrcPQf4noNJlHSyHY7vtkEemCX
+n/SAFbIPBwQBHmQyeYfDSO+Dl9DuuuERiCRXvPsufsJziCqcug5zJZLiflHBjFC83KzY1+kXakA
jdRQNJnjjyIcB1xZ8fUXdO3nTL70ixP8s4eq1aczRx76Avym5F2otvn1U1kdYI2oo3VGapj39TN6
oeBdL4aM95pG6NEmXrXzK3bwk69Ub0VTYBue0+Fhm1b/YlMnkqmhDFsn+WCNOy1efuEpECRHBCPt
jjobOjHAc0txYo1zgdlDYwAWP72z1j2FTpLo6wXJntJr/QFMOQ+JBQCvVq0Jyd38lLBuA0O8Dmhu
BaqWbkO4I/O8cMMt4oYlb0XJuOjLvyWcFXzjAaYysopHJKc24ZFVGUwey+Q9WwCQI1ZxW0EzFti3
7BaVzWGtRGJKhqPC6dLGHQzibLbMb4Z/KlK59igPHWZXzJc3OzCRk/+45wRKd0cFumrkYqCA9bsN
3pgtKf1NnavlNbcEKnGBD5UFqGVYuxZRp/GLakeqWwaZHeCWzwG43pPxtht/+9qFAAuzbT8eWojr
b2fDHh8yU7KzSia4jDM4qqNzWQTWzMRTWYHeHwq9QgMtMjRIi2wy+KhYO8v2JTFtPKbLc+aPD71H
PXr1lDSppOtAODAf4iUONxPe4AGvp6CRuk7O2y2YsOqD2Kdycm+b+SGmLLT8Z1FKaPKrhT5VRcNd
4SLRtp0eS868jomeYQWeA1OIJhTGXMfFlNvWC8ahTDPm5k94a18ZywA7bOab3ZuBR+LKfX0Uh0o5
Sy6npDexLPcKdbQf4lvS272P1mopdEMI8yOxHRwJZoBbh9q/HBLeji0gUFrX4bOBaei9C4PfVZLg
b250KxUVM7onpAcnGr7KaJbzW//D/bcIPs82cf6gCgKLRPEIxmNDCEK5KBjhhXWajqe7OFWi+Eyo
Es7mk5EeCCb37c1+tglyRHbE5pTPQAE0xMlBenzhFttlESep5Z/L2kgrdvcsj48ShGsFWF7Rc3hX
x/pQ3HUAiTM1MNs6ecCkJrGLYrJme3FKIZna9b38Vb1Yvntxar28LRODBuZW4ED3jstmHzBEyph0
rctizJWlQ1jPJReQ79SXXE799oRxsuggDXV2fjVl/G97gSJwc/BBOxudRfvbKUEyYHPKwBVq/YW4
aTiCN5zJZlRb1gpazNbHB/V0qhHyOCudALoSarEfIQh/E9acJZk+VsL/Tn+JYh4Pzq+teWLsukxv
L5e7RM+yvDfYrdTWtwzVlFVQj6ywNIGcAzNFXtvTMJwZcOmp5mu31hxppKx0IeUHtIcFCmzLY25b
RQjLJkKoZ1nP4T/EfNFplfwZ0il3uOGd+Mvs+RgbQQOHECpoyJ8loPV4wg2dqTCgQAPFF5sabzEz
ltSpOVTivNnSEk5N+b/nhBONcBPwH3mKtYIMPlS0Lsu84tb03yN1WozjtvP0NfANdSY3ESu9k7i5
8CdJATUNNURivKM8JADypoKIJTjH/tmY1vqIUd+wZlhAwMNxf5UT/tHbbgQC4NeUTD5tZQUuS0qs
Szoc2BMBR1vhCiQygEx8Glj6+aFRn1lVGlo2e0ZnY8GoTUOeoBmHyRsVZyFxMmq9YQPNrTYhWBWH
6QTY+9UXMvGrC7FF852t1rOeqBmMqJfuhDnSG3CGujMTrd6drXpXUoH5EU9LIB/sQg/7uCxBMsCt
RUFNLKsCbx8YkKgQUEwFn6/rZs1D0mcQEaop5Pck0lRYgxoK2EEDQ7Fxe9Fdf7PLMgaDz4ZwEt9K
vRkLNkU3oMuh8fuabuG6qJd7tFdO6BS7QkOVG/2NEFuYSDRza/aPwqR21Ms141o+TLYU9m1Lzum4
dr97ofPWtP95C8/z1m8zaNkvL6FcnMr2MSe1Ay9jfWtkiY9Tt+cYN5R4gsRvIr4AzPwOVLYUxD69
6HzZKbf0ie31/Ke2JyvyHhCL9942hw66dCnpZkXLhDL9FYqUG3qhh4Qjllep4r2nRyLdGoE2gz4T
vdnATxe0V6n/zZXg3qCA8e3+lZ4U7ngHJKtgGQ8/66ZUI1BlLdOEv1MyzcR+sv8cySFTO3jBdqlV
oxffmM7GuQb2Wvy3es+9hXaYfdUMJQShdYPvAHwZ61AZFqPB7IM9rv5jSkgm70+7Pfn32pBoTQhs
VNyygRCa8cNeWb07JCe4XeEF+sjYxtrZLHlsJ9D+qIysPVh37eQBmgW44o5z+IxUNv2hEkIpOTCc
Bs7MityDCN1uwHAkw3g5b2dnYvJLfBy/hpr8zBWhDYxL/xTkObj3UkJcXIYeWZdmauDz8HEyQu7C
Z1C8hqcVofsJImEb6EUPYaSq+ZwR9sIxQWGalHbitMzDzfVDTxcTGync6hr1JTw1Tb0BFYfQedI4
jUUWZNwLXdRdnlYdKUp4ARGmbxTnsfw8gOq4QkdYAEVMYxCMqESlVKu+UC5Z5t4/Tz2zioJdWEmx
Yq6hVTvcs3T9iUu2nEM9k6hyhM8+nr3a8Ghk/gBzXmW2EwO0xlJeyF3clTnSE3ZbcrsiXf97ztQ6
tjTxbbwXrpQbj9ry63aKY6uc/+/BCY1VaZLP+nF3+IS1RRqwlJhEZsqzfpRod7KHoyNOGWUWw0pC
N4H4tREDsZi+VnskoAp1Pd16603mn0LyEBhUba5WjoUL6zqbx/vTA+6SkVgGrVeZBwPUB+ZMkKk5
1t1L6ZpFeZr/Cv7gxSq9liPRyP072aU2RZ+bNppbrpZIvdVimgHpDpFINPlc8Ge864XKZVJiclxR
23c+3+ObuHBdbLhnGdt3gAVnkxgrMJqQbYGo9rgeQuKKdU1WSHe4GJcWefkrb0ZTvwFDR0B4if/W
EP7FeBLI0eZ1MCTlGfCpMwm4wZfVGlx780XXK5WdJxkYuDpi6uogAhXUggGbfDM63m8x7RBPkMuQ
vjFlU/LcZLnwFPHkgP/c+dr/VlZDXrE/7bdvahJxdie/ahSJozhLqx6nFngNwq+NOMRqf/TtUar3
2R6KBkpokhPUFb6E+fPhnnNIG1Ssph4aF+RjZ0i/fzt0mM28pyLIuFQR40iuFE52PJSBJjp5EK/w
beUUGC4qlvYyJIvhMv+eNKgmCDmCcfh5FzMHfVH6s2PqDtvAo+ZXL/T2QfQPMwCw1hi0Eid5ODDJ
nf8bSMwQb3xCDFYX9cnDzN7n2rze8Y2XvctPVE4PRls/J2gQrO1QXxjeBKdqSB6GiGG78Ra+d596
/+q9qrs0RsCvXTf4NVERZ5rePiJbsyohFvBq5UKgFfmHDsIpCMQB6ldPz3/1w2626637mhzsXdv8
+0S1MifdoZoh71c3fQZnSB5R58CbS2DAyFanU5vYL9JQx2iHqVrtQ19xakYZg74zDyMT8QJq5zqz
c+ecBPyTmQx7uNocCtZ1OI3RurtojjOxXg32E+nQ006mSOxN9y7DCvWMVQ4xBSIsN3yqEfN/4Ej8
SJxsy12SSBNzq19+3k07EmRJCMGjlAFvcrYoV3/PtZvITrAp2Erpnai0mQ3Nalipw/E1Fz9mtpwn
ctpICaJ6DBYeb9E2DYprPsu8TbpbGisb040xKombQwSPR2kqqAhEekk9mlANDsyx6YrTKSmtJsRW
vsL5IrPEUP2XIk54Qs4R3YiFvMYjK2hMyquAo0pt41CyTXggFGUnoMTWFp7IxissydfWyWpiWk5x
Ys7pSP6wCTMfWow4r6k83liWzp8zIimpzD4KzrnYL3elfLNkivqvd5nKcv0gvWKCrsPMHjbEIDgN
7Ue+2Vy5fuhyXh34h2hP+hfWXGvkYc3mBUpOCxAEBCSdDUqpJCzZGAq/R7tghjIuAjrBSgohRFj2
IsHcnFCt3CNbpsenmG98+lLuEcSqD7lcTMCxAdwHN36WL3efXtFLHjxyrlR4hI34YwB1KGj5GuCH
Z9EUZIsGFApx2Q/Uywt7a+mKA6btGtFK8VkN/EzqJL42207zs5Ha5p1WCG1raY/M05nMZvJKEokL
H8vFYJuwFHv4OatZ+wdwOdYlABBStzbN2rkIQ03m7PydfIguHU9isH2z/ZZFD8WzIWBExqqWTtqs
/4BOGNx3f7to5oa15Ds90xBmDM4vfxy1Hio5R94tsmkj8CLDEVKsBhHNoTrHkSCr4hHtA8J4Wcc1
3W0ZCJwX41lzxxeeQ/akr2zs5M/DEkb2LTriIXTJ7/pBAy6i8oEFhOF1VvtN7XAHtchtyQ2/XFmE
YDrkv8s5BS5iuJDvTwE6lFPJTsJDqMrdShRrH+MEbgFotaStF5i2mFc9Se8+tdOt7EOm1i5c5I1K
J/WCKwHGe4HL10yKXTKU2Bpu/IpmT4U0zTzRDjDf/1uAlhy0LoNs2/+CQXaA9vzdy+OGqeHtw2L5
vL0LEeESgqrnF5x3VxmcrMfakmAiio6npSCBnY6+Wh4LVAnF0pYiRE8R30kpx5C7PUAWBRAT4wlN
bsatcbfey6eYPjRbQKtUFAqEwJy4LqjZBTc9Bbk2oxha2sy8galJVxUPGSHXRpuU6zMs69wMcLWl
wBzhh6gjycVWXqU2sWmKUxKxdRJ/EIUgjDDjDafouC7hSvrgabfWcA/+BHAIzxNEkTEfmvRjQGWE
KyAZdqj1OQav+hKZOHJS0mk74eNiyw+4s5eJlYvVnFhY65Sw2xmSGfU8grDhchcXZU1LV3rQ5/Gn
YPix87LxpJecNquY2a1Fh2+z8x6mJdl6LYm0aUCKQ2D3AF86rjWRdzK6yTEzBBv+4KTwA7ueKMe4
bIMc9yfc79KA+uOhnwRI3qtC3LnTLC5r2kMY0N7eckxVzkbQWkHxcNRFq/DX2o0dJozOTj1DZyY1
oPq8csUpVJAOqO0FGo9Qqv6WD5kSjf26mQDv4SawkpUx0Mru6ALZie/m6Xwy7N6dIQt4ppLJWRM3
d3PCaiGiDfsk7LvkKRmpDALD03WcnYV5oOwg7lDei7qjVxixOo1qA/teldIO9nJtmiTRYzZWSqNv
7RE885lQHDLGBjlwgp1W45PaIM2efdRVfMRja2j2+93S8R20nbHR3zwm3SsswdvsGBk0NKtvRkEH
f4Z5jW7uPqaUYvfdDUIwTXrfnNidpZQcS1HJHJvwF6KNh+qH1L07tUQEtYtjzJiN82I4TlT6za2/
+sG85O/9kgZ7EglSJoerCTxzV2iUdQVnoJxedEasYei2bk3BuTBjCLbwl4URqV3sl8myEm7hUV5m
eU/XFoL+kXPd1Fomo4DqERv31WYAfOCih8MnGQFsClc/n1k2/UXc/tVB31IBl9MlzN5sOfu+s0sx
kxJxpzX8Xa+NXelRZCZS8+xkQz5OyDhXcgIXIuoIP9ikk9zS2PvHpN1DEWviVebVrOGqysH6TDo1
xvPfqvy9NSkkNI+10u+o0pvkxtBZi2kAbRQtwyo/7j7FWCupPQw9NKhCvTPrDNQmC/jhVEc8u5s5
BVn9phHySFXZgWkwmV1WvakyKklN/+nOxZMj2Se1rFlkUKFbGPbe1czrIpWn7DGazsgbunfWarN5
zNms0cuc30eWVC9SPcMr/7Cpj0eqSwV6qssOxDSOKqH589HJsiu2giVBt5vNns2/J/UZo2ffw4v6
ch614DYO3aQ9ukVqFZTZ8nsDUXDYkYigwQrf4NlWV4Ew8mMInetgBQBUXCrext/usugTryRn+dDC
0yEoQp8tGgoXhVh561Ne2DG7fWmlL9rpOvXCmWiaztvgbr/8Eh+JdWPYWDw0ak/wWRctMgW94CVA
ndHLIwDcZrzRnjlag9yGopTq0YRUri273DmJHO8GaXFpL0Qo1hUXgriNFuY1hCzWZWPGXcgPRZPm
axRAzKXou/BgUjvzURnAkVT2rSCJ+Ym15Af0Y/d50xAfu2Y5LNQKbO/TuOkAQnvgdF44POLOJtiS
Mw9z7uYmVbH5L8C4sRBrcue/3JJugUjKnsaAbZArEaYkH/ALONkqSGfA8tPBZp7Btgbx4lxUpHsC
yP2LexFlFjA83ippFiJQQ/N3ecuoATD5GMmrU8tR8SQ1aRY5BGzsWRFT6jCLoU+67ZXxLiZmawRf
DiCAes33Q+JS7oTWqHEIXbEKSiIqeRR2rPUyPiMQKwie9TcXYOf0JDPb19wftsbuiEghl37VdSFU
LxEePAGRhStGKg440H3lQvOiEFIWT3jTrEjmctyGnzSF6E/GBjASUCblHsmK/lT715oQkNfv1Q7x
JOXqypbTunHlmMzznnxo50HJ+BM58Y0UKbCnNfdOoEo71XMkVU6REI7NCa/vROA07C3oqhrgzuOb
1hu5JSBtXveH2Gs3tvRKm3P8aDdrJtjqBvvNQWJ1mm7ftaGevACn3xQtOA3vMHRO7YUQDTiRlkES
F3KHF49XsHapeknTFvcS6BiYUFAJit5S+EEWqW+e/Y31Fw495PjUr1f6HaYSPVqAdxUAtlY9YZ3L
2H4k1MO3f+hdMi44vZtfHc3r3BUtlmieNBwW9z7xLUV98uQ8oiG9LozmwDIYqFW+m4+MdVMGLcZS
LnQmLt9083OkbJnyH8Wxy87Yuu85Iu+QUq2dOL3eM73nPKbQ2Wcc6mAdK0rZ8Xgjoi3UcDcElF2K
fAuc1C6onuErN1SWeBTL7HaLs6Fp7NqUrHTlk+7ULAfl1T9Xl+uwAeEXsgkmkg1+Q92DNc5hZt5C
znfaX/jfd8IklFNk3k3PDzWrwBHEOl++IgEb8c+KXpi5Jyq/Tz8Gzlwjr9STTohv5PtbyNjWinyA
VIuMwVD8+A7rB09ulGz2xjoU09OgnH6p9x6jw24ZVYLJravgFlFKtTRFgthuFPSUkaxJYVo8r/g+
/nRgS88MJvpN7Sk8DkYqu9Mk7cPvBB85WQ96+zxizaCY17eE3vJtE1mS2rZeYWNPx1FzN/dB1r0m
eXnr9BkpGzGMZhqpCF3CgW13fqK8QFBK/Eo/Eb2P7Up1Qon/V2QX+HEQodQLVY4V5E8ff2SYmwKS
8zdgwwkBGmkuXpuu2d3DMCzE1eOBvRCdzJxmGlBMLxDeg4QwUdS5MsqBp0/vVwmpdvfdat5BuIlQ
rLIdVhWjMs14rX7z56PprK8RQYHlXIuTlrRlA++gdsERYeLe/mmBvZeC0LnOg50pniCui9Fo5ePf
9e8Utj/Ok1/JHHPs1tqGiA3kXW3f1rITVwM4KHih7POcQ7AQrA+bNux6Q4d01EwubHt8JumU76Ps
3Q/+8sUmxeJbiJp7B2OdOqUAw0ICzREcWnSH/snRRdUafed39N5h6jwyocFXmSiKiQOZspGAIuKD
N9LIxShdjkUJck0R1pI/kKtvFURAK4jESAEMTzx64lu/VOra33VLcPY1seBDEN+SV/hWm4hstvcW
UdUQqwYzK3+roGyGehUkYhYsMftVQ3HX134LEEybRpy/YFmRzGWhaXvxFfBhPixO0kPArZQikKSU
AgZNW0YuZpxnmrzknmf4wr0669B3mZIjc9AS9YfTBFwogJS182XEZX6IjnkmXPEUWWWkGjQlPNDQ
+15z5p+TODRY8QEIvMRHxfoh8VHu+pt/sUfzJOrXiYvu7ZOeBOYxPXHiLEVVUP4r9zlVDnI48EVg
s5B9C2ikakUsqr9CQKpzGeqfhsQTsbuy2DVccPI3rSb5RViOsAXvg6h8wTjA6yXfF59pGGLMViDr
8q2VNpbnC3HcCH+txMj9bLuK6b+54RbHocsfwigVhTdJyfh0eb1Oj9Qw+cxL7r16k/MPB0+00ro3
GmKD1ibzMtECWgTnj5ZBruLq17yRIi+XiXyhv9f5IAXCf6mCEiC5JWZKA1oQ6Utoh9yT23PIcn71
ZlzWwl9VrySIy6U7ApTA+QuclhHePgsgeOKq6MAiKs5z5S8Lu58j+rbdN9o71Ws6JnLsnj1OuFx9
4zeNJCkzb/FtR6UgdqvPUlufQjl1168JxBbAip6FVDDuOZTgiShTGOj7IR/BT8aRb2IQl0X77D6+
EwRy/9i/6nEFZEvXgrHUlMiofqoLhtXsiOnxbjb4u3XD/vrbzF3+jnWIIITaCe5NpCyFub/KTiRF
jaSPXhmI6qtwA45nHNN7h3Hpaclby0cbWCXQMJp66XKYm3xEjAjHSnUu2w7+uoqyuF5z3SP/sToi
I/G6vxkEHYsf8STVUc+T4dwm1EQkyVrSJunnvP3Cuhoq7SofmLRcTFF9HnMGOJiAtT1Wo258683n
77WLX+c9RkR8MhWYpllD7iEmUaIyoSLrpTxepe5qrzaz+u6tZPvWYyX8ugWdCS4D8P9LsPgwXFBH
Qp4Um4WDWYAol5LtZJw5Fk0/fHPp19Otm5IyhpqEgWYXajk6TPLaqUdCm3mGDl1ohGM1jr+8k8Z3
CuQgZObRtwTTg6+L6EUaRFa1F4xNmFIr9u5yS20AXKAE9tPVQf1CHOMimM+0sUqq8Z8vlvg2aCDv
yW3pfY0a6FcxTIjKFTbTNXkjaoxhvc5LR26eTgJfrJHmcGrRJh8mzh0MsA2QF5w6CZLPW0lhH1bE
UV/OK+wuS79aldU+hvUe5dgy1WR4NTEYvlvo8or9UrzmulmRhJ+LiFqWOW/XcrZVm6Ri8Akj8uhb
HqvYS/NHBZlsRVQlrILmBwFBvECppOHOQJ8P7/Nn3Y/Nmh58xNpDQ5J/mlEyed0vycYm2fSspQG5
hdcCnWUGLh/TVdWoLKA1OhSDszQrxpt2sIu5yzPjvK+UjhGzRfcrgu2z6/Dtnz9hCDQuJKRfRp5p
F9ETcdLllcqhMOMFn2FSiQucX1zwDSHA3whN1XiM9g+ckR76Q3Ibpv4++HhTGqfXJrtM1xyEU7l2
E6ltEXUICRhQV7gU6j5xXjaGV7PKqsknK8hvtw1qxJLRScZ5OaFYTXH2sZIspp52kfEUJjDWLNfM
cBTyYGsxDi/STyGq43fHkFwDmHBWE2IQYzN1vhTLDMN9R43++xsrAvTV5UThriyNY5ZOlBscvTxV
+7Ml2wL/QQiogaBKhiM34zDO1L8Ju5m7EHo5zMuIX75RULMLT7SUC8rxTWhe/c9UanFowxcKyRSv
h6zJf0Ptk/9B1g/85nB8PXghKkdVSblpacBidRpsiwJnfm6RsIFCjLMfNVU4KqSFancBubhNK1CT
7LDA4/G/J38+yZgJTw+WJPZMdQvY2JCkSa0+vHdghPl3XNZ3gWiWBYcyH1Moj74x3x7PTZBb3eUT
wYJVyoVs+6mH4GTCMSzGN+xMmcvXN/OoJZetNQc6IPEw0T7akJOLZTsITA2wlpcniAbEuxYYNR73
e5u3CIQ/wHmzkk3EDfE4veyNvxTED/EOomejP3Ncp4SQ/1QRsU8IUKBsPZVvCbmPWhnypHGZpl/s
r+Al4So3FstrTAh6nXWyXEdMLelrQUxXHHJ70NpHa9aIKKngaLKKiUilt9Cs5QcecNXVi6ITDLAd
lzBN7yF90QHRky5K2AYP1BzXxjFedUy2UZ6hR1lAj4uuSO7TlZqRo8QQkPcixyHlO2g2nRFq+hLJ
uRWA6kw1gmofk6j0Uv9gKIn0Uf8y2CMRsmyJ7dPgBotbyCiblKCLe+avq9OamKIlENJhn714sM94
KnNqF2/0krKkLw1a1yzHIhOq0fAuXARSKboVnNYAxjxG4+p75Nr2wCNSvRrM5dcLdU0Uc1mWniD9
bCsJvGLAVOR2LX/0bNL9Zp+YgO+Io3MeGfusTTXrdqxBlVZay/sMQre32TXMLMirqDxVDZ3Bm4w1
F7dIyeVNgKBAVE2wN+5SQATo0Vk4Qk/nGtSETlUXnox9EC9UMkO5eDj5mTtnotxMU4PN8vijN4OY
4U/Vy1UzLhFrfPTHLNrbulI4R/OAPTNWwHUDMslBR7CEhbkqw+Bh+vsK2LCPD07AUXbInOkLxbU5
zFJk60gmqVAqOKHVkzyslfB3T+iNQh+cqnKdh6MeYAF0iS9JHkSf8dRC8KkhrOT1TZSX9LZGuZwn
hEOX8SRiEvIfG9ln8uZPj8oP6QqvX70u0agvuvDTmBVIu13Dv1jFWrehTwDTTzce9MogsB78SDno
4wPhj6tT9m/Jzxi/2qEOGcyugbGaqsVWg17ibFFWzaUTK1QtrGcWEZEDOPmwrdnzG2JWvZtPqg3+
cLWzPRyfr38E85GkZj270tjp/VuBejBe8PoOUWnDu86MTB0HWgIROIGhRt77Wgqaw8Sw7h2AKd6B
r4HtsZZdgFdgfk/fCBbvFcm/Ov0jpDT1JDJGU3v/PmuQn4RlRStvQ94AAfTgFQrU3qv26QKu9lsw
l9iENlGE6BgQ1jRzbcox60Q1JTQ9SCJ9nGVidIYF+GPCaQT+L+1TwxNOy+6sofAf87FlhqR2baUJ
WEt1pc1YKNFQNwZU8UW5G8mE2Yb078Xh1L/tyk5IB1PRinjJly1Nxz2+IuD35cVoCx4BRLKtlOw6
3EIch0wKt6szi7TnDme/Q6J3rO1ZDuPzWM3lSIHu+mtp8laR6cf/d9LJgSjZIGGaN6UAiQdcsnIE
4DAWUQHSe3qEVHF/F3Pd5x+dYitQRZytZtLj8qdkJeL/YvjlD5tSVo86UrtCIl+4yAf7G1c3LSmf
PJSbhYOET17QNwxxLURw5WMRz+1dMO8xc4/sCqDVATzh4N9lh3Oqf9ph62VTEVA+56pv3VPlvgZa
bztKeyQbEcV3gHKopb68ielwGCP9NWNgKZOR25XNZUdRNooHIf06QQy/+6WSbj8PvHze9se8msLf
BDlys+k+TrGik23Ehek/2otA9Xfd9ZsmxyyRW7QMNQXsM4vLIwHKDFhHlJLVeIMaPApnvbTa9lLc
mUbzf6tFn8kHMglpzRqNpO59qm1VSmQ6RnY/NAisbET3uEyDml42bckleOx6zlbBo8v2v2d18e1W
qRfEibCNrhlUcrJHqEuESXNAVzL5cimBZlpKaNF/+7oXDcXGLTDODshxTNHNaxCeStyMB6xo49GB
goqQtBjmy0qo0Y55Da4yMoqph+ZofEbirZsR2Y8XXIM5Go1eSzuu6x/dQo7KTehzx4Ji4XHPGKe8
jSmguE5Fokh09on+lPTIztckrZxTgqkYolVokBmL+d50PA5nc+uTXQtW+IBYUlex5dUr8OBbLoef
8AEy9aBc1sI+6DyOsT9QWkwERxHqRRdsPXrcg9ON9QMtUh/L0hkZHq1F94VjzHY3xnw4DvelEFkZ
nhc4uRoxe8Qz754zcKT8zG0Cqh14OmlH1jn3mkPC7D5iWnfVdvXX4ospBdvutAyrjsHqGqAjsr0B
lOb3hJRZcrMa1L0rznMaUc0hx3TofWGtADPJFpYDkcCt7wpFT2WwmGt0qI8uA9jIgautRlgJqJ1D
WqeBAu635XhNYIJzWd0ClUeNiCxgykAQqDy+3MfDua7LTUiuLDFwbwQR3JouJr7s4P7w9tEXAGV2
+WaqvlnKeLD8F71nulN5K6/O2yCGzyoLaznuW2wAmLZUJFhj7xVIuag6MCpDRqwWJUwwEuhv6A2V
XPRdLEP8mpSmfJ1VoxtOuFNTnsfXG3n3c4UcbvEFEf5s5NWQfeNFo2pp2w9AAPiWjBLcGLU9cE1V
2oOgAKTcDnUKaCUKpgDqc+Ufs7bsDCnWN/oAuhOp1/v9KKPQPK6nL9RH1OW7w1fEuOFiHA+h8FyC
xmfdT6tr1EHl+l7EtK1t+om01128A7GitwqdYZrXhDxZ7ncNk+VW04f87UDRgO87Ej7g0dqD85I9
DNKs0Atvd/mRrlAbj0vNQ1s2RmjvMZnnTNSQJGOcp7luUz8I6GQyWnlJ7gh6KGenkznGnQK7pUTR
pXLIQZLNHOUuC6JrFMIiJxHDDCGScXW9pTyFLsAOs6ohNEB8Cq6U0ncCM/kru5WJ3rQpWT5k2u0l
VOyv35Jb9dAOiZfR3Se4bu2ZE5lJdhgEpFqRESKRO4xJ2gL3UvmAqW0jLw4wk9CA1Sk+ew1KwhNI
p9EMxk7nlbL0gC2msOIo3ivMvU45yQ50Oobfq/E0vqcDASjLh18K+dqeJ0pauXXU7TosAao8h4vz
I+g8blJJ1mUuKtNMgqdYKAAdBOubL3DQOnPTuax4324h6aJNokUZxMK3UkGLlHYXFWz4g8I/hhK5
S0JRh127lJZAdwWKOPfToVc4LpzvM1QEw2ly/ZFpkxvrQvC/vGwJUarWuY1slKpGUNJsgCtb0ze8
CbVpaehkHvFF7dSUcIDdJ2A7CYVjy/sAqxkQcJHaFG2etb0HLMJmarOYpzlcKWY7h/Q9OaS8jTQ4
AUjM5JMyPPrX7m+l8d8RkVXwvuo+d45xOP5msaISK0Hwm7Zpq25zuIpUWdZjbNTABLJ3a1SNmVIw
1OJ4oG7l9ORHoCbGZI+bb51tsL8xtyWwU+aEHH55VMX142AIX7vNXB6tpeE/RXGG4hjyC5IFoYcR
QwY+TEToThxkdr+zlL8xGioPJ7yGxzJmc2fma/PPirpRm8N47/5fauA7vGKS308Jk2fL5JbLL1SM
Gcz5KHId7kSZASMoE1snkP4apx+Ydfj4PiVmbxIXkNMBqQgB8L0d+6iU2wbzmXkxsIi1Gn3dE4Qk
TAlhTSuTKJOLg1quALw5gnIo/y7oGh5Haj3x8SfTSu4V/kmMdbWCcHqz/Qc6b3g53Xr/q0MAoiN9
cMVGxPgKDZRqVMAeLckYFivXODj190lPiXmGPKcTDTd6ezqoQxMj/8CsvgejC+dlAlWq5ZZITMy+
eLdwHtaksNA98fQNgnl0wA4DpUqB87HIXZLMKmEgNh9z81eYNWCApqJjj9rgvof13WBKJJ+SsyyB
hTJPAUT0fuzf64G5aDrf3pfFTJ2qq/jdHwOc/RhCq0mhXA1YdeEcqF/rkNC8TT+mVzoezKVz/zeK
9OiS46SRFazopDiYH0BgRwbFopb9J3xi+YoQLMndat5KnX1XkGDRaAfvCuFR0SENRa8PqkdSi4Ha
csxSnzU0kVnlHFMFqFJ6OjFZt28chTCQIBNKcuTpIe9RfN04fVPM+R706s8vW4G3IDfe09Ivtcw8
v3xdV05rX/UduMHwPKaaV9+io9sEo7XtDUGBiMiGyAl9YO4nTj3znjZlUDb7ZJydRYRrNnq87iJT
oNaLaBBW/oYEgqYf4eOfSbp614hlzlrDHF2W8vrGimzzUcl9nxWRW30PSW+30oNtOtz7o1MypgSf
LeHWd8d60o3zXOAUdPEloQKh+E6rNL53T2pPbYo/0a6TDYCwYHdZ2Ll2Ra0JipxLK2kDMnXbFV84
NsBK9h8eTo/IuXiHVNAeYWpvh1sztafvE44X4x2nt3fONU5bJ2af/H7WrSI/1Bc6Xb6R2XMc/b6Z
Uf2JhSvoVXUSgeQnjUsMqrQ8C6lQdYkPEyvpObC1wx3iGlty4+cESaoQujm0+CShpq15do1ApbWT
1QF3uMrFsXHZZs5tWLXqaMOInrxDkZo0KhQYG9GQlayRQb/EiMsk3IMvpUmJox35CYBwJ1t4PS7D
v2ZZvnyzxRPDUiRrvk+wl03iUL8995Gqs8V5yYPWGpW2FoKnEHr3LLiCUNMXVJcuN63FzJAwSgwd
T3V6SmYFodE5bRRGmlplC5wxdua/acDevnGoVfGH9wptrKJMbWqqQZAvPvFyeEPJ24+q5akUT1nn
+dgnBSLYqVaCAyaObMwt4uBNF1gBDv2/8Zo9oovz+1X8vDpFyyN6KbyYMR/+XiCL2LD8GgUkVAKT
EQu5cNL5siGL85mDyh+KBByMqmg+vNejbvKDZlDRfl+5RLsjIxHPX9Bs97Dbaw4pqR9ezDnuoOyf
6Vr1O4uogHKOaDFLLhn9dw3y3JYWS9yj+xBqFTBgezwqV6qYENWKNspEh5qLz8+muk/E6Bm5Um92
SyCfTOnSq3TvjR9BEyZhgNB4BDi+DJOlHF18cqulUdqoTzWydAkB6I3dJamREM1Vjs90FUaNxd/s
Gi3rWwfBxzjPtrqbUMbPCdy9LQXa3ty47WaIiI8xhakIVDwsR5DyOWlhrpbN6XyxYVDXrxijV5ZG
Aoh+n+vfbv0a84AVlEB42NHIrBBJgCDPy8UbEc2F0KCE05x3L16jgthemcfLPlndXLao9Pyl3M0x
anAC58kHBodMBadmSRaNAHnvsJ9cfu5QsKAFMKZFTn2BwrXWEPtqEB1dx/1F23yD+2JZQiAM++Sl
lyw95URykZiJLyzeVaQaZqwv0TIBxqccgS/zLRsQNtBEBoq7tG22ZvBhH3fwRO0MMBOKePXtqFPw
kFqYYxUBGLKHweeq7/k8dnxI/A3DN8GfaLQ3RKrO4o3YC2tYAvdQNf1FZYPEH4lr2wTZy0dy2d0l
cUSLe2kGyolzfe3yb5xdJJ6HHCHtAfyV8/NKISnrWSpVP0mz09TSJnxpag4X46s1xELkqjJBB0ci
qpsWXZl2G4UJIesFBrjnKjRJ3EVw6MmCWAiThHpdq2/bXqlNBzie8QO1ckhit2D8YnCwa3+P+eej
iLvTXz1Cxoj40urm8QGxptE5NexS0wWhCbWBm7lZJ2DARyjMTRUTgwo4+7xa7QuGo7lC6kLQjlgf
LLFpSnYwOr/fH8yB+avb5ZBjWX4+9D3YZYifgdUc78j8oE9jxaU7UZptX782ID5LYGl3ZG8dT7dd
VtQxQMAv/Mw0xCmX3m6C7nRQtIJI9M0DliHJe6avjTvNwGWkvChUqN4eHToetgIxchL6iebnMPKW
yV/HseVC47mKXzRpp553e8vfthmeoHIW+Cf7H+6bH4ANqjs6D+jln0qQ5KFs+QkfsfLCwB8N4FMI
wO+0Pa6Q6q+cJwlhCqr6ePjXsC+KMuJK6o6OCWEyABv4ZclD7um7t3X2ohi4LA5c3QX5uSeHaaiq
UzlrVsO1b535JOOCBeCpCFn9aiyFRPVjcpzoOeRWqrQDhJBpGvZ2kL2htJKWtUolrn2olPg4OHNZ
WsS/b+zGV+eaSJsmEBC0gRgm062Nz2L/6eqH6Kbk0z6/VGZvzcx75E6i9nQMYxShyLXr7c6mPkBU
msXn5C4y5cr9lNtim3Yr/oX6tamJWvUmjdz61y6cZVLqjIM7TBqPyNS5WV4EQ5jMDyUs2m8VxaaE
i68IQbU2V/sNNToPX464pkVMTxIUFKxK+y/psGfsTUuWqkeiQ4SMywiDMB0fCsZ32/+4/Q89OLmI
DfedLcBCCt44Owa43hqU+3MnDtJAvTjT75pPpiG38DNpgRscTbEAw+r0H4kEaQEPMFK8EigTEweX
zsSc1uZVYKIjWIwpzthI5Nab9XYTZjPSZniyTZj9pbXoXa6MqVPvCEg/AtFSUa4p5mxoYuO6/SSG
1A52V8yCRblK52yBahRbhzPaldiATxuASOVp0uIeEtsjCU4avzANYZumJ3ESvuD7Nze9X9pqfahO
Kwy/cmgE4SI6k+t5b8n3rI0iGlspFbWsZJwJd86I+USvBpQvew06R0NqJTNWiwIujzmrh+9rtTOx
wY0xijKjOLClCeQ1E2En6J8x0JWiYm9HdFUoMfFYlZs8P0g5IRzaf4MUm6g22FEMYJvRnlHoZyiM
Mjh5kmV7i8HYbRqJ32KEq6cLACb3RfetYpIo6Au36vXt5GbKV4vHmEp9AL7EOpIISoY3htZBbdpi
QnX8NvVdUdsITMHWHIqCAvcxkmtYKPOJaTQIomqrzGtDln2ZoHnmVBiFkG2oHcmKzLn8hJA2CeCC
2znVqy0r8nf1KazoFA3m75dTQYqdJRnfn8DcT/J0tm/p5BvHYvS5iqSzyBf4jhcn9xvu8zxJuIcp
mnBxa1VV0icMNsrW+2OswdsbrxNIcmvI5yg4j805QvtLZYFvNqhC9r6HpLchnVRuiIofwf+uGf0T
m35w8khVbzXZENNKhFBn4izQwzeD1LXSUinwKZSj9jH8UqE9HV93Zm6tZEp2CCBj2X7Y3Z5l4RgV
9eoFeu2ufEdb3btvKFeLFfVb4CWvN7ZFqbib+CAiDmv4xNVP9OfNnFZKfF2h/Xx4I1WYJuIQTVmV
CUtbtJWpDswErltzM1S8HajnGKozsbPYBtFOSy9xEv/oEk7f1BJ0aJ8j8OlktyBbpJc+KHHB6my6
bFuL9sped9SmQpnFU9gq7RHp1Wjn2qPaE7fmt9Kpn5mCgA7DbFMcV8s6q9FQ26C2MkdYi2Qfk6j7
E+8eiCFHtpJ9FWoBvRerVdf2/F00wWrBkSu/cNrG5BkaNwF/RR+7pwPcCmCr9OJgl7aV1hcH+xWF
2ipdFosd88Tn2G2hT+/LJQOtO7WSxQZudzw+O4Q1sYlNUOpRoR7DgNcgdb1vKzZ6Xi5cjMfUAalu
aUm4FiSRhTUaoyI0N26bl1JKTJpCj5lLXBj9WAW66oBDVJH2JfasBe1sqYb0bzDJ1dKfjoGeEF3z
1SOtZntbEkuClyh5SKxyEdQL4QmBSrYIpWHjIn42YVr2CTBOO1rRP/yNTAHvC9Js6ItvlDrC6kdH
X2F576Tad27v1g2etPrEMAzY73RrtC80gqgUjKdDs9gU0gVHwNbU2KSKqPBBLBwxQAv2WU7dsSdm
Ycr27X6APKknxuSHu2jNxxT4F9Ojuodf27WXHOJrA9lNdSU/+xX1s34NIE2fUmCPesz6NjmgR68c
VKLW6ojk49mHfXeLByoEQRrghrRXtxhmJFLaCL/pozGDP31r431vQBI7rhddeF5foRUyMjxHoNt7
LeWTA62gBAiKq1NfSCGv7udi6PQd2WvLIjAJMMSSlQdb+SpEXjbZXa32T44bA6Zn6pH3bDcO71FJ
/kYH5Xia+nwetNsSpNwKW5HhGRtxQcfM5bG3HKnlJCYRUcrG46BvIV1KcDpIzyc5Tvr7bRG9THy7
zv7u+P1TR/5tjj8K/Kveo/0E11J8T45XeqT4GWshg58nCq023A+f+/bUYpeSM84wxgtBikRRI8Nk
paMjFEJ6RyGpjDW7owixap45ggP0HiHktNFx+mS+rkOeSc1pV7FHmz7u6yZOe2UsDrRLSFbRH+KC
ZX/bTPIsyyfuzbGDNym+WduJM1q7vks09hUexXMhnegSdBBuU0Ij27wdd/ndNyEOCHgiiediioEH
+VhJ54+JXaY5psF7z+IahRmZt3nhaE93Vr01+NDpt9B2wZ+wM9N87R1sYfmCuUPoszU39C+Pi3+c
SkxNVeVw2fqHxowwQoQ0/7BKMXsJv0rNErFUV0Z44BcqD65Iag1H8+mtguQpvTrADBI6xjI1acs0
c1QkVM2bdEpj/N4Kwk4iYdu1gyB51C0gKzQwVk8O2QIYnWThqK63Fjbp3fNHyU5B8CKAZznrMK8V
j6IGx+GEvBEmu2lfp3cROCHnCJhyjJuxa95Z3e+YCWhZdcZDb1vOQamYOaZqrP+ipX6X+ghNpd7G
yeIePO93D8mXNWKVleUPt3zYdjlvxTk3cwsu+QPZZQhXc/QJ7QhXbu4wDqFXDNcts+hTcduBBOTa
8BCZaUby1L6AFYuFJl78An9KcJd23roHFbH++viSVsxZLUMixLRXnlrXQDDcSjbL76qNcefh+YAO
+xvMnBz+vpo9QzPntwibNNjissK50Scf60yzyEc8XtLUPxvf7GToXfDOtl4Tpt0zY7aw2MnGpBCJ
Ztn8HIw8JjQswl4rq0QhWTFIuMTSZ5KSVlCuA8DULCePIUVozQdmCcSp9PmzJqKi19d1hp28gGgt
CfMTgRXJhlM98wxJCZaY7rMOq+zCMg8aB+n1YGhdB/LlwrsKmAmHoERAhLi53WCOeiHOuwZcdUxm
NuDwrUh7Hjm7S9whlB9UKDSPnf54+I6IXHcHjpcLGafmin1FJaV3YM0XZgUd5A3jLUjZIr3NW2Py
oc0687zkRKFO73QpPKyt/0hqzlJT5ud02+ltSD4ObzKECDAbW/vVJRgL+lNTzP8SxwoLchPd+UMB
vID90TaigTIV1TxU7aKvWeFV56+b8jRe9IC8IldukEHoqFCVdEBT5HxcEaMZYNYLaTjkWLv4XUFU
qzDHmEd9eMe0vbXmZlDW05CHAp1778JxGM0G5VvbvvEsu+j23i+JU3v5DqQInHZpIqBdAujI9ZFs
6U7TRoHnIDBARU935PhYzVQ2N9A1O42Ag8UEYR6l1zHEeYoh+oWjiFZEsEakrKoQ1i+rCrBZ+QOo
neZOrmw64l8E+gt9vGrsHP5mzbCvQPT32nQOMMXeIerdZ3xYYfy3dHAC0WpefFmKDgBjS02N5R7R
i5Loh7E6fD5j0FsoQN7p4Wdsi5thKOo5sPskm74UeDkXgPXqBGR+IA8ze9t/CteUQAQBTvo3EQwx
xPBFh/ddqvvnKMA/AzrMvTe+zVsa2GUG0Qb1smCe9aaUlcq8BmyZJ96mvHUCgX9LIsDcFhoz2th0
vvUKV5DBKfA9ctcrNqRymXT/PXnLr25WQYDsHCkSkpc55Y4nWW1VgP0Jwdh5pCEXV9rNXEuheG7T
m1Ck8SSef6xi96Jf/Fn5XPrDbOSAWtFu1q62WQI0SCjFCHTSZS+AidA4ciFH46keWNrEoUyMHl0v
0jSPc8DSJ2nixk0T7xR+jZ3/ub5sp7XHxRLwCeuUNfNw2J2e67yrhcT7ooVcDqY/Sr9oCqpECk3G
61vnhYgXPxUWX3yC0FSKYmeFgjsp4nXR32r+C+OCoerz9ILixOtzIDgaWHJwzehLgfS550+UA0qe
7ycUSW5CmKqZBX09UBLXG2f1xyM+EMsEKAexOEtxoJ4F2jYfkhLGwRcSS6WES95QLYmivmZdmCYs
opLMzGuv/cvISNFfCvjK3nALSqmI2zpH2b1aa4g0x6+HSwc7BliHjw5AQMH8n94iAaaTk+gnDEsv
6CK2dAEGTAYEQrLYdn8a9vEx14tI+TzK9l6VnWUDc/nt+hXPHvqyFHEy2egpVrwgobT5WMDbHu0s
b0mq3C/BU0bd1xuhch97R0RekIJXYgC5OWFj/19eXkLdbiFa6frtBQii4zbhPgAlGvQ+J2CS3BFF
Hdnah58ieBoP/vC3XmIUAXygBnPzeWUrYtQkogvG0nINkabeTiryNzRD/vyNNf4re3P3NN/5nD86
f32ZwObRubsEWdV5mGjU6LQBdVmeWvIwMF/gbYkmWef5ZrH8CS/gQJ6caDLUslRIApxV1zXQenBf
p2bXbXiQSfs5hx6bmA5oBFlTdQEmzELZAduD2+sxqYsqLL2hfPNQBaSNKe/HdudHRy30ROFTCtW6
Km1vFwLwmo8N4sgqQWjoHZMilMC5vGLTSGdfXwJlEa5G5/TE+bm3hFtJ0fnQseRv3DBwKHamTUX5
AO5fwjxbcsodXrqnWBBfmd6a+9t1CXu+iteiFTqtxvpBU7kHtaBziQNtItB52qQ0gsP+w1jgzQzq
eDyXOMLf48kzJZoruWE13YZSTHi5JMU0VulSpWaUiAYxBhMcWzdqUh2rWjQQQcHZyDJdfluIO10M
CyC8I79pUNPzkmVXN7jrYxYC8FFlGMVrCySMG4U7/zCuE8agYQiEAb5YCWliXhmqe6xxZdCflvKH
F+RoaT9DMZJakFXcfn9ZDPJqsnf+4DPoJoZ9tP0bSjBooxpG+PqPSVvEHWQQXJm50MXBNNxIAFMz
2LdK/4XmPH+RD6EOfw8dzUFhBYBPaENJAlyc3GjMLbyUPtC3QbaPj9V7nSa7RvGr3X3JWmQN9Qvq
RaFG/TsAt3mJHh+U3oO/eh9dVsOxRcVtNXsP0oNpb8kO/WkLSP+wIQak0hseYv3X3dA3o5EjF0y7
c05BLY3YtqfNPddIXHThivqgtjRi8lChhpbNVWwLKqRWTMYtK7B9/Ka7tX/bF2Vtw7h3aca4E+ho
90tdJD1yIu7GOYp22vKc86/2w0DF2+nwGP/64rZPyeezX0a6Aetx0H6AeZkSBvJbAUJAPL6kcjmD
6vZaD2FbreMT1dugTZi65nlQkPOFVhC2TlCsaQHfcKh2uIog03FpVN5aegx84xqtJx+SZMmsfR2F
bGHqreyHbqptZ9/KPHBQ9pERtd0B0c5+9oTt5ZdlVeuwlG9al26svzPT+RmKNbrDOKP07mJ1/0w/
fzDjg5dAXIGglZtiGH2+hv+s4DrBEgQZ18RKnDER1WXN/PydVdlJF7fH8vRhE8jqz3NuQQVfzJek
LLxvRAGIlffY89/C4gOm56MRtmFsmKUUtL/GZX1Mw1XdKm/KXybfmn2oYZFq7l9/WZxymotbTKqT
Yrk7KuIz3+zpTrs9sVkkz6ZREP7QAx72ajridS6bolckFEAK8ILC2N/v9zd853LbAf9gsLrc9c8k
SYGxS59gghKAwQffgzmZv6X1HdbNVNZJCtdO7ol2hfkOdZTPbT4oT+mtaAJerJLX6PawSiRM8znU
s4zmFyCZGI5ItsGt09K/unYv+sAmL6ScPboQmjv4tVn1s/KBvGiFe8MvasVOyuF4B5Wvb8fmzLdf
Iqpvr8Q65O2v1Gcgc06UJVVOJUrX3klbdhtbJ7P/NUYgW0Y5yN7E9R5gWatef+FDiUBHTcw+3bvS
uwV0MIxrl584RUh5xq5ET++wCvgEIOH83x2OOntQ/ruUjlo0FWxySAwJxMTUG9XsGtYaUdtuMRP/
eiy3x3pCkV0kHwmzovL4a6xBsMU1uNlxKGKIBIHAWVgMkiKwyBJQnyGfmA1zYfHYR8rGcz2tceWh
/cIYs53RR06jarE6hlycjv1ffXRsV13Y5tz9vMJvx43VZSTz6rXSgni2gwGwhJT45LKAb8iWwuCV
fUO9lSXB3HPCttIjjebhG9KeRYse/GlQfBM/NIalm8RmApmBBbG8/KDdGi88sgaoLXNW8g97ZhYv
FY8d2aupaIW1G2sb3FQ/+Sw07SrAxY3Lp2yYAYgNeI1kp7an74dKJhDPv/ujRPkE8snz+vbgU57x
rszk7QE8HYefg53riwC90YmzwYn9TeI9vKUuD9Bp7rhl5NtZ+/yqYaI6/5Q/pjMsXRbFAbSzffvT
08lGpeQXxxvLkWYyKWenksAqa91hWLvx0f+/PBwMaN6fsOI4dYwifiESL5SLXKhV6NdDpWqwBph+
lwTHaSUHMEVjk1IlIoDYlsxj97ZPOI7zgAF4XsEDkIWsVR+bNA/OfLMPaleD/q1IcBYKdAt1gtzq
b53K6Z1M9G6eSqOdkfzVeJaKa5qvCKBvv3pNEQIWd229652mxjB6Q+zSYvWNEjgKzi2Pms68lBbp
N06x/OHNeCKAZoTjn3cBgmTpsMHjKI+mJGMBdxvZR+kRfJkBdk/vp+0chkNkzjRAET4fW8mAhPf1
a20AYEPliVXh6jYdK3NDGmm8t0s6F8lHt6q4SwxNBP0x/Wnx2axkiPpgEuU1yFUOlN11vC9KU96M
ShaQ8TjzAFiWHJ9TO+LQ4XqZ9uSKLfXizBInGhfq5CDh0VtjfyAwxDQYCzQe8PuzwkpBztxEW1mi
AuHwrKphyfsax5ycyRUfHEUB52TG9z4iYERUMV4e5LXEvtepPmZhC2UPYU2WjqeBE37MqMDawL3P
8fNSjAmucBrWHx0J6cdEtvzBYV733KTGQHZX0LYFKzKvS0Dj9ZORZ40B79zOuwhHaJ2JebHcfUDg
fq8LxsxpMejtcfNshsmy5PfUPjf5d2hOcdiyfLpSdSf4nwSmSCBSYMBg/gLl0mGtiWc9IAAKy8Gm
nX0i+j6ZHb8f2DcJWCrpseShG5r8Q/nafgaqP9Z0a5JMpYVnpZY3NnyJG4FrfwbvQlJ/mIX9/OSr
r11gWxCs7Y9h6AvHBZlJgqSK6P/jU6Z4cpFTvqJeP0HtGL5gJqxWEEvmBhlNNOC7i34pS38/FwRE
BtI8WufepfDHZmNYC9VT3oPWXv6SSW94YeCSKoWU7EdWPLBKtegTqlgZiYLxfMay1NMSSFuSf/68
2mzIUeO1zm1YlSmgzEwkZe2sELU7PE03ukAOFXHXJWugAPSHcVlB3V2BvWjaEVnWGLnr8+2FUlns
SJbtUQ6Bcupuxb3gY11LT8t1a+TbQsb8mPne/8npQjBdY8AgIURiVA2KpAJsiYeomAFpPW1+JulG
qlgfwR0AaWKVXCxe5/DpKKTmC7optaekUUArhR+gAv8CYlAo/3OWLpIzn+/3dq1whWjDqAgBnsG+
S5tZwwjcThksEldgKmPEVyfiKUP2ql9pD7XJKtyqICZyKExdimWWOkbgTdWacxL/o6YkY0wi4exy
6lF4uWY5gIifuMGT/XOAH+za/owusXcSrdEnYqe5zzvwLwl+KFtoOPAuZLfpc8Lxg/f1Dxgyrbv9
Lwn4MLHwPQKOYM7vMR+7lXSCo1vleU3HNJS80p8M6vKMrgNd3TL+uKt/fIDQ3JHh4nGMa6BtgQdg
KaPYqH+sJa9ctPyC14PuW17r86V4g2i5nDeaHwThcndpNIoocI9qJH8lg7WO9B6Uo6fRxawcbdH6
tGAC6BWj+wRJ+yeyKU5TCfmbywLxEZHH9qc71glMvK8GaYP59IwipEX2NhkpMqG0OjTSeVubwhYm
nA1967mNzpFORm/q0jRDayfTTGRmzNTd3PAHdJVBVhBHxWu9AJXxbUp3tP226tYcW4bP40N4kuS7
tuEq3CMz8BQ6Jh/VoXRiMi4MqwoMwGzy8aPG/Bec7uDJ9DR2HkbwVx7XIjCAUMuXEyyD7+TmMq3r
z3Kv6d+Dnt+xQtqiKkn9bGILAxy8ePN2tojVcrsobo0q96BMHB60mlE4OwvXwTwpdEaYG9lCzU4D
saiVJHYCRTmSeLK9LtMxxrkxaNYZss876qcc+ZZPQMJszsb6iACDT/ODCEsdlZhXHasEG+LOUWyx
qJ2hh/y4/XZdNb3wqFPYmrwdM5jrT3SrYWuPR1WnOEDYktmqnvMeTwy/+kvSWgPwxJOTo0SeoUbu
/2MMSAeD+x3JCzUbje+grl6UPjnooxu0O3AgUO5xrT5i66Mu4K8Ff4YUvFQeZeO8MYf0VzLcV4W1
lB6flHIlcZvVNo/patD+ruJ+zb8EVCCthOc0jt4MrJ04RY+NZFTW4IQSUCdsaPzSV3KMaZwkexLl
ZQRPdmYQt8HIY1t29oFxjGOQ3vcS/ws4at9g5NQKTV2NMDrAmj24+4RXu0Yx/i0y+dvBeofx9RHx
0COMAPr7HxxpBKtXniu2ji0t0mCOX+/4CVuOnb7M6Xg+2tod7ZYX0CNG69zYrlcGE39ppRjdPMFi
1RwO9EHtlhMGXydTJuHqCRl5ZKENb7DB89PbVN8rDxcQDpMRXo9CDToZHD8KLn7aMYokbNJGooyd
lBbd82aDd/FcpXJOKzxHeNHxnFwO6YZKL84CsPXzWtVRoUryAmNmGEypjVBIgdsBPswU7Vw9yTeo
vUOaltS0ToSJdOnArVDxcBGAx+UHQ7OFV21b7zestQ24M3Q42TPTMiHzxluyngoqTwwCJw2WkFjO
RvAUZUyD3HPi1dB/y3cCLyVIiyQG51dIHN8bKfre0YpEvh8Z+9+fSLXYh8pojt3wJ33nooe4vF/J
PWdYVjXNWn7LpkTwB5vrcn5s0tPsxTPBvjIucfCMyaeJp3jiRJOE8rRm9g0yez5Ci+F4pDRJssvo
Ix1fdKo/e/XIR85XLyq9CJomj0ahOphSwyMRp2OYgi62EiPpw6RJCVU/74mSOGaBSEdSwJIMkuA1
tlLgqyGNXBdu8PRl7b0Sg+S6Q+TZplhBrWufLaROKW0af6qAqNmM4tdFaBDb9UCcUxI1GsrH/iFV
zJXSM2gMzQ/n32pTmdoAdQi0D8rqyl6LlRSnrh5T4Y7zm2sP6vCkU1wYeJkmcvYh7GkHtN8aN0ex
lKVNeWWQ7p9Osy24r+GDWJ2/jvTaSkNY5rbCGixx8rfBlYPvb3MPN/m8aLvdCiaW4OwQFSGzYtin
n4mKcHAg9KYMFBhV4h/o0Q2tNQ+ncO8hFSikGk9qtzEc1/6v4/1e/eMvqcggbX+q5CvJR1566SGF
rLHoJddw6nkE87EZVeXzjJNFU9maraFoWC4CK/D2Rga2za0SVry7F+wb278NGYcieOPIkTte9k6j
69AsseVstE/slpbVq+MlF0SgoaQcY1JOCO13D1mw6O6xLI8kgqUpnVmujbhse3pEpKOql/U4Vnk3
VYdX7McIox7gM0EVajthPwI25uGPVHdTpZjS58P0l80wFnECw0y9ABPPBuDWgc8Cq22Q5tC1JwWs
H91yH0dxUKnpqb6Y9i8cbdkUWescHLEq1HTMpwe08Llb0eDUGmOOsVZuX8mJY+oOYRopWRXCl66B
mbkfNEhfw2HiCH+CUb4ol3dp6kvzJbnC2Xh8tRtflze4XeQO/TT/EERPu7V1U7smQOK/v5aG7mZq
rKnDKRPQWJ3EiwRnQRAeA/MjG52TGqEbAeCLkHHQHJ2P6eRBioRlyzBWzDDIaF/EazZBrQHF39Ad
qSBOfaFGzKL75cH8uG1Xho0/I+//kloV+tDkLreaP7Jvw3gs2jYOkdbYO0g6B7xQG4OQJ5dJisvx
ihhzHCDQnnBoJ9GILG8WRX6B+lpkxFkKmOkO6NhHyyWzFKBiCvbkOx8VrOtaCh0C/DnqujdKV9UO
GdiYqB9gDEUUUH4XLatyqX2HSbKBOQnLFsUmZ0zkga2ER6YafZrL8o0uXooXzlz/1GnWsQD2/J+5
kokxROXnGf8N4hFsLxcy2DX2QOaEOEz/NWSw0J//0ftTVnL4JINmXygApxikySHr3NVoJe2dXOGA
KvQFh2GmGTXfbVwlcjNgqYF0YoDYClp3E5lb1T9GaWooFq/9wbbD4gKeHKge+oet2y1M2hYpXlls
6bedkN4WOz0CLo74/+VWJBumRpORA3zP7FIXuXZ9E3gqrbXY5Ib0dk1GrlzpKB5Im4NPXp8WjAxr
nziqAw5pPUA3HwvPvQgz9D6P6T3tnXzhvjtmrww5G7QC8mnbumdVrLh3N+4VtGwO4u4AdfNIN+YM
bQxEuaXIs0TgVR0zfh9NmjiZ91eaCpSxqGlzjsTa5tlwFk1MipRKEocqf5g/CdSyvYAT3zxWV3ML
VLZgizigUOD/67dJc15IelOQSKIwTEqkXJ/751qtXuj/Tzev+fkwEGU2tuel1zDi7MCk3EiwxlS9
8X3Kfgw3sC3brE41s8OBB8LpL2xrczt/zZ31aT3G6UdsSOQaIhjAQ7N6bMvkROC/kbG2qGSJcIHw
qq9TovczqpbRk+C2LjSaRv3Yrnbv9exOepgQMKOOedH/btn0pUJjrHibaWOVe/Oce3zJGDqQCMom
sSnJ3r/j7MGAQ8sBckuDTGLT1Lus8OuzLxaqZItixZ1z8Svqon3SoSd61kzU+0sIOqj/4xoIhXEt
GyXXwcc/tfdExOQE2ztgQnn9tvDvdV+epOv1zN6U4nai46819tErVHQBvtEVrTwYwknBb2jnJOMM
3+s+QFtDK0eODzdX42Ng7fFE9vM9GitK9n8NpaQR16r3kEksA2eze15orRf7tfukmmO/nGTgmscl
yusjXfIAfazGMHVCEJJbfuMSeDW8ek+usQds2xDxCrsuh5G2WYWEUujBLU3uu3/VLyV1IgFtBxBv
Kq69K3cPniebGIzU6vyAxyBxZxWVyy7V3nM0RgkJIe0M85GHJocAt6NEEaIAsDYklKePYxPjon/r
tNLVOoBrUyhkE9GDVKtLT8aFxSxhZnHIaEsyCuGYdCRE6vItMwGi1oE1T4JrJ7SgbchaCbTm7IDu
6EaWb2380Mcoqq91IopfQnSgCbG5zwDTUFjRVfqZxV2h8xblzGkH4XGze2U81qyKnbqzOZ71wJ43
2LxlXBmIxxc2gSMQBLV/rJTfhyGVEIHHgQX5AxmijJSltGTXoDNbVit+DC+xedJHFgKar252z5Ws
DG/v2G532zqVzy5IzhuAcnsK8I7pnEMB7B/N+V3Na1CDIGWkYRlcu6FOJGDG3mcWkvV5dxm7sxL1
g/uvBgT+gCJtU6S8WIQuujVwM/0RXgVyCixUf8B0yK6wrCzO/RwBCgk3txzBmPK+8w9lvSdK/88q
aojrndX7yY38+cIYMRf5ixa+Cu4qUOfUhSkOXQZuCdwFwoC7aD4UAqX0VKOYp4neBJpbV2Yeiyeq
okoB/ynx5FVz497xm9zby9K+tKzGIdhColPUL0JIfqbb5Sv7BKW6d3dMV/Fd6aRxEJMiAPulM8sy
XQvimS4FpmgQms77QCTyN3rOrMzqXn3NVBJXdtE8iCxJwHh7SOwIoz/jmj6Ud3hwl98H2Tx/7Vqx
qoYtmSoh7CQdo3oiypvEwMbtfJ92E9oY7g4lo0R4P0BaglCC/gGoG6izsK+57fbJuxwtgJEniIsE
lCjwnXNF3rYOUMt8cPmKTsz9T3wjhh7G7keBHpkgkYOJ+Hk6T22fD+bPcWm1X1Q8Yi77HSmpPrQF
z3dUwQZ5WfG9X0sfd0XY7s3n5daiELiGjksA42MlLvNyr+iAmEkrDFYFwrkGLhsFD3YSdrPgzP0N
Fb4IO57DZQdwaeHknNsEqkhQjjMWKLs6chpoxLToIPy3ZrvQr3OR1EnUpP6pwJDpkWlQN5KtmQI2
5xAnq4rmwLSLUsNHHhGnpBUsk6jVXZOxYhYSMgNxFEnvKqgQAKgke6tGnblOCWBDlN7iux7NEErA
+5kEOgeASw7T3qd6b8ojTs9+DtPlJTUZ6w/uTePr+9Wjsx1klNlsS+OELNt/JPIiyAUvLTnygGlX
W7dCqjNuZJJpSYoDnn5W4dTIOoI+37trVjmFxt0fueVkqsDdsfVb/gpjSFciJ4yrID5uTGCp3nEJ
cNXBqKMM4GJDOz90Rybsyx8ZO33opSopkRgrgOmGse7HwCuB6iF6kJ//l+rt25hAjP5vgiy42az4
0TTlnpxmx7s6VQD9hkIgA73PJJknUpH+WtomyVv5J1d0pDnwBE0W32+bx9Zr/IQqpzkVwlHqHYs0
ZSZrs+tEQKx871U0TG7iq63K3iXRjF69tYKXLsh+DPQRKeVkXIHlENLXD2rTXZdLRVhCKQr07DaN
Aeyw3kpfmZMJs+HWvNKkIsFVHnF83i1ytundxPANTjQDr/SfLEOYft2oIW3KOdn9t4rG/EEBSCuS
M+qR0EAUq5UCwbGQPGzTZl+fp/OtH0W3TDjXVNleawzvlIKu6XDOC0hC9t2Bj87fgoAImV8pxOdW
6IE4UxnZitMTO22O6R80lvHMYEUeS+ef+QBA+sJ6QS/0ERUagZZRXMlo+JyILBaQbHOVE9frn6MX
1k3gDAptnYqjJRuMIyDjwz9XfU5LyjOa/pj8aKtA763lQCbSPBtCJwx/3lyBMEg1ZbHVJ/bl3+Ss
RMi0x5tv9wnU4KrSmrYygvGj91v60RCTMRHrv3GMdB4Gk6oRzfjULbxdLcBNV/rBEaB5Hz/exual
2m32YDVfj2lBJY/xVNRocoxCx/99BTh4kITKSn6HA6igRkPZLR+6W6Dkfxx/81UnbAUXWulpRnDN
PtH3lEO/WajXNNSLJ16x/g9EqihZ2XkHFes/uJdrtYQWWm/wO4w/gHW8zP1/ECZ3C4o5Qc1TV5Vj
x542CISopQhNk4G0QjssTB9fF2is8UWEau94sfQ4RSbStNJqnjKrlcIeR9qvDRf4XdQ22Fcjbtmm
PcGlvDxohuxQRs+DF3J+k146MsbSowbUMmNvrv+8ELxt/8DOI50p4RrDVDVhqZBZkcCiOZELciXY
ZUS4iJENpJK7Db0X4HldU0ccuk7UZVF+rm0PLxjPq+CpwXoAMRfVecDXrmdPN1Hpe9JVdEeihMb0
ShyuQVCH6v4+ZHni1pMltZeVDY9H1sE2NPtzvUn8NEYWLDMKNPFmgabXIpbzrWCmqqTbwp1+0tqM
1Jvi/cvfy7JhE97mFzXbp1pgNiiRQV9gmjsb6/uvtjL3UDCcC3l9SFl5FUtAEApo7RyGXC8xzkO0
tSwK2/3waH6p0c8j5bF/jdFv3t3SOymZtSLFqhVA+UWcrynj19QOf71sSQ1gxC85A4bfGYVALcF1
fW/NcsBLu61sIqdGuiZRbizrjO9lrp0ouEUxa5MCODl1eIeCZeRvZSoVGZR4xpzwncMhKMsl0YzL
pvzLc89yMG+JA+3n07j+UdiTrWbdb2CtlAI9YQ+/v8dIzvEOepxB00CNwVjZqhmkZWHvv6JTX5WO
DvcEvCpKGY/6a6z7XxW4QcoMvGJox7A67Qcx5x2L2QuUtioMuVZIxPStVehlWVeBN3EXcSx4jboH
5PtO6wgIfobPOy8FBBJ2s9EJ1Ptg6/y2yonX0fw6jb7lz2NuCohRHNHFr4jiSfHYHdlVmD2WPX3Y
hYRrzW/ct+1M//FCkQAXsDCkpPzfwfKg4HA6F9vWkEYPWt1jE/IUlDNThfWfXRXxcM0VYr4elza1
akb039BSzwzQd161eGykFUcyxtfxqjhRseX694Ju+5zbF+dEOR6vv4Ymv8eDS5IyBMSZ9fEa3ZCd
lDIxVAe4IZQtvzcAMeEOQGnCJvcr7Mbn6PSM9Jh0bGqcgO+qO5AlAliuu3bRrObmaqh/5ACPRiCb
5aMvGSpNmdeizcwuWVRBQARMluTuypfrkTRZzxY16wdgGh51ecB9/eadrrIgPWag2CJUQo0GWvyk
aruBRex/HQ29/ER8RFm1n8pTs0fKmwTSTf2NaMM4RdQkwRFrAWv2tWirjwMJPV3fLI7GttmpfQWb
BpUOPnOVi/70sdWJUWAKmxrkwxylAN/44D9WwHsNZp4CgtceNQR/M4BrXa8Dggn2XfLAGrK0r5lF
UhoK6LYvD1Y+5zpuEgomTIciRzwkcCdH0F8Tful6Lia6YwgxKUeM7TIVUkAnHcDNEvkJYrgFQxip
wruioGtwCp5NiM56gsaSQbRNGf28DqsBYcOF6MFQJ+FLG3/8v7ZzK41cm/4I+52uUMKtH/9vs6kO
wqyEK0EM79dFdTXBURKNnN+2oq+WvGSFUjrgvbwVgI6gvWgHf/3HGPQA2D3OHj2FUHPKBzKofI5s
r59BQf9OzC6rB3OwQUG5t6gbjzoxBhWq7tbtfxKap+1HMOtv7oQU3p4vxQGMj41tTx6S/zokeEd3
deX6bpDWy5/cg80mR9dX6e6HnWLLPagAoDsIwf6AKSBhPlB6BggPyKUFL8Fu28KyUBVBoS8bzbJi
MmqsnBfNGL1kS0zC8+mYfuIxNiX8HZBus5Nxf0jIemjhCbYVkS5CuZspZJWsjuAV1Q2yEs4QDMQO
g69rYx0lsZzEao/fTAg6elPtMmldiky6lIS0AsF809UijAxanbLnTr/fv1E7GV+vFkBqDeML9xFv
gj6+0we/29NXkBERYJQpe714JprVPxjY3UL96shj+9iK80dwmMHR2FVEecMGmEKFYH4liAInRQjK
XsRbSZSy/VWMlWk4IjzZ9KhxxKOAaktaVOPwb8SDwR+FfgmHpWcJZHeO4o2xgdACAwdbAYl/egCo
xCUWQjXcVgW1RUbD5GdRoNXc4yBC1AUa9Yf0r28BGYFLK2E4Ze0JQJMr02HETljXtzwOTz4UcdkE
cQRmtg9YSOTNNgBRECXaCmmQV/ImIq+1KegneSxDorltbXCCWjb/v/dVhEscULzWzTGsbaVj2qW4
KflpXv2+1ouNIuBoJgQQ6YSUpcv/dntWynjeA+2J+qWr10dY3mS0SIKyG97ofR5oYFc4tYJANhhl
SW74FO0VNHKrLrqfeb5rS+yWucLsLIyDODazBoLq18nhyk0Hp6N3s1dLj6y5jU5QsR4EbyQ56vUn
HgEgiBAZC+Y5rg5bvPh08TDdvYPpNunjIOh3v43ZpOwBd/3vgFuBvWbxebEg0/oVgPYIWClqXG7m
l/2L8vp+NHXBiDshCCGOO9RoalRnhXJljj/PQWAvAygug1ax8OxKoAKQiQfhzo2IfPdPc2zjKEvf
JcacYC1ycKmc3DpNPFYVz5IfDI5wWKWb1ZhzU1MCYeJHYTQ6jsITLhOOEGS895VM22CZJjKQHJwN
dCQ3O/XsXK1QHlbVzDFJGtphtzxBnTRwQPojQpRmWHMQ75N+8VGnwVxfqY52oPkYzsMiAa59DPkv
+NaJYZ8BPzHfYJkWqRx++XDBHSsxyU3maFZhWJ5qyEfzUjrIbzzJ15jowtZh3QnAx9Mg2LNNz28E
LwymmH6z5p74J8G0fhAeCqTSexxHsFU/Bv/VYJn5Or4ZEWgQj1xOhk93/7g1q2+pMiOvdWv4KeUH
6oM8XFIVK7T4z1U/hhBnHIhEW/Jd+qu9mdUYVKUIPCDstkNYOqRnEi2nRNmTlIRwhg/Z5rXE8d+M
opBBtfnUv7SZbZ4Eh5koZA/ik9YxQeXz5sAGogIDubU1AP0ClagllYCLk1hi5/hqu892+tOmBS28
JFgFHPC3QntyoQieWkC1XAQZjVopud65V+0jt1vsP8nvUCKTGNFCWQGGXKMZN5KOHSa61og9Ztjo
KNqZsGgKoGATEJZIGxP2FMUM9NvllGB2Cp+NmQIcHCXgamKlF3FBpXhjWDB3ZwTspG4VE6e33zgK
cdpJ71xNJADm8Go3SWlRk1Z6buwF8SWh71HTYB3YKGJle6I2ON1jFXZgoTu9tzWvIkVDiXleCpPw
uEeavpuZzoHViiChPVXKTjdPeGGDjhyemhVnv/FJeCr28G9ZQgo0H165Ut0SEsklhqTlraIpLAL2
ze5NgWDVBTPsUltUgO3ssNPwnM0wRcmPbRLe6eTAcL/vcZt1JsEY2LuuzwPN2Av1LgfGC1pZcD+j
0b/ZRclrqxVNXx3P+/7wTw9P0sWoN66k2ZxImKQw5u7G5BI4qBPecKEiKNj3Zmck46DvvBvfv88k
ocl/OzZGPKZRtA4oQGSk39MkIYmHxh4jdGplFgdWaW/krSwocOSAsPAya4P7YqA87mWvbZMmh/et
2F5ZSyMnndOxUVghzB+1TyXZFGTiQ8xRi2cryNQSjQRrjBB13iFFZRHMQB2SWCHab/8esWD4aNKf
htVN0fh4bYDptAfAaMSRdTyi5qouYoxq7DHz9DVcQ9LzFaKuNX2MqBKLg8+v5HIOBSkuNLixvqUq
n/aU49gQCL39G8VYY6yVsDLf4bDTQH1mNVi36wJ/84vx1rb62XYsUcNYZ/Pq6x5DjvlLry8B89OP
kBFUjZisAF21ky+B/QiJcv0RfNWAi9JKlf6gEhJv6Ke8P5NOY5O+5WxuXemLuGo/Mb6+lIAGXo+o
xt3c7cKdIOGqfsmXYgDu5PrO6A0E77fSijH7yCkRL2b9uMe9/OXpcyelEkZwerFzhN2mpSD6d6kR
h6R/wYmxdt3r/QZi0Vq52hiKw0JOczkNPNOoOWugZ2bkwa1gvGFySPMMTi0KGA5xLJLl0AG22cRL
GKuIeg/PIKBTSGKJfkwg1FJIY63Eje3uG2uJBF38zfC1W0t6LFtPGkrX6+7/fBg7TBWBTGIJur/F
drpU7JO6gnpkpBGUg8pUBKYJmZnqDOTUufjysL4t6s/+owgPDjcVJSviKb9X1kckegEGdnev6oOF
+FVXhQsI/0yuCw6O26o6dn1QuvWV+2tXnVIJWrAH5q1OzMRz/2aItQrL4Z5+QZ8IQGFh8uZEVxh6
SjR9HSTVV2zx1u7mzaeE/towQ7ID6v8eL2T7LUR3i5du/YnM2vabO3GrTZxlSagXX+hZuPmdn/Ae
ry6nIBUZRDYurl04TQZ/zSaMSfVF/vuF7YG3CQpxQ09EyYNKk1tBHuTlN2fbTMc3N2p7Ahg/9TOY
mcMUr/1XuvE2CUUtIPZ5Q2/rK5p/yFJcvbPRULCVs8SZRkoRgKaf4h3xCVjvfOHr3/AuK9LD0zDz
1e1CZT1QOV7geRAuglVDGPazP8RabUQC5LVFbXECKRZsCcHpSeRxC8tsz/mOWsa2EXrVu+Se/f2W
oPYbblxgD4d0JNjyRXU99iOVFjI7MW4l/BL1YUvsrQLn3BlTFQaTEji7w1Ixfwugzky0MXHNKUwc
lnT+JKQqb0Xl3SRpFw4DMfVWJT1Pa+Eyzk1GtO+JetAOsCUzd33gnLPRB8VUL2UOtbhr40qoKeZX
tbtBNFYj/zMP3MtlKSceR1WD27uLEW/rmHmh5lLe29JlqxaXUNqNe+x4Hl7oqoMc9Pv2AM04qmcV
OhrhOc88n3+81JyvqkSjco93zp0TBp2vYr/qon3aYk6B+qKh/HfO9GeztSP+gO3sUGxAW/eOXCqy
/uYzPqRhbP1VGWCaXPUlsjuXc0glz581i2juUB7qN5GOQVdos600MNRy/+uf62w0oW+na2JYy3T3
YoYzcy94VdErH/hMNXv8ziuTyasWgEb4GQOlGU6Aq6jgzwzNVgvSxYnoSGDGyQS29atgCPFtNoiG
uycKSS8snm+mMTzEs+S7eiGnk4N7Cijk+mfQjdAiGCDZv8lsekbHQY3wRAIfDnc41gQQp0j9HpLJ
hPJ8p636gHBjlxP8nU5P9ZzyGKD52/SCr6f+EcbMMNJ3F59VpnGjcoEaBrcvZzhui4fodebbvuY7
yh4oMHRZowQdXS4xTIsV2tsIiaFtnyZrMHt9780A45FvH6Jpy4kMpzE550IF/yUdn8AQ0O7ftUqi
RjiHrvNtJWBX9xKpq215JV2QnrcyAHhh29pJXQ6WTYVtsXG3fYr0+FffIU2rJrGevaOFqWggryGU
SLjOpZZ+5iz6uqnsHNSq4Ri9SXm8YHCnljx+l/zDDZgy0ivzpUeaeOpUvuwOQbzja0FptMD4ipYZ
NPsQQXBfajTpBukO2BwtLrKsgZ4ABq/MmRYNPhII5GLWaodIs0ND+MAvSRoc4uEG5CXrdbIa1A3W
AAQ98No5840cvTuszDKfywuh7OKYaSZcFuLFXQ5al75hJJK+nBuWAHU2NRYt+5mSBroy9+kinRk2
latvYdm2vGxm0gEg90kiB8I0Br6i2eZVpwR397LKk9xK+Yt44VABYvniR6/fD7yfn31dN1KmR+Ec
eyoBjAI/IEbYmjdzudusDWZDP+bB5DHkSDMfYorZDk7nRIgnP0C1r2kLczOTANGZDGT9QO+KNam4
TLbaV7qhfRhA67DT3bqAnDAiv+baMXgyNy8q52JKqRNXs8njB9dV0AYCcVO1IrbYpsJQYNCxYk7o
BZTnGm/vFjhoIdbQnILEoyhNO/wJGmWdgclf+zA/gwQxhIzdSq3oFvPKmhroitft8cEZaPVnHq20
YPVzrsqWektNs8/WufcS5j50iBwyaGJLmPDRqEoX5AoiBCwOwcTHJeSSDDD6534qzgE4TG5rtU5S
fEUxm071E3L0NOhQdQrbKrJxgiJGwGj4yyFzfOUFmy1uX8eAQgp03nwIVkxhCHun+SFKhFYCKG0u
u2CK8ChczB4EWoyZyg7V9YjhMOYu1vYRAqLUhINE/UHGNs49JvmVmdYgwybpREdzY2rpSQQ8Rorf
YS3DuzvUPB+sMXzYau2iklcyCNTh64Qo6rjVwvEOK2/dYbfOcmkem1+TUM1pAWNtzqQ7+kIrJ6it
egUHFbogC2+BC8FvCsDirwP1+gLXtfI4MFqvs1SQtX5ZFseW1WbOv+aa9hAxZbNEXctqaeBC1TwT
PPSwwcyqwc/4XIrr+1BfUHC2kp6CB6mpG8ce5JPgDJLI8o1mK7bhBhRcCFNdOTzZixsvkeE12TQJ
xtt1T6GuYoWMMBdpfpHPUHy1Tla+av2REmP1DFSw1ct7N21LM+xZURU2SSYbFInp5OwHDclsH9lT
hpJE47V83IfGOQg3fnyOsyBKMKyY8PpXA0ACYoUsF+iHyk+46LZ219rjsd29tz3jcFaqUvmTExLA
j0+IcNMQbRo/CqJrRRgd2Q1rCjrS3PZnQ1/H7mQpE29gnRsRnpdw0091B8m0koKm9ck/GdgSJGG7
FuqlG8+szduaJ175xcWuQFONVs4SVihEI6ezjc8EZ+2+swV5Ntka4XOo8frzuKRSOMgOfS472WAm
asnU+F7rkSJ5ZEuvQ9Az6PUN/9ry568vCGtoeu+vgCTky4ULeZWFx+nrWn9o3ixhlVEqcIzQBE2X
VqNEqdUx5Le4gq+jsxpRPdgc4gERhg3k5vZ080vPiUHYRedPnWxX3FaofasvFS74zwHDBv6I9nl3
jRgH12+CVtkHcJLH3Y7jC9zcuSGCWe0bGLIiON2GtWe4c3y7kthkDjHwyGGDn0iguxvFzmhem8zy
U102Se6H5QEFt98oCjfg6WSwz5NH0NixRI0UsxpQZLTErRmwTHfyN0s14rZvrxHTvlOYKd8iQP9X
se8QpBPHN7eN4GSEQ+gGlKGxC7UrCiktqG0jGnE3uTDbXoqHimiIflC5GnCeBtLsWzhNV8L26oBg
zovMvx7Vog/DPy53cRIV1XGXAfijS3t87RxK3EY975dd1Jm1jrYZgPf4sHPu1SMToKwqqtTUgBPR
wF7SegA8c/f19lsvRNVUEbcidPf+Litr38uTPC4DbdGSHbk/DF5BCJ+O3tl4Zohzj0JT+MRfX07i
BD3PR7D69I2dRygaQBs5qOi7yf9YkBOmOSUHUnLkhh+7L8ML7E7cbK6e96FE8AVJ1FQHRwOTVcKP
IhH5SGtzcNych1j1Tq006xsNX8Cflcfx+6AVvaEdtU8EmKPvIt+QI0OzsEEhMFWyux+WfM/ucFNZ
/VYonL5seIkfAJ4cfrhc1bObol5Vzh7fw1+IRwVrMuTy1PwgoT9Sbi9pNSn/s3Lnbgx666TemvoA
pjKXyag+oFxaKefWD9jU6MIJBpojsNaVHlCqa1ujkLd12xRz/cSvwKD45Q7x9kMLshJNDtqqT6GM
AWm/ulGt/5pjlvdmZTdCHqBT1NwPe9cov2N7fQ7dTCJyTYHSn0RG2YcGuohHN3i3ucHW4eY8pLFt
R5a7ipKBCPSvMzrbPSf/IJprcr8bVsVoz+1JHYiZDxnvBx+M5JdoTur5nTK6yd9ZQYjWHakvRHmA
Smtgu+iMLd/AFxfcQ5fxCpdc9AWGSLLGsTrs9MduwP6obpD8V//tTiEWl5rg274YUAsQI/z87TXB
RhWH0pEBSqqQO8dz+E4bbn3q0aJnvdSGAUVXlQJOaoaZ+/iEjb5v6/TSAe/k2ydV5a7uwh28QZcc
BuXvudEx7SOlY/Ak664m5ZpfT6FFERge4Q1uZay/pWih9HdrXLOFaC+0jakij/omEEqje6cpwV3U
dlyqq/TrlTFS4YVIixN1AD28OMM0VedAvKFLRO9qcatxTl7zJ0JDYzF5PcXHqF6n7vVuIexPmiOP
7SoHRLVHLzeVeuPgSetgfBitGauj2oCSqkL9E6MxXxWvZy+6EBZRHC+GbU01N90PLIhW3vg7qpJt
e5j0t/0+ONbDI5TSPvUHZ9AO6Us85OTY7qxD4JeHfUs6otioTF5wL+ejGaXbgaeczj8UbyaJDCtn
b5vPB1p3qdPl/Bqu1m/AJFC0UzhcdEGNe8RKbCTrqPOEdroNLiYJUfO0Viu5Xmek1CXuelvLfbF3
D7BvWWLu0Z6JEqvBMV/0PMv3Cw4WlJYz7D+42nALgk0hSzbrCm7HJHmnl+FteDqkFdKME+KOJerD
sWqYxWZJ5jEyRBoSeTzODiW44njO0Vp1vjNOs6bck2lWvi2JkXa6cMJUK+FRoPO/xUI/aSd5u0dP
y/uEPaYHDls9/fPmNJZcAvNtUaO5BB4gjsac0UVmpn8zOwtliBI0rNqHVSennU4TlwkcjESY+D42
piJYz1Vsk1Jw7Qk4eUpURoF/nMjaUsqV6cGcUU0dA03JVtzz4Q5pRJhov8y7fqciAr530u/NaBrN
ruAzy84yDrHIE58/dZR53pTkI6U69bGEx3Ut88Yc3gBVG0/EFYpEKawdrXVAugujyKs+e1gOwXVd
wXIkJbjp4wcIW5RKPGZVARK8CYj5kmYcS5Knjsf6K0xGnU7ji/w7JhRtiansWfppj8wrH/vfcy8x
CpNJ/0EsdXMCYOqEnVFoM6Ns0rRR6FNBGVbC5Ojvpu8x8H/50MphMBD8ac/1JtZpnkVVXz5WHTPD
GIOg4aMFP0n9XXNW4i/SvzKR5iSdd0IH4xE2roxXvpqUDb7KudNGQlLs6AomjfVIeBq3Me7i2Md8
N/cxshuIHYoqloydgze4VdmfFJUsDURgGA7rV0riHsoxPFafFvLyy6vKJUgaWwoqui9aKJXSAOfJ
fE5/ccin24bc24t+c5iw0MRmVa1Tblycis0spPzkNdAuaztmIF6+NPbJsFHx7g/MV1W24KbESpZT
ezUeUnGdXVhDWNx0QUun1/GgVofkFelZZgtyTAId2R8r9Pt228L1VPCfrA8SlOb/x6zTC3ltxXb0
oCAMnN2LqXjx+oM8qPwBZfKw0DRlgBT992j6LVL8Mp/05ca6N6UxCCuZAjLdcDYzyf9m/CcQZMcc
SnRfq6F8GION88OqtmljFALwTDkhBU+EZO7OevSe7O6BXAVfRjUOSPUmjrIAu1U+Z7s/GAhxYpfT
tDokhtARSRqMt0vVBxFCSWJaba7+9OshDTGZVtr4ZqRCkkoN0QAv1zsTlft9WqKhSGsYAvIfc3Hr
UU61+Q3QRkEyZEHHYIE+FbxF40Txujs4RherFykk31w1ynUXSuq20/BIBk06Fm0I+2sXvSS5IR3X
moS3OYV5ti69Yv88axnj2pFsRt60wkAzlt0oY1P/NbeYkWhN52d6dsx87qrNQ8uIv51NDQy7xYKe
oREPOzLRYyVovoH8fmdwydxS+rnfOGn7NM+GnWO/ztZpzRf/uBS7tErXrTAK0GA13h/9kCUIuinR
aRYYNefYQSp1WUOhwJvyhAlYRHnaXThAo/vyZJ9sJsk4sWyzGWej25pUJSv1jdzFBHJHxv+64ca9
UKYZ96Uxtos7d7cy/73Ej5je7O76V95ebPER4HDT0A1dDBExwE7SV9aQgGBCKPxWsLwzCnfKjQyx
1DErtd7ooQ5ahJvgCobr+pp9piFJcm4e0LUqRyATFMku5A0zc4qizfFomZkFyW+a0JxFnLMm2KHA
1Tvw8elnXEjl9vlykOpXU3eVHzzQ/Khq8HH8lOgnjQtdAwAZ5Tb2a5wbP/vkTnXDlCmfhZ36SwyC
WSnYI496RC9kRgMvFAlO6HmKlvzTLFRbUEUnXcBScNttL7+czD2fsY2M2C7nZzcapLv09ssBvuw0
cTbnLLGAMdmXiRXMPOT1kjnAO+2BwOnePscZYUr9gEbIUpEcF/Xzru6U9A7Ssl1wm8Cx0dIprnQk
hOfvbYHUzKFDxBGqXHlFguL9wL8xTm70gmj0TlxJETNXeaYBc+asgt9s8mWqNFqEvZxQ1IvGZqEI
YZKwVyK8QfuVozAcVGMqnGv3ucGFzgd5teUupXsbPEE2lGzPIehPAvUr/KN+n9VvM3IGFULEltQA
UgdRPlS2y5RDviHFj8+nyygnzUK3lzI2WUQrynTy4ISdb+nfW2YY3fGwFXPeibKGH7EgBd7tuuhZ
wF184DEDa+JKtP2ubhMCHYWpaZn4foTm8qeTNLDZEE/Hg3OAmOUKK3UAw9pLReYogrKoJ/GH2exp
zRwXGDchDvZeyPkUEAV3Ym4Soh+L5ZrRTcQmnTZb4lzVjIJympGasWzLjC1TJNFQ5hcD1sTrTCxd
lnk+Sqqx+T3Di1eS6hbY1IIWGFW9n9yzDREAc4wHzD7MxvjVlVLMPa5u49Jw9sdzYic7mGVGRKnu
XF1/8EiPIAu1tznUvy5QL6I0Ly+iypStyzV+wG8rPAVEdXJgCe3i4gReNPueqClZBhby+PCn3iqe
584YDEbmcG6NXRF1TTetawjp18lkWG8wkN2KUq2TZV5ugg5cyPUgrSK+TL22JFMILtdxF/9q7ZqV
WBB9R0ykfz8mXsK6n2Te6iM8gVPFilkkcfH3eFIZdXRwOC9L3jx7TRvn7cYYb0wFkAEKTkFVDXUc
COegeHH0Yz4NCFCJZFM1MB1VUyAJgCoAjrICnRULVdqNs5e/IQOwDvlU4f0Rz6cNpIDY9Ruyda0v
T0RtcxPgo7q0in4ja2RRQQkEjTnMVgKxB3Y/WtLCKHX5nSDIkOIhO/3HtsfQzGFDqD4OOmuevq7F
rwTHIS5eIpITquxV+raK7PnELggiNRM2DxcsySp6oFLzIGPkwm2j1+YDIkZ6sV7efHJZ+auvWUv9
hf8D2VakZ5+f29AlhXq49JRbPeQ8QDkz0U5lhlZ9cIKJorDl0OpymnuLbvq4QYuA323ojNAwriOO
xH1usMOyIELdBYng5DP2klgO45E598+ZhLL9KMpUkYm3lBCn+V6B9c0Aq/TQVh8wRfQ0eOmylDtK
3KuXZxMp5iHhq4wXJi14gpcefguF/r7t2TvbcGr9hQpJH8cfTqzUbr79O/Q6wQW+IdUuGg62bu87
f/N017RKS7+VqTbRKvmtAcjU6gKgFBQgirjPMMUk+z7ZjFwLC7wn5B/AcP0ZPtm7RR0HSvz+luxp
RGjJci03oMbiSSKLSsfPkpSD1wQiuOfCnCwsJTWUxaIIXM9/0NOaME/CtO3kFBZGdNML9nzGDYDE
hFWz8uJ6gdgSnhPWuB+Oz6FtCAyQ8LAH+/5N1y7QFY4VCVWFRjKT76LeXdkrTTU+XSqPTID3JWP+
alnLziWnqB4FGrc/YfaKv0U39ZGzNphJ/qm4tLYZxVuVVEpx4o2hxRsZE9OmOzmFUGj8UG7cSASM
cTBn7A4qPBTPACBfwDphvBMN7LORI6XdLjIBZKgTK8z2Y620uQhrNz6b2QyOY6G9FTnB+m4nQXhM
tdE7ZYdfv36xhhQ5X0995Fpa/AruiwJbZfP04Xv3MqT0o9d27x+D+xiGhug1tSIMToVJJy0qd9eB
rvAmX1tC/atS94kWqytECsXDYGu2WbDjL7XQ5JVaF0iDpAyicSOi/VJqZ7+aY0msKNOAiyAo+uM2
ubceT9wDgChtBUVnhqlJJ01L7LdMjhX6swIGoNb+QtyozilEDKBwPDCP4G10nHsdBcYv47kEwsYC
jCEtvRIW5y4ev9q9735Sb68deoeyBOMgIMfQaJtns8lucsDWKO4hqlGMXdzUSBW5swpqoiwnOdkO
iMo4BwhtTAqczX+jU44T+df5MRTQo4hyDCgl0Nf2P17ORYbamSB40LcQ4DDs3MGbjE36XV3fzJwV
jGDYYqGiUceF93a0odCXoYnvQYSGdfmoQyeENDPnxjp+jA3jcXVCHlwmf/5e8dOoC/WQSSz63TpF
tJ6nWd2/DIBTtChCvAWmInXCEWuuaqfFyBMX6R6iKrTUtbbDt6DIcDy30xtrIK7rGwIBaA9K+8t0
auaNZb+mb2NoCW4Ygx+1UPnxDkBm1l5rgH8n24Y0l7XhXjC1h+1T4EebBFyQmLG1xDQR9Ee9AisC
xmCl1G91TCskNKTG1Bbe//fDRsHlHwFTG2FVZmZK7kFFPHbNl7IUBrZE0POpPrQbbL2Uu/5RQ3S5
SPqVXOYX2cwRRJSPQgGM2l5g+FvRs2G+6HJxmNLjLZsrvDEV6IZxELRgGweJIBZlVabvSHYYeoXm
/zSJd0OMu4RycrKSlSlLJsYMm7g0vxUTq1UcZwoXXFpmzhtVSYfse/TRR981H1sZ/jncMGYfCNgv
6iqEfPJ9UWYoV1oGlx1tjB5TnGOWsw8vLFCnqRzA3bbQ5eyftqScsnQ82UMmeKc8ey0G6kaiU4g+
hJ5G88b7iYik/YfuPGiNAMukQbQ4rOW/OVnk9M38R3smFrl1XbFXVcnqvncLwtAOegWuIZDOhEMv
MS0lmmTeuTvFPoh3uS154HMTDUKAnIgU26hluWg9s6nUnAQlUfZpMLGHdsrrIM+1Yf4FVncN2A6o
jlMYiWC8dOti3Ey12U3I1yrvuE8lImP1jGBOkGFEzIRjsJc0ypkNvwP7FUOxbeennMaKmHcUF1E9
vtp10XUVzNV9PFoiGc32FzyLzZC6vZc9gQR4nwKJ57ds50AUQIAWnF54H6jIm1FD9O2HKOhMy+AZ
m+0sjAWpW6FZfpaOMV31AjC80H8zQRq/9OEf3iEm1QyAe0Vtw714bJtUYl5Z7zNhtb6mbb0N/P2H
7SV3TSd4NSorovTyfOyqqRqN3wd8ZrQlI1aFe01JdzPoor2WoftOp8pRioAUZFCNS7XsWOkOUkAI
rgyabXNsuAaCG3xmTvRbM19c9xlMbtJ8n0nKs27K5+mEEtrZB4q8FUsauL6n1DnTi3R9KrGheRXo
4fXJvqg4cQ7RwQlHxEVMR+jaMHvueykRcybGNVWUyyiQVOjIlOssqXxArch7eA1goBrj05OMZxRL
9Eh40zjEQlYtmDHWDog5NxB+GFB1V3CgfVYkAnSnPDH5gQD2zXcXB6EwD4qqrI/qTgRNQXRJEDh0
4TeSpjulH3Tcmhmrw8RjeythFptGgBhAPM1cYDiNpWcUOXYyToUupKQHpaG6y3ZcSpGMebbUrzfz
0SoZxXwBBXPT7Ps0HRzkPHjt/2QpPspBczDHMPnxSThSafQtuyw+AvL9qhe9Jjw84yDhmlMy7iF2
ma1wjrOdvaz70Ya3iFrUcm6wzJdZeHbp10sgI7kXcSDVQjplUcHBlK5RbIr+eDadtc5E3bKRBHgP
SXpntQxxZUzzMso6r3f30fNfeB3rpV4PE/WbWIGmdsGEdVH3gTGY+NJaJ0MQAfBQpDeYlfgJBZvi
0rB2yXxhgNfyZPFkvLm42lWZWhuv87CE3IJB6hDUkwjtxQWVRbeMVP41aWTQdhocuZbzxRrc5QGR
5QG86APcp+vKsc0oec2S+butweYZ9g8D9sVf2KTltVlY+HSjc+k409krOLGEOe8kHw3vO197q2en
JBMAHcDwzenwRHhzy4YadTIRvU8WW5zE00soKldpe0HWrPfhgz8jmuWtJaU73R9wdwc2Gh5/nTSJ
8vI3f7C7KjKGYIOWgHtgkBa3jiP8j8jg3fVJz82x4BCcz4y47m5Bz1DOqh5qdvcufrAQm/rluLk0
MG3KaVnCbCEs+bQ+OI+/qHaT8fDFWxKsTU00PhUrohlVB3bw6vcOGO47dlC5X6cbtDQejVckinaF
AsOPzjGgmSZJF39c9Ju/Sau0DwUg4KeA7+YAMvOw8tiNX2tvAb5mRXbDCmnlRyMGPjG92vzEOGcs
+yrX+ag46XZjkoEELTi0xfATR3DfhZRJHmi/FlaGgoB2rlZk68EQ+MZliHaKULSrVCBHojFt0oP3
iryWscYEQIGp5c7gcBzwU0EQvuNDDZSL5aL5T1Ag/ejL5vjPcbQvEEwhwy5pLn+N00I6S8mIMlqt
Zq0PiLtlS45tbRNcBNhGajUjlL+eCnnv87N2R2qQ0J+HbPGilqKgQP0dNN7zA3bDXOWPseQt4a8S
uiwECZgKqL7UyfIx8mF8ye7X7dLrbVaiPvOk4vzO5j020rc8Fre3dOoU9lODM900QQiXfDrlFFH2
D7RILHQVHB5pMEsQqyiAfxwJBCUD14T/2bulCKkzoyEgnthWeG7UwydgyUtlX+/u6lhehbvXz+dw
2sDUGg94BmVf5WLHqeEALamOE7FdMaqSLzUTFVoJmECJGbttt3ewTm4wjMf2LWd60tVyH3xJ9lZM
wqrqn6K1nAJcP6BslelgRFmX1gnwI8oUUBslYlwiRaHwh+0EfLNDLHgikYqZQC85Uc+f3hcCo9WM
HJwR/iytillClzEEwp/qSUK/9lOB9v/Myw7MIHp011ceIzkBfkDgPOndc/G+Z87vP8RKVu35dOgF
26bLkmTCJqolAayLjoDgIrVjEbwGf2FckwRYBtQaDEWJdnbscbDAnO7SoD6dVlwUtGgNlPbLZUiY
ICkRxdj24x0hOGB7Ra/j76ZQF5NHVD/NTEXu0Y8HTHtAVu7siOBVqRn6fcjR7YH+rahtLKLmW/1g
R9fABHD+UlWr0Fekn8d8CDYO8PMjobzkSt4jzRpdwlZiuSCWAIHwRjuMOvvWo9bdDC/15WR9pcTz
+UF3Ci/HzZRPC5xUvIiuGHMrREirf07ClilayYAucrKZ6JAgjDWzDhCD7PkMLNG9HwtyebboYI9U
g8lSBxvLhSdrgistInhMtT8R1MfsPmyUzJPayoWdpsQ46YIVUYTZ3xNx9LfBB13eIolG993zpEaf
xGn12hAEpWsbNWB/gWbaQOerRQWfzcGafCPUOfUKSvsTItuhJ4bPUY8MmgYqVRacv0iDnwBjM8Ug
z5JXVyC732h2PxlW2hQFDMT0KXblBsYifWKhSgTWTVB9oFk1cTuPKsu+77n3P0f0vW5A40oAnMgy
7Y30PskZstFyCN/aEeFnJxpBAm0AmnigRDUktCG9jkIFzCBT/yrbmJKDG1d58TTDEovmRYj/U1+7
df+60TQlLE0X0oKby1IL4TTxNvQigqeESOmkHyWj2zGejBPlDF6UDfqti5x2Z+uuW/7WGnQXD3U0
+bPXsELSm4xGrpaWMa46splTvteek5eclVIYE3lHecIbs20VuEYjPpYr3ANIBr0w9p4IN9Hium7s
4D6/irlVzMJ6rbOID/RoE3IxIzuPjcJsPwwtJPWadwZi0Nx9SlM1R5ERRJjgt/HPw0UGp9ke3bBe
vfgwjG65H14MzxnDuluUuWYHPYLXc3TgGm003dEoPLjtHJ55aQJ2T2BetCwjh+pjzzJGti1RTuBW
6MW3dgR2RFnH5X3Bhr9Vneo7qh4ni/uqJTYv6b7PPerBhTjWeyutOc+Ea6P3nyJMwv/4D7OXu21Z
gNbhJY9MBDIROmZL0F3p2tfTrE+CVl/YNR0Rsbkfr9dTTtgydSNvGQQtbkP/U1cPSRgmyqtNpGRE
7G9lEDONijwI5PNzVmclyR8Pww78y/mVHpeqyXrMO4hoE0vphcJFpnZKV1n5umoPy+maKUrrKD+S
R2YqP2/6AZDkfCPl8ivOxDlwq+KxABhVMsumfOVmNZuHrVPAHmnQr27WTGD6ZRl+ZHdh+VHqvtUE
dfrABqqvgjKbTYaOgcLLF5huu+SQTyUD969NYd3SDsh1QtGNj01U9FXwkGV20zEAfSClW3/feC1R
EW9ZLZ9HqClhChpX0WPdmclxxOVPBs2DFHgf5CrV78s1BkMG4oCCvYJj6D9nStYnXZWUwtNqy7kk
23mMFVc2+hzY9ti/SNiPjPTMFH2ytwm/CEkN9gdK0rJ80wg9MlMY6KBa79IeOQkxJyukJ+s6m4e3
Tz43XX6G5uN0nM6Rv9YTWuNlIv0wrb0gT8rT17xyARcLIg40l795xLWhxkzUqWopVjcqlfMXkSLg
pFkBQjXbh0wwxBwe6PVrBEFXz8JzHZ2pnehXgFuWBVAEIU21kwAGQufOwI9nNCIkGKktO3YfXrJa
kraoopAzG8YasbSdMiYX8PRZBqoq1YrqsAzErSwMCTpvc/iFAEoTxRU1W+IgZX/N0ClsKBOXAd6K
ysurtvN3XA5zBth/O5118WzMGq9T96vXX8dYmrEHZ6cdt8s4HrP1/Yut2eDb/CdzBr3k99pdKGH2
fdDX1FpOPP5Z1r1Ly7ZTDCG4TISWC3wbZYYD04YJFgjkl/caf4fsRq6ycF5yzjWXHO1zjUkfCa0e
0shZICgnsLkzGMtCkSl5Lz2DEs1f/OWL+vL3RKZFfPjklG7khhQMGosiu6wdBqxNHOzgacXWZ4bI
gvfrZX4saPd4Q+AdNzJARZGMNEvE7pbGS5d5gpGZoozJwNb8dHaT+fazLlwxvyeELeBGSJftspvZ
oaA+z9AvD6IqTF9YFweIwbXOgVWaltOGqbKcCZ3ncjan2vMIUWIrnOZl0AVBIR1yrjD1cMsSKPOu
43anWFjLgcJp+rgYbBiZXe3Uh1ZYbvJeQioCzK1gEKTJqnFbshkrYDxqPeRE/X0yWqTrwGwvdKb0
JBZRKuNaBsAiKB/VtpDMv3fyeMp7JGL1BygqvHxSL5LIiRb2fJv4d99ivGfEdwUvvhIM9xIpdQD9
e7pjcQamL+VxUnAWEGIr2bQAZNL1ORQqCfhUSgOtKzFrrDIuyGXgfjMPiZVmeqO8G43nHVm6o5nd
05HGR9wRpe8590LIhq2tgonIDbrK9qBI0jR3hfeuwroKZN4aQuGPgr74wIRpdMDKGGpRZusiC9GQ
tJ3rZCM1gwEHFFtI3q8hI+wcAHMchP5sVfVwNXPDRJPky4lda5mN7RqxeP40ch/t8PVsr0zs/kYx
xReP54oV2p5OAcMiSQ9Vy/BE6GMfv9Y8f6R8dcbiJdeUlVEEoMRkryGy7Z0BnzQzbFQDN77THy4+
ISMMODOcefeoI/3Ja4zncj3Es2Jw0ZvD5GyJEta/ifLaMcxqJ8UvQ05zwVkIWe7OWfPBnEFrPYIx
/DqkIONoTCs0u+F3tSORvPsy43MZobTqi4cT7qWsK0a86We1WWnChYpRHb3iRJEYhuKdG/gawNtS
tzfh1XuedzkZErSbG7xfu9eX0LdSUtxDnPRUrQTqyIZ0THylDA+0cuwPG1elvxzkHqSEG1MSWVU1
asuYNqikVuy4W42PPXc/OpjaYubG+yno1ObUrZSMd/hkPLBYodBcOX8hhKyIFYsmI1jnKpCznCSp
xqDXKtmq6EzYMkQ47WDkC9835ib4UKzfw6M5zI9RAfdrAilWt9rMQmzIHO/II2pD5qswLLw1XZdc
YXAfUdXoSkA4qKqjfyOA88na3Vaj99WSDBz1XDC58xo3qTicslOeksooeSw37Ysl7yP4oQVMGy1p
McuRAjtZLc3c0dnF3CIVOQH85dGxAM2xEOn1q5lGj9P54ZVoFscdCFo+IxcNPYWqMRqsRs8nUtKZ
/j+166LXiGjRvOv/R7R1O1lEJQCX57jRisxR8u6uY3TLBjroinVPSl9eYykww0qe/s3mmK91iDwr
aC/w47gf/0a0+dJiLYqOCFcIMBF90x3QFosCTZ+kyHf41OS8Wfu7LirUTUb+MXWTB81FvlCI1rNM
V0oMapC3p6xCdZMTbCj5AP41eYrQ49xDvc2j0FCPjLfk1zTSGNolYtC2yEFBoYzqt2KPRg+QUKFy
N3zVUbpq54nk8G7cRlty6r627+F1FoINt/9vIlQ/K/rnih/byrnzKa+sOZgDog060sZDa5fG+MI2
eJjV5Njdl1xBbSjMnDz3Zs/TAZmAoBaizT23OGk5hT2/26POhKy2yjnjN3sjHIzwmKs26y2Y8w1t
ORH0EXDfT8OrN7hfGGAHY8gJU1EiYddgSjnbs+a55ypAwH2UsWwIvWUMmYRetdDhEba7xeXbLug6
pIdFpCT+rBk43hg+CyNxhHEtZYRz8q1QUlT86XAdiILBnlwW8Te81dA/av+0U4xD4/cOZgFNj4rb
FBPzKb2YcZ7hD/jCRRTGndW0wBv0dyuGeCjV1WhZUktXMLxasTofqoI5dBzmJaKRL8nnIvatQLr4
leXM6ClzsIF6IapBHgVOWhQIDmvam9yFbs7EFsonHj2A0AoNSKo7ONRpeZyJ2hZr8+usF6WsJcTa
LdHPk56BiOsU0P1lWT5MOLsdyCCMIIRcLSEs2k99b/8s+sO9WRl5jz1W/I5BH0g9QIQrF8nbvN3l
Do0YNvH2TbhvI6LYpI1wVU1CufgyjJzCs3+8yTK9lTK6MtqA0HSYmr0BFGlXskNfYm0sHp2mrB3R
IR9n5oCHFwg+xOw1ztgev/B2MhzngZpwa2yBz3bQdtjuLKlmeaLfLBS7quCMwOkxa417jlZenHCk
yrwVevJsh7e8/rmJPnkGdvCvOcYJW6ebttC7N4D/dTmkDXc5rmdWYlNaMii09aRQgNx+2lO6rMzh
IIVCnTMs+cITcUX0SYG/cj/QXPd/Psyu2D/qxqLEWBS2i0aQXEorWZjtbThOOelpbkgYYuvobhnW
7VK24OrzgDUGwZuCnqyB0twE0YppzCY5ciIK7LvIeCcDpoNgPit//Ws3gL9p9OTcD7fMzeHl7EiK
XOHzZ+ssZDudSvDlXrvzzXfMi6DAe47lvl2pf4SAjA00c0ZWlVk6TrxNwFlmNuOplhK/qYsr4O2i
3SA99jYToPXhJS2IT/E18lxa70/LJ7b9Q66Uws07uH5Nw6XPRXkbkzeLSWIyrPByonbz4uyscPDK
3kO9001juOsFFDM2I5fngmFvVUlAB1kCxE8/Onz7IwuK6T489Jx9SJRurbr6TBiBmi52PeXAPjHs
Mn+LojLOsDlzaGkn2QHwWvCz+z9iuUfd2mbhevX6O5sNITel3wp3pIPK6S6C7s7GhmiGXESCCdwQ
GdJgFSRgpv3vh32L5EDRc/yqwJy6Qz3vvtC7084jOHnHWmc1gH8B8K9Q/Wn4SdgVgRDri3jyUmDP
zn5mLgUvsyypX5S8XhPJLKvBHeo7cq5icsGzLYJwblfu9CtvLNm9Gn+U5zQ6QCWmkQIjoPwL3IY6
BrQIh6mOfxUj9+/U5RqgVx2/fA/eL1Ubfw2GuX30/MPmfZoYBYRcq85FDiAWGXzjuVtqouQyEINf
QRHVDIUZvLOPgMbva71Ywidgky0E4xnew7zaGP7rTDvFfLbTVMkScky9ci1FEm0gJwDfqO40RSrR
YVRc+I2JcPWkvZTZr07iWb2lwzLM1leqETLUIm6/SJwerlzCUza1HXkvNsOHtmB8ukpojaG8FLKi
At9liiGMuLeMb7eBrKpKDN8Daiix4O51oVlPtuFHbbeWeGGkXGxYuV7+TY99L6OyhVpLX/d1oNnb
Pv9kpOHeNrBxk0MXzdnu52d8nXtwj40uEVmdkiYIfhkqzvTW6SBCYtxIftx98liRVN+z/GERNRxX
fEmd52pxN9idsEldO1JLupAZETKl+HEOFzvbAKev/pfDzU/Z3skkY8CDnhnQ80FRgcQfaag2NlZA
nacePuOOTXreVVK62kO3PiITuEbR14J8MDrM4cTQe7048oocosJq5SgFvSvm94cpbxkmpl29mtk7
shHxXc28/rYTkVHKLEKJd1KJrUEVrP85CMxNTV7vZCALm+R/fY3xhUklHaRI77ATw8Y6ITfzdjgQ
4HwQRXcEDQLsUbgmwi3EMO7g0k/Oz7pEQ9u4va5fuNc1D72zzV9//o+SjOXiskyWk5NV5Xz6mj7t
XmSm86LXIMGzU/VpeBq8seFLvr5bfGT/IDB6R813fh4CpePEHOeFFMbezyYouE5yaSQ8y1Gi+1/o
5VD3oreJxZv7GQzOJfrs3Q3ApKTRcJmB+wjIsGtWYpYrlK5ELhZz4CK0hqYCVysGnjdCc/1Chc3P
v8yOO3iA57GAEgAKk3TNUS/ZdmrvP7rUGiscL70bHa2hxkZovSf5xQ/sLvfti1Jda+fpIbFdpPFs
9L4ZArGlBOoYSklSLo5X2wPg7Km6u3ikoAfQV2gtM2JEr4yIdlbcOiVO01nfv2OXqEFVn9YHC8uO
wFi1GxCejCahahgRyyhjKkpVmV8yL+1fJZbh357JPJIG8Qmxi9Fv8ngQmkqYiKux2YaqWHCnQRG6
iVBHzGl8ZEkutaQbhFeKDZMX8AQL9eKTR0qcof6Cnd03Vukt6akVl6Za6UcsrZc1k4kFxS9MUahU
r+qriefsXuOXYatQzHeucrdwTwTF0Z/aMXPRbjhSk0cDA2Ja39Ge1F1w6k3RePZEQZqme1xM0Nbl
7ItBq10FzMvnYfkuO85XMlnD9K+gAouWp+VvY7sTCvr8bTr2Id98dm0o3pstSnkHqmmwkg4Vz2kD
PN3kVQC7IwgPfACPQUo5q9VXVH4xNkQXNJor5iHvX+EQG0tezX8c67CFkXqDTFxIxrHMNT2TNq3k
erficVJz3ohR7KHM3/dSUokkagF6colj6Yg0Cc0gdDWrcOKtdnlgq/qBgtr6JGftae707v6isECT
Ur+BL4SpVyeZXPLoaa8TiRqf5vdjXNUEvHohwZc78fkadRA4kqjzj+12V9MVAMs6m4E2tKqrK7L7
052BfW2idv37NuT76xlGmGCi/SWg/yV0r/PpIPoOBaOR0V3EHu+wSUgXMhnODtjb+JHAI9UjA/rE
XF09qmwH+pZo+J0UZuGKo0itZxRPURoi8uTkv6gIeeWYJXCtsToq0Z3LG9M3/s5y9hdVcNwvvbPO
OznOYuosRXE9RXJrqiEuWaFLkRPvt81j8ebz9FgeFfMvMgu8N1Ki+B7iuds64Lee0KeF5cWyBdyG
u+0xWi3iIANLZmGMah5vKnXvHp+RlAXvgOOYlTCHD3Nea04QO5b7qTSTvn30QDqRY3z9ROIkujhk
k7Yfb8A3StBzBCGGqDXIhPkPyMRoMYFc2nmU9kkxkNyceQAJBLoYeyC2sEZNDbSmY0sSAcupSaBM
bE4SsfpyYmJzVLcRIE0eza6E63wkpZWazAuw/ZW8pCS8B7SeuS/xeNk2+VDfNh1KXh0RKLnHbrT0
MoRNsZJI9/YPGUNJKw9+DPRjeIYPJ0ZEvj+Nqew9PQ0CIDoPgq15yPySpR08VRdzsYd2IO5ujqM0
VQvU+ZGQWIlmNInqJ5ZNPOkVtPUTbfzIM5r/uHHS3YGrfIpfN2NIaX1kMElZEMeJ0U09nJqx2fME
0E+y8XnpQs91mEOBoLWJPvN9G4AmSDp0hw28ck+JmZYEfXbcrnaskV5jfghgmt+JV71eHMSprQip
nRDBxtdONOXx0ZMuSW1PsXMI0zFgneIFrArP1fgKMAJCD9eHnJw9zLgX5x3KcMNkM/9W8ky21pH1
DVZIHOnGNfY18wcjhHCLQuuphyKQbh6Y5jYI/AC6yIA5iAYUi+9BAV/8oxnljbsekFxx+6T3SFU5
9NVqvG4JBfS7/6a3xZlat4n7ox/W67vW1xhd0MwJi2iJ8wLqSnyy8NCcRs7hdN1yR2AKQFi8b9V2
GBTiJ8cXUYr+SG0uorioW+53tgxz+iEQPji3g0Htqo3wF3wdgzgoY4aEq5J3NtIChq0RZGJ/P0xZ
GXHHUMKVv7J7LVN32NBR/rcmxbJde4S1DomdLWJRBh/QNqv0OmCEmOJ8nllGRw7HDRCV67mnqGOw
/krXUXW0qXUE+qsQqZQwrA0oHFq11O4kPjtZ4/hDIDCrjna//tM0YlLbE1A/ltwV9ynhXyrPvlsM
6AJ/fpN/t7gLvdR+mgBYRC401zq7OobsVZhh0tu7VxtjBMfOKoD9iuP323AiWTAOiApqf65JrEny
ZQy6o0V67mnS1G0YSKxn5GA3IxSDW+glTAs8pVaYVRdwY0HjnPrhxTwKrEWvNJcVnJ4m4FteYs8R
SNHG86YWY+qoKCpXhwPEPE+KywOiUJ1VUVYTq+OF7tlVf5tY/YHeOQQliGnYovvhqY4quCiMmsld
ZYi6ye+Ox04+ja+wO5BDyREoJKHHxSeZdBV0qk4eAgOGnysyN0j9Mvp/r2dSwc0+m4BN5yb2lOW+
U/Ok/oMsVYIdPJJPt4nSfl+IIIjgSuv4BtUfOlYxcxkcpWJi2j9Wf44EHzYZpmTdOtFH6+R86FPY
DlmHa04CC2xxTlxn9iQegC0Q4MJ7Y1AbCCsWnFveGYj+yTzn9MuDVyQuPVX7ljkJN//TPuN1bL0p
nokdG6hBXAOGyHDiV9fpBV+74zbxpaej9vpUctyKK/r9qxlnxEcfrbU5LFh4zY+u9XZB55kjoDV/
9J2EcaQ8vFtTV/f5ug3Y6jay3e6zi7ENfefWTmmgcnGwKBgQgwARvnPah9sKiK1XQzQK9i8y5ms7
/9EToxBCmh2xSXzMFb0yPlBaONtODlt+R/Xj9FtRM2egV2KHXaxdCB4KdFk/I7Il96DzNz1A874q
1/8bZIu8rnbte+y53Xjv+8zS3bKrqZN2p6aVvHzldj0ek0nwn/rjw0VCV7nP2K8RZNxG4gvQu4Kr
dLwzhPuv0eIULa0kz6ZeBTX1hsPsz/xhspuxh1B4kGi5o5PeuVxKmEEGxAGQtRgTLCgRyDjLznBS
1xIT72r0XCd7ne3MnRmc8nDdhSUOfk0OPIl85yTHv+0MXorQZy7IX42Q+MN2nYPUptRjnYTAowYC
iHk+cECH8+uDHZm5kB58vNCq3od8zu5Ta5ym/fuu1RH+tSncCGSn2PP6qpR6AZS1WFAYB2INyUTh
XMmPQAHsX2IkIoKz1cTPHhr1LHakiZTidWO/DTrtpkxpGEffO+hhz/0UglDR/vZoPckrUZGxpxZ8
Cqyk8gjitp2KGE2PlwSkQv5AmnQUKBO/bL9MXCUEIFIncW0W/KfdweN5FWqW7Q8ctu5BE4T9JWhj
1Dfeh1T5tD73DYMA2NO1FmpNrBERee7dBC39wbdzkY0KVQOYHCkNeFVqva2jE3HKj1KzN7gtSzwi
C1TJGZNhBJVrw5y1c++XeN3Vmcmm0lfJohQkWYyTJ6RcCttO3NCvnLS3+jvPRo0m6nxWfl4cZjAF
Q8NMo2yuLDU4h80AgoQYnKM3/vO3FDztClJUVxCBv3dITOCIRL6g3s0PVvfTtmYnLVdDXkGszu1L
Z0j7EbdQ1NeyJRQwsTRICzKaf4thDVzUejiwTev0aG1psUYs4NZ4QUe9+CNFmOO2GlspUQfnqj1g
YL9rBVbcahJDVU21x8q8og2uR0C2e8GXGWk0DPtRUZOQi4/13HTRR4Jx53N3Czv/HhZ11hLgbPUS
3ztD0zBUs1TzA4/uMHwjp60pAt8H3EKMO82+ltsFox5xmAxPQ9amX6r2kWBtaF2WJjWJ8Mn4tihD
ptJvka3FWuxmXd42xHaStVyfTXHWBl7HJagaEIpA+g0QvPaJzDMXFjyQuV9/3/HABDo7aPvjIitW
bkyHyC+p1k8bEQoyOGTkd3g+4nZQmxowty9yicRioIdk1rlTId9CTQRt93z9YPOTcwewe05bS/o/
4WZBNZRfvsye+Mq0hm0yqu5x0iC+UY8DkgxfBzDVWeOAV/4NzgutElUWDZm2S27tyGCrpuArNxF+
bqbMoxNqbiGTkU/fBcl8uPbhH87NPYAM71OGrrqh1tvYxTgf8wYLWeDCESzYgY8zaY7fLG2PHiE/
avyZx5oNUSRrHitr9JA3NkHDTLHURNzsRtMsAy6g0F5aWyTJYqsa2E7YtVcaFjNip3wqri32wyV3
ilnp5cFIlcr4wo9Xe0iyTcF1aYN5OEY/MgOU8BeZnxw84G048F7BRQDDe+v8tV7irXNppUpk+B40
js+yZcTc9jbZ/od0l+LOtGH9vlhxymlGBn1Szada+uJsAgV9uNBWgW9JYwu6WLAhJEGO+zOTxWU/
o5MgXgW+Usaby1KsG6FmNHT+BetRCMhmDA/pjIkBYp/moCQXOmkPXodo4ZJBlYMFwLpe7kbdmBK/
4yGAvS/gfRuRg48cfaLHuTckpCFdYvVZ7QsHsXDr5nWl80Xleg5zlcarUCGt7J/nXUXCW3ebHhlA
SkJ5RkBoakh8QII2vRmuBygplGRGNHtDMdGNQRDWjinQar0IwYNalfu85ibNOL7t4fnTpvFvJqJ1
429lyXzaZPFLbbDC9Uhy+dSCPBmxYBzHQvP+I745YTLyagkYCDQ9c+Hnz6cZ1rNihg+gH8L9Ed9n
a1woISPkBWVCpOUNX42u5vwf91D5Y+MjViWUa8APzH492VYhlGXyyyIsyA4nu6iQAtgO8JLIgH+y
6RU61jsIHONSZvr7D/ClrZy423vXzsmiTMl/GdBAdzo5U56cKdraafdAMZEwZLINo3BemMu6AWEE
0tdIV+T2jJMySLSmKQbPFY+kcXQAeNH3oFLdOe+jh6nrDLhsdW0kaJ8BZNma78y09raBNR5FRYB5
ZNSsmHtPxhrUE8wOqGhD707Hl2WqTIULq4PqMJCizBtQASHOp/NPBKDxyC+zvt3yB9t1aGE4h9yr
XEdpMaaFup/lrE98QDd2lGaZXWvAPP2BlYRNtGIRAOAOXgSuxOleNvQQCjSNfRm+n6cZT4+H+83q
x2o/PyFAXtESE2hFDbwTXdvnhVDtElCFPOjtNxorR9rmpm07ATITjkPYrwLmgwxSaSDVZzMtSLmd
PHNU3S7LIhWKTBmKml3ytrUoFST+wpvsMATgi6Baz5MA4wbo3AvtU+FkRV8foLO/4dYdTbSE5gUN
e2LjVkJA4dOrrBvCh1D/j8jx8qLqCqlz1IGpcX690urJBwKDB03WREXmV/tSYElNMIpoqy+oJ6lO
peYgzC7Fp1Q6gqqg9aRGShl3oWU6KDZPWMyRvDndfXVdoYKLTzOyULHMo2kvgypOCWkj2+elJEOY
I26ck046PgXavma8zBwYyADln0jIbzJz8KGKLFp9Ykmgco79f9UUMUKrIHED2RLVOTZQ3mRZExkr
E0RGez4HO+cJc9y3B7NY+eu/BugD0nk/eXp2sGnxePYwreAMXVQc0OHSrAqfvXPEo9xlle3l2Cjd
+PstvC7+OfDYC6EaNRtxz5MpiTni3nVUjx8CFOLc/DO6lj5NCj/nANED7SB9YV6jclkruifF84o6
1NIYS0vbQw0WeE9SIlX/YnEnR3hu3tPAix4UtgMSKDmWx0TNJSOPrPJIMh0uXwWHNQLhECgDAPkv
bv5k92c2ScbqgXNl9XidAijr/qcv7tPwCOv2SUWxA0yqbstSNOPA3oI1zWsfB+igLdqv3gO74Dm1
COCNrOhdS1VT7XQ56tSkoCgLSBrvsJHWyYg20yZjtBZZgCf2ZU/27FYMONxAxJxzMrX1joYv4nkj
ghJWhBMS1JkvPcg61QfSUFWsuQVb+dvZkykHdPHrmltV7UdLsrBhGPG3jp9VU58T9mqnq819VF1b
owXkuWp87vXVFzN2mJv4e8xcojMANxrsov7C61oVlVx0A5VCGvC2HvDoQkvXkDorfhF0eYjvBHP/
RcdvXlrfIJjMFheWwLpb5STfARtyCxpcp6GOs9KoG8OxJqklwURtAYAMhCU1ZPXA+T/d3ln9z/vy
kwapPdnqcYvbtnpGGTaUIxWv9Xw3aJ3fiJxmgj0QqqndBLQukTnpOjHinXKnSj1Nj5sVAkxtHEz2
nkSB+kBz/3mJWrEXKvamVALDOxiM135dDdJXY2Sh5sgpNyoPNDdYJjgEV9vI65z8jxrmABLcUqxQ
H01/VIY84W+KgISnq2U2Iwa4gQ8YQeOXY12u6NDtkGvp1TPQaCLsPsxHnxcsUTEYx64RntlKV+yB
hS9egYTe8+sZPtCyq/bqcHOmyFbAdwPuo+1+3pEEwHAI0GK2tkUxe+pCoKErMVnoMXAzDHNU3vHj
vRH4K5gYrb3iayKDMNOwk9vNiwavCZLigjP5CvCdiGrZNCciIMHwcsPzs7z1b2XUH2R6TJO9Jeit
dQ7UEv+SwqNcW9iOEsC0is9WdGPgSzezJI74VB1ZzYr17kh6FDfM8rKQimeNfx6xIkqC6MybsAoT
xpw3354tf0GrcHHn+YivKuIjUrxyw1DGopzd7JnK2LB0GRY22FT+QpaGB7YEo7oxy+Oepe85nC6c
oxdy98hzkushukveYriFtENNfxHe71D1h598uVuxSECjm8R4ytMsuH785Yl8bw61Kloi3ei6MJ45
nu9iE8BzGyBfQIw+hLoFQhMINjkhve7J5C/hi2VhxaSaN0D8SNcBLM/Y0bVFleQaBLqy7bBdyQAN
6nGrALt/SRyRrSW1IbLBq8JduoqnvZ5JYeeiXKQikXnjroiNeh8PTSptMR5kPqvgAr3rUyH+l416
N7nXEoRxqXZalpHo5QGimxx1Xl4YMj+aF9dbkaeN1+/rpi1gV6F5ZiVk3YvckA9D+3PxS6qb2e78
J4zYcFTVpL5qrWT8l7vhRa6jpp3BTXJCKmFIhX0fUA4aL1gUWrtz3I0NQk4Mqlh8xyXnX/noWJQX
5szGle2A5LnHxzlreiKkUjx/N2eq/tU7hl+K3CEbzcj7uXEcJHNS3985foYb00BbW/253xkJzX4C
hkHLJHs0xua++j5vHlmq/BBZi37xqqIqBAcRwzyBACRB1i6s8NOFojv7UjAdda8u7lR8axbe7m+I
TNizu6MiD4q3hUEJ19az2y3U5lUFoCq7WB3pw++Z6j5cZIEVcYVaKqOkiTLxguuXhunPUhQR72UD
4kC9XHoa+os8tiLckc0HUC8a7+VUkYQyCxC0XdCe35s9bdDnlyqaJ1eTyIRJ9aP9G3fpsdejOVpL
cPd4EFP+YOo75R/UoINISEzcixlmJ4CNEqjXfBhyc8ZUj/Qf8FwhgkLVw19nYC/x7pTWsmYUn3++
yMpFpn28mJeVJumQAVURWkrOxetxPkCfF9YwmLFeckaMreVuiHnZapQ04BvvICpzkurRPGZuCoCP
GInWYe2rG82W2+qtd5ex3COEFr9RD9su8rPUSCjMmwAvc1SeolY9KcqDH+9tVFM6BzJP9QNOBUp8
OeH5BKmmtUNBioDT74VKsvo/kRq7O8r3SlzIReHBPY2gXtSSfYZNmWqvUnTkLTnBcgNuSMCWIo8F
+Sds24rK29GMnn1ID+2Z+lBUNFxebz/OPvLIVPUug86cd66vBccJnbiDLU+wWznPsrERxD4k+jsl
PfZmd7ATZu71t/nV5iWGzw9gx0lLPXEScNPMLS2/1huP2c2aYLH55/CIQdU5yk1t4E48TigK8dCj
xx0AIjaDEL2EudIN4zG9+eVSHXYKWHgXF5e8zgglwduCNQrR0sYLvf4/uIM1mamyuuBzlO0pfMpY
JVC/GopZ1n2v/kHq9vW1P9CoMViDG+3HMZNAWAUNEJKy22RZR5dHX1xejuOSTojv6Y0YwKjY3xNA
h7EgsvG21dquCJNXMWgf42H61PTKANeG74bzOOq3rSQfsxhX4ZvWFh9ZKdG5X8FBoFRoZC+n8XaY
qCi2Sxxx4lK2Aee2jX0q17U4y7LYBwpmWpVzItqULu2uPqc9KD9TwPPIHflZ6IOpdKToBN+1/95J
nXlQS4lISbDyQ9+j3cZgQLEpbR/UamaYu6OjVK/vhYvmf4i0AlMwermY5BfuNSl8MIvbIwIUeaK/
jE65XXPVBL396PInlGtUp/UKvnifFwAdZ/WAj6lEVVAln0E0AO64mTPvjaCmD2fD9KVM6ocO3g+O
m0D2vZh827XPUtAavSnNTWGzuVoaS3cU760J6HW+ei7w2tN6ICxM1fEqe93iM7naUHLrExTqxkDg
hpFwn7e6viFKlkAxTT4JGYl9e4/8Z4kloYfHpoIHFaSFB9AJ6D0Q75VbKhOizso0XdWTpNfYR7KP
dhA68ejJ0uJLQiQ5VC+C+lGJXi7sEQMTBt4OjoJYETs1PXb3ax2099JWZaB/reZ8y2KJ80Ifbadj
dIgpmpvOwgvtShtreUEPOpoWXmk1Jk+0PPiOcqyg1Mc70KlG9P8GpcDTYU5iVXtBJCuHcC/JzFtB
b8LQmN90qLgZraNFhYJDNPpnMuiBAwBrkkSqOVG8acM0APRTv225bTmz2S7GsBhRbe3Fn0CmcHMP
yAdmgNW/kJ9BKQq9gTXxZbJkno7cUXYMoHrytbiKdUJUGWfqv+9r/AXBE+rOJ6ll90g0alrQ2wA4
GCX/jtEEVF+APN8JtTScz+NKmIDaIlZbsO5D7TyoGBMCkGZgFT6JEeHiX7iTJpK6cDl4gyWfVGzl
BKBXJVsqXBOdd1NB462X+y4odN1bEJdWKVMEDvgIb0aYRvhFTV0CFfe0c2FmXe0kLy8jRL1uzhxF
iJLRYC+Kak5t4l8MVyCX/6ZDVYBmmjZR8JAOF+4+1/YwlaYuQGQQCxCl6pmv6U4/AUs4l0rnr+Kj
jTSR5PN5Wq+89Gm7LTQAYAxG724Vfi8LJ5+N7cCWFRPhRPOsc4fV8vqXR1s9jnC0AcPD/qG9ZMb/
ALw34bhDoglJJbd5+cjRd4B07PTR32p00J7T1XvowqvZ2zH0DxVcFt7R1J3UCbGkihLR2Npym2th
92STjx0AGunPmh6T7cXQMlfkqVwvvsdUMqYSD4yWnyRMOpoSt0KnqkBoUYopt5DFiGxzpTWeHAuI
1k+LMfs7BaYcpz61ijfIzmtX3WdxXKuGcZ0qsmrBYmJFw/eAMehSNNJh3eM8w/hSRVntCHAJlIjr
1Y0cnM3NOJ/uVQTcqhn56ejje6lZHbG+zR/+bK39zt4BAaQNkH5DiO/ITHj+lPLJnQbe1sAnddb8
sTocS2k+RgDSetKhlGGxf7gHmRbmxZCnvBF/cICsmVJMy+SOWsEYI7cyWRrbZgfroR71q2yVu2pz
nBbxJuNTHUZJrKeKrdtWyoUBSKiOXSLk7DJ/b6lr/WYPQ5Sa9cfhc4Rd2LInDfCxjpWJmbKfFkzK
CSM6GwU3T3Dp7CiMbxe0tR/p45wBXPlRHcdxbux0JEO+55moB23yba6/yX62mf0NGZG8HJA2KmiE
wUHkTFfu+K7pPFAZLH0xLAF9yvkV9XpBj2XJb5HUfaGFMqtZ7Tbp687GB2fTNz6JbobW/frC/ZQn
qb6pBGPygjquZHpHXNYQ5Q6rQ88qAKC1n9zpMVWAYkXi3WTJsGFXehKAQdWlOPxZXNJXuucs44Ni
VfAe1QIdHhFg0wJ+Zm1gVwwfu3e1DqIR9Nlqgh02XmuaxNAh1Kd86aPu4ZqUh95a0tAsnmP+O6OM
vO9YVJEGJFqeaA2NW2REjnRheBwQdrL+QyqNdsideGXTmXUAuBVweglq4F+yL7Z3C6UF5hDfdGT0
fviumsUdbfF88d6r+HU3+zvnY4c9mAZR020RbG5Gy4cKP/TNoPFi5p3QmJecr+erWF9cPAMiy+/z
wH2xfx0s4ojM5wYX02WtYmdRNrFZC/4fnDxoEzGSscs/2mwQWGCibDhHlLX0TqjLsCe/HMmh75xB
7G5BSKCNT3e6Jwbku0GTLJUSoCSWL359mH0Kp53mQhYTHL4HiVt2exHnaKBZPlRfyBOdnhBtG72P
croWvHrw1gtRvovZ5armbhf6Q0xtOEwPU+hSZ2gHQ/59b9m17zSn95OjuWI9f+GW5VG+JDt3CN/N
nxlXpLAGmYnJYMPTNl8Klu9AVNRWiPtXZgFgHM2QyDYXwLccoz1PCu4zOYmhWG3Nf5l4ZcLuIZMQ
UCP+tm3enw47zjzVezH0sQa7qAW7pOANli4HslCJV+t0wWZiraiwUTyM8sCVhHD+qmBsFckxoR52
PgB08gpQedGjiCqDJXj7REw/cIwdFNJEDJnPss1tFxUUnPe6nQ44E6jxyBhE/z+D6D3M26+8NFr/
8pJOmUUL2s6I+3sCXebh9FVWiqNBhu1U9Nc8GoeSJ6wwtQXlmJaVx/er4vX3aeFxAbLRWe9qey/Y
41GobNxM6dOf1imJ54MGXoxLnIDqj6TRmgoWNlJysX9YdoNSDopP2t7f2XO1vMsGBy2zNkU4mg9P
7zXyzwzluhqDPhKt4VDvEI0lUvmpw2iM4/piOgNmj5RpdL9LVu6EABfIFf8XUJlD/jVFaXNTe+x+
TsNJ1yNATu0gG6JE3ISJ3Nn/JVTuaDOXi+MYAP7OGC2fHP8/hObBDAxk+rl/M+N+UUJ981OzUWvx
FAMR3GYG1Fzc58Vx7goMoIKUmZmxceUY62fo+pTVZwGD5iuGdLvtXbc1c4SZ1hm63mhUNd4nhr2Q
gqf2KhzmmYZiolyJNMnuIXC+IASyJlRh9Lt56SwARTlooWZm1R0l6VSzQA4YEh84qlWAIYn71JB6
EnHsVzMGxMkiufQxHVPOIsKkrWcxf3GuknSglAr/TNqYuxchS5A3ivbTGJthpjUaNFBgcp/un14T
keovum+csGTIl+wMgVgUWquUC50lhjkysSazyj0brz2PZQme20vNHpk+xdDpTUCHuAf+QIut5lxh
vXEyr/ZifAa6w6VrupDLAStruAH1yXNsZqd91xFIaTO7MCxhI9QDuytc5OrvtbwZORyGQTt3JM3N
Z8kFSwJcrJkzNS0fzlG/YHyf7aL8hmO3kufL2DZdgHaBylws2I/6oOtpdnbYyhrxSzJQX/IkwB8Q
as/PRKF8OwzwjuEZaTStAv5Gqy0vmW+A8kXS7euQ0ou0gF46/qy1OT2VMAT9b7dcrtS3XIstWMVl
YUPwAu1z68pik1WZdNSAjCnnKkpPVOV/3sWSxY9jFBo+DQl0WKvUpoysh1rcvFUtjaz3SqdBxgrx
NZxCaHmWhNrwJU+C1wUa/tjANdRBugKwfJBHuC4byg+k+PajpDQu30cx3XC6+4ZVeWa9Zaprvs0J
VrlfWIdOOwGaFoKFgWTdk4d3woiO5ypVvTJ2BN3CxoXeRK/jpogHwNDum3BXaMGbyDEiiPm1hxbR
lvpa1dq1puMpiDZ0HBKxnb7NfK76OEJ0Iq5ZyCWyDFHpwJjIGQXYwLAY3cCEbRXR2PKDo7OG5Yyn
tNJk9Qf+wMubuZxzdBRrOWshxHhiVGiMCKqwizQ230Vy19NfwOHx9PLeineXmloHCgJ4vyjVGk9O
bPyeR3QqLY+R6JahmpYYePrmOfoMFhHr4bvR1rduDMc0W33j8VW2gI7fK6X6ugkzkPy/grkuR9np
I/9VKS7mk3hoS/ra/rrdVZMkPK4pKY/nAEns0W31iOmxGQR9JDKU50iC7MOhmMw7YOWSPJV5ixY3
98Mjn75cWJeTZBNF5ZA8+DLNvRSwgMf7+L7HGChHNHoR0F4tMpmtEJw9c83Bpu01Dw6jNjWjTHDD
dB2vVTpNbjcItJJW6dN8uQ2Mj9Zx3h7UX4RwirgqUtSKVVlpmwvb+6VB4sazp0PnMq81hKi6HhwK
pMza6Smm5/zLc4PApknIwqWcCyNwSWZpGvqPxYQUsnD1BnxS8M1UzRjDroycTvAepLT1XvMowT+q
HAhU99guomzOhCwg5Y/6FJWX4+YKqt/dNliK/Yje+z7OL7k//K4fR+dulUO5sRV0Hh6ZuzgWK6ZE
13FOtatWCAiw4jMiocs+ILEDmmUqn4rIRlLV5uHuPkKpGCg5JFcxnndgTga+TarN/pAtwGi85Z3l
E+FajCAKONh5z7imJx7YRYIGa19OoOnr4UVQQxVNxLuQ/7F8aI9IfV3tg97bC/vvqNGFG9vKPmA+
WW8wpawNtkWzMrSKj9LeI3D8lP7ArT8+1kby4y6X7WDNrpWYJ31p0uM/4kM5LmePftXE0rf66i5m
ljlN1HDcQxZotI1hu7KSBsWevJRI9c9ju/t1UsJWYJx0hJU174UBJnfQ95wq0Zd89uIgfZEJNJiV
q9Tm46AKOIOa4IdAsjyJa2fIbaalBu+NtZBWUiMFykXs+dKjRQcW3ovuEGTPe2gIj6yb00gJbY35
93/IHOuJ8mvQeeooZvZvdCD7R8ayqpOgBNokk42qFnxDhdo6Z6bMBDSyKXq59ouTVzC3LFn9HcLM
daWFQKFRnpx8bfzwxbFuKwppA/OodyOPz31H2wljjX4iW7bPWCvq3Foj9WYd8A+7GSgpBxDM205r
sva4bICmXAboNP+dJg8haWa7Ykg++mldItchnO5V/c6uf0O4Q12cRE6aViAC5n+vFXhXbk2aUvfo
K/93/CEVBbXFmoJ6T2iaPwin4UJdyFSDHftnPidyiSVlCnyxRtsDXca7BvPrJdp3b90G4SpWt8bj
M8ZC0CNZXHKMvfYBfPo0tDUi2YaAP4GOsxyo2gd+dI8x4ONCHRF35oNFta47Tdl+LkW0D939qQiq
ZENDKODS0GW4Hljzezdh3XNGUALDKjPemhhoh2wQnZdhQ1L/eka3lZDt2gFpwvaLGEv8oXQmXtv5
KYKvi2/KaPEGn0hqDP+YPMu0NySKPUrfTlJbM9dkm8r75VtFy3b8jX4HBejsGrH1u6e6HPpveVS6
febacH6rdZhwmPJuTKgHHDhrv8NUSeDNe7oBSMOe3sEVRwLBRoMTnIrl613XreSHbBlYn4Jc/ECj
ld7Y2387HIL3+9q0L0F2Fu0lxymYfG5sM12UtHD9sSJAsh8Wn9dM+yzyKdhwL6CjGHodJPT/EDhY
q0Ny2t98zXBuLWwCD/pNaTs3ZCRRjpXKKIytpx0lTZwDs10qUIAo7glOKoLewQvBvSX+ht5df5te
El1ZqfKCrt7Hk00//IlzGMTLa4jbBHRB0fPW/dzHBeXd5rvYSFBXcQxc2nhQZqnK975EiJkixgDw
XntJ2lc2wDazWhCL4Mg0u/v6fBK5onzxz8xmSFsHpOg5DWOtlbWq8+93WB9kBnF5UIIwRhChM9o6
dRmCrwCAxNP61bXKkQH/TPgmwn6rM14EBj5UCkJCc2G1TFEwAaA8JTsFHEEyeGk5l7MFQIUgRaVt
TZBy+T/KPh0S+tAXk21i8skoSimQOOwOwNa4S+BErWbGG5V7WERjkVkCTLDntkXC8JYJXF9yNWV6
/I2pbPvsuF1ZGMyk2fKH/fcLoKCEZjBqomskA/vN4TJ9PmTmbrYazwYZE+NZ3BNWCLzbXtQ+0nsz
mmRn4ldEgwaJgMc1qOS+04LCg+i5SIgbdTjZeY1TbhU/5FxqSv+jk5xWqgtnokhJg2urXhmTuvk3
z3jcEiOc3zkcCC1kg4KMp+DV8C58hpQyc7etpWSyPZxD5iJrJLCQJ8tx1tD8MA5z5hnVJ4cO+Lmj
0gjEqOQkXHteNzGGYjd+LchsQbswpouuUMH5T/YPV+59hm+O132A06QpNrLe+7q2bIjoA3F3Exuz
UDC2QCicQypc9oTVIZsM4OnaF0Bc75MkMtAp5aKnoaGXMxwC3Q7jlNmr0+zWEeR6cRxHgv/dzgZG
LNFAj6Mg47bEbW8RZhCj0S2eDkhkzFRQeKBugXyvAVafeXqAMgR4mOG19TpMGsraY0w1c2KUCYXz
bFJUvoohm9LDKs1j8ZvhyJEI0ELt6MwId9P1Glwgv4P+2a+6Uj4qQZ8fI7kesc1F8v2ixfbSYLiJ
eDk5LbI1RCI8A0JYVFXRQUUgZKbnJzaMPlcXW3RMuwyrIkHJbsymMH+UiVMg6Nk2cmXUjhTpbHVm
cDUR7a3fOgH1oJS+kLfKxT3twFI4U6M4ivz/+lCmhSwL8A6LY5zr/YnTJdSrISOSspmeYN6SyfrF
nnxcLawNf8ERl8o0Hed34HrhkqUU23+N2Dm1GqjYfiKZJzIDf4axkxRfVYOJJP1jHO12W4abJMfU
DpgYYneayc40bccnVCSq9eDv/K9gT8fmoScb4/ruQgetJu96ykfIT8Xyt3YeiwR/a//rBtlOtt7O
4mjg8nPTvFPZP4z8nxrRYADNMqMrfX0u6tuSNZs0vrEfb3mvVIAciYbP6Ft3nwOJQg9QG62WD4dO
u0psdD3XqX9JzA+3ywQoYAi4lt35pKLthQkH6NXNu+8LKU+xz+BM6q2Fwm8lpsJI5VdQ29J8/c+B
GQ/WYY2ssRXhM2kJ+adl3QrfQFR2pFU43Vx80NcvZB/zpJB6AuARlMvmhy1yJ/+L+5tOOAgFnNbd
N6pyc9TYnBSzb4s9IJ5D1elAIbgZ3/JFjKymkZxhzL1+QVMOgBg8P5h4J6dES7XnsM7ZqSibAJLG
r68mntRem05pE/UCkhas0jCiEHqOUg+wmsjebuwQCeQzD/hr6BKDe2n34a+qpz5jMBYX0yOKyTNX
3fdqqv7L9Pa/9JObH0Y9+X+6BEmU3fDRRl1p/iq2qI7QbeBdlaO7n7GkA0SVwxVWDCIj/n2er8KU
On7tm3uOavnEp2pSd5y1C0fkhJvLVxiN0MYoRDqHFa2GLFRqFkISwKh8ZzTjeN8+lKKn0eWzrUwy
8l3CorWIJ+1YhD0VAOn4Hkyn/DsVrg+cGbt8kHmGR+7R2KFg9nBFl7dnU8s5KVI0CFAZGSazuR6e
Ct2kizieB+K5DZ4SBXfsarDCrPMN4C8MVUrJe5ug8c4d5K0VMfGHvkub/Pn7qB8fn3PQyNJlPBd6
ET08V8vzQsrD0FOY6TxsVzezK/+zs7+2uGOvp76t/OR0tqHi4XUCp70r0q2zHHrDTww4aN32s1NS
6ecq70v6dfGwtSxHfiYAfdthj8UApM9Ah7q0lo+Qna16tHpRKrrVNt5jo/jxvn552X+5+CX1mvwl
cZedm5QT6QZ29WKML6vvlnR9ih6p+7i2TaowAORmvyzuBOBMDpRvYES5StGNuQf9+nhedxDBr6t0
VJxMLQdWGZaXVqWVY8bv2OtAj+/CWAPZ20Oa6ro3c79aSyoLny9rt3frUV+Sp7jnpB8BNHw/yDY5
P8Z2S9ZOMgiisUGKI3PsnSYj1yRpbHN3R5mJuGZvvaR1JGZhiFKjenVLrd8dE66BvGFmnr/4PIm5
aTiu0WHivFXXo5/kRv81rwVIOvWo+57tjP6uXHdQP7vtmKi66oIfnxOh/ByZPnByj7n25Ki8xSQJ
mZEFY97TPToZKSFB7nn9rwAlyBwITpyne1+1mA/ZOZpZ9icWqk63cJVIjom0HCGjNgwQnGKOQyGf
ws4yyJdD69YupeIBsaWAiylnZz7TEEsEzi5xq6+qO8zAhLYmalQGi2syl7t4ISfnpUl06/GGYsKy
mhInaVqi6oIzAJ04C/gXmD3WvTyBFCZ3BZGdgOPRRyd6nYZIfIj8vZ5px88z7b8VVZWt1Y9ROFNS
C76FeJq6l2Y5ytpWOkCsiXxiUBgXW6bQTA3rB+dE6VPinwGfQNqtiV7vCivT5cLCaHMgiD6tKiLA
KXgfJcEdewY0vY2vaL1EVt2BYML9EzlujhIq1CEMg3YP/tbw/l//UGcuGsN68mgf3u4mu8J1gAz1
nsx+C9DAiuc3MCnR8C7aRF/IjYssOYNNT404co5USbTs8KzQZjtG1URDBd0SPQyA1HOcC7tgwjr+
y2HkkiRJwJybWPvIbjOkiHlkEHAUhf/kOm04qJGVoh1piaHDYcw59yna+jQWSYLxCKxaCYA1VtW+
EciXkcU4vp7fjti9LefeHkJEmJ64kvHMWVaC9sz+uy+rFK2eikFc6PLR+VWwsCc+HS85OU705V8r
Tc7Oy6oejcpvXl3C5+rBmiAh0lwxI8QGUC1HJeTmFoRBWT342R67YbuXSbPJP/jG5pamUfxgY5rb
ZIMkA8R4YkHiR34nRhNx2cGLJQ7c9QxbEdZCn+oePqbflE5oJFkJyhKFUIdwAF0JORsrUhGacQVK
nrEM0/SSD1f6TfPnPG4MlUgUTg36NhsGB+GIP6e/EX5VjWhfFVp1Jt0wOeGnZ/nWe1EpYugYkaXX
wHWN1L8d+5o52P4HOaovGkQhNQKi+gYvRvsDJbhMJdaiKMx/0dYtZP3mlj6XAUAu5gbMXshqeDI5
UXJ5d2wUhi+SEwinBqxxY8vT2vB7o4GgwP+7URssh98KeStH19Byj+03kwnrGWkgUG0Gg0qKRALl
RKGI7X9YqYuejnyx4KQ3wVYDLKd6a0ro0Q5QFELTLDD3vwCwwALPYi7iW78opYZXLAiETMxKNfea
kGoCItlOyjxhCWe8X4ew0GDhYp2mAWNjUNq1JpxmvO6GD31J1jCqQ7E3e4RXjqRe1ly4SqrjrQkr
ulpmsUs/U1w1/WkOmdahe682miPaPUQCzz9r2OyJaH2c9Y2gK5vNaHqzGJ+V/giEUYe3DIwAskgo
DbhvYy5xi49wxXHNJTMbGx/snyu51RTytDlrYmcOB6vamnv6TiXEjlbcfILlVcxHUZl0/4QUbLIO
ko+eFRAi6/+gi7rCgmBiPo9Ps6lvZsvZgxmVCY4ny3jdPTh48uk934ucd9uhERAJkraGjo3I8NWN
HWDRRsHrA13EMQgE5VHzGDiKS1E+ypIN/rBewDxqq2fKcw9ztiYHKTBx5eHM/ZsrrtQ3hVb8xdEx
fbSiWfxgQAhpFcXBLACMR+gUt0wtGISabkjVkCD6xPC4dq6G6uJpFPLsWJDwScTFTpE3hPCqqwWw
b/lZxicB2VW0h4s7kn/GbGrOAU2mpavCsXJCNvSL25Ra+snWGzAfEoQp1LdH5BZeOGsX6djeTOl0
kagN+OJfTO8zq931eXxq6+/Y3Y8WtlYmrbMbqVXUST9owdrvstndO8+LTiXyDqadyiHBR2Zw17hN
9rcBtn4fvcWBV+/ft4NzxVl/uMSgBH1rDPqAmu+fvqCg4Eyns5QAn3CO1i2BcPORhIb1JfKdojRX
jbJAuEyjzhMeg3Lrmbw/uOKWZdfv38je+gnNg+AZhMhvt1hhNXrrQJ+oxD/XqPRzUCKyfG2qf9bh
nJqJFsOuFi9Xtis7tPjISdAtVpAGeIido73MOUAXPyk0kHB0yW6uAC90iGwT/8DjkZZssDSgoWCv
CL/TTzeuVevRwDOYnj930ywNensK2IKWefNLzUynriA8p5E7vN5P+WgIfYQ03uh/zGGtKfcYrjYI
5OfdoNN3TGsUCcP/H2azQaid0vudT7CcPPQSywc9pJUECMO1NfcNVx1KyzQxUxdyDgtV3lUKtJAR
+aslksveailC8T3fH7aOcGjm4VFx4mGbcRrTTDr33y9kLODuW6y5Uyfzb5ioo8Csb7uUi4ykHmat
VKOCxa4OiQvvBNeyG3UF8v/Y1nCctDvaB3hfgWxmFDlyDmK4HmbFkw4Ieo/fkOhCtBUzrsLr/JRI
QGjBPbx3HdWjO61zflWtrBN4rOTWeJr1nVlpnvm6CS60FMHr1RpyLtUj94rCQALQePPFB4mxFPR2
mVyalZdhUzfhLNdYwelrGqnx8LSYfxtxPlOWVao1/FBJsb240U8O9Ua1ViHG9q79nl+M3wPtKiCb
LWkbwwcWTGBYabbWzknVNXta7dqJKp10PXJ50k0aRa1f467QlLDd59fCgG2UfV18g4Vvk2ilkx2C
yy6E636YlgovU+VYtUQXm4KtkYRCc5a/6gOlmyajRYpfXOIbKsNObZ7fAb0FEQSNcI3I++1hsk/M
CmnJcLwPoqHjUKoLi3LNsDrV5GBTFFpqxVDtpcSTQBQGhtTvCXmanPC7C4FugO0KWH0VGMP5UBWH
xBh1zRNfQKC0LJqkQwH6LjiFYiiiDAOkfdbCzBsMSRUUU/cTag3RwMyOlGq5EUJIAmWSZHHCoCX4
WvXPZ2npNZHi52UB7H71Qt29HpYSzvGKOll07DVA7UTPjSHODqw146Z13O8WHRu+1flg7kXfyCa/
w/8kYQCM5aFlJ1J7UGC5vDmLUToWI3fN1IHNREpxEd5N+BwCLGhpnt3M2KOi346760xd+Rzjv6yA
FTI07ib25o/UKjBZBONxY1scLNaQuRvnO/JGkfAw/cnCgdTMKQjBeuI+cTDsVxLWplb6paxNaPtb
v1V3jhjvAXk05+IXfAIMfAb/MTgnOZ8dtex/TLH83Z2aiZ3i4jKAKco/mvLnEz0sbzgKqYMP/UOA
nMm6pduXYJG9X+/Z8xY2RIHRb4Vx12khOCncNwjDs8CYOc23vzAMQTX9s6yxdD72bz6F6YM1au1n
5bXvqNkJAozckSsuKHqFmy7wGi9uaGYdGGKgVS1O4rwAT66ATRy240POXK7ZoNGSC4vFczJteYMl
kUgpu2aluWqyA4E4taNQlMSuwtKMY/GqNN9aiqprM72f+u0zlGoH2ogZFhsybxpW+v0MZ+OJgIoJ
nS8z2C5kWbxeJ3olOSoC7i3CqToaBKHG/S/fHr/SFH136Twu3uqupK1Ntpm96eKJ4IYNtioXN1bd
hfrCd85VxDM2+hO+cQOwjA72ixPLeeR4ZWbZfG2yDf4gbq/mYN6+XlStvxsk/1LzSJ7RRSf+c45A
D4auzhuatbnk97p1ATiJfZ4QI9YPKlR3bArqpGvxEjQEX5P/TjA0iGeThN/oWwA5E84VDrzoeITK
KxTO8IWjRGbqf6EM0IdD9F1Z9r++RmfonyPxbqTfJax/XJxCaBWQvGwu5p9hTCZ5dCXFR06dQ45+
G/QQwQgyUAGwrJ3utyXejwRAuXXruheuijJ8jlP4FvyB0Rn8kCPSlD5FFqF4/0igkmzZL9AiM+U7
z+QP5hAe4E8uUbuecMG/opmCsp9ZOx7YzECCf9PaVQyUkDdhYl0wbBawf2rYxJcCuO6kxmKObem+
NCRcW7ZrKhD4O3ZUVFw11QI/NDSaZp6bmueeJl9eqtx5rPZxP5c+ngHi5qaU2aAmjht6m5ZIf1aL
Gdn1IJkz6PpOYf8QHDRxnGP1rYgyNmprt4XJzr++7Muf/fz86afR9GbO3iB6KgcI4aShv2fzqUsN
F2NXq4zC+J6BsZpwPCEcMQ0niM2c2LsqemcZUWqWzOUHRVlUECwJ48D277WTIvfdALw94BWyicwW
7xx91FPQW2n0l4xT4p5HdTAGaJ7smzFkHrcU/2rTRj3p0HHJa23BPnUJ6kX1DARhykSDTgvvHs5g
O84U1pMevo3b/OQ0UgUui7/ZGUCQF8ey52Y9VdDswbUfSxJyvZq5OH7PQXPgxGXB3/Qy+6nGWa7b
nmGL+6Iil1hvAV5n0J2aQXfrkGSK0/oQzNzRy/69BYxVFFfCgWsjLKUEoxzZydmWLqKxk8iFm5Mj
IiQKR287Dpg9T4PiecxNLPm7htmcRRZM8sZdWwylOE6SA/xsrX9dNzCA3blig44g1WGVbHnPtokJ
F9LyjafZ9i8t82LEeBqzhReNkS4XIGaiROQ8FqeoKJ94kaAOFcCOxfTphL4QLoNdLYreMblziNQt
nc0tdXjysdz5o+x9E8S7FftelyZsXm890uuFqHCLroulHO7LBcv39qIZsMu99hr3K80do8rUXMoW
G6tdupe4CgDZKaFA2bN1G7DwKKTMR1W7UlXGVhN58H6ALCy4XrXCEt1e7SSW9G+PG2TPKb6CgKnA
tzFOE4GJ/JeN9CYZ+bSZzm/UC+4r0M2A49TopRnEtn+pVklcPQWH3+J+5dVaUF8U4eCAtZxPf7Yx
q/IbaGTZyPAQ4ztdi4I6nWTqsIKiC/Of4KLjisqes31QDrpr6DgKNdin64q22C0uwxgbX2Wu9+vA
tmWaMf50abBbx1AWWemYWvMp/H1W2YOTKAlNnL4m3WxWCpXgbGz0OhoKlkrwhWmR/nYkl6tJ2uUb
4QFwP/VDyYno9Mh6RefZYJVscIBCtxf27m1BxDTCWLbzJgAs0f2tC4dTfKYvdrSJkCV7Nyg5Cr/w
O5zGsVA8Gm3VxqCcHK9RS2HkvSH7j6iaf4ySDGt8CHy/fwYHMra1K4Kemgj3DbFzSmdShAegDcbB
iRrrAxhHUvsM6i2c3oL3TK5+ZZBbmXL4Pqg3oi3k6QlQK3GbCLtL5ux9AXBSpse/abNWHJT1gov2
Cc6b7/Dy0FHytJhYMXRAYkxsAJ3mbw0TpWc506miZbX7whmL4o9HWqRky9diObX8ln6rLMzWOgGK
m7A9QWXr6BDZHWkcYTxuxKOcRU2FIAOq+tf4DdOQG0oDMn1PZpADgecDKSX+ehF73qOSk0yvo0ZD
jVQMztE5GjUdwaHwGFJuW08glGPbR1SyMFxLj6sSgzR+/KPnJ5kXOyfhWam9heGMR6PSIin8QH/v
PayqUznBOyo7YhyA447BwKb7a0soFLaON9/QcIICGXij72bMy4U0O7DIUEVnnCu130LzOjEed6gU
smsQNfpdpBe1blM5YdCd5s0KTDJt8Ddm53ZQVFT1KjKBn0iAloRmqj4SIwWsadDVin/YNk3HeKEY
TvfQZnmaPTOoIY9JS9WLnERerVobGMPPFkIMjzRKOJe/bnvG9QxSzH9QJUDDZhYvXjIilOnypBNo
+fUz//oGzOggqfZGhz47G7uvmqUFqmdMsjONvDV6bugQDBm+1iC5OxZS5NWr4NXpkh1BZm0FZbYW
kgQSuqMJZjSIBMTq3CR0tDleE3wJOOEHDoUsGDZWk0MNqVcssL6YHEerz6IVPOHGqnmR63OTUKWa
AuU4AkK5pkfzIo25hQ0LFH2iHSL16vURXbeZYQL9OsOOW/CRvy//pXZsG+w8PTpfbSzfGXSYq0OF
UyIh3E63k1gY7P/40+BfemVn26VEETQlKYuIocDSa1+342onaPCki/Cu+4ZZJ2Oayf3WNCtJY/aE
VrXhICYJ/ymjEkCf9SMFQDAwFL3OHPjWa1avy9N1r0F2n45UEvCoTfeB5New0mw0EaL3/ErtXV8v
iFWUSB39mu9Yc0GJd/Izef4UsfEqKNWRVajOoi6ahB0OQuNPkk5l4a9KuH4w9wSbeWbBtzXH1C9S
lFm8vBfXGMlG/QkuXUo47UxzX1rF4VTmQpLtYKnOL2M8avWDcwvbszUanzRGJInUod8MqUxceDkZ
xgCzt8gQ7OBioRhA50JndlntrPGT2b3DAKE85kHm0EX4U7HceDaPD5wf/aG9pgHcKccZbjIwda5j
SHulcpbRneUgRSZxlnX4hIKzWIJFN6WKul3TPlxv5h+9r12jcfj2sdqQ5vTgEy0suMAq5ALMkudq
BdgYhIEt5Mu62M/AFgX58ycPZauK8pAScUXKdlhIsrwbF/PA6aWJ4NHtuKopqMeKvGbXQHXRXqIv
K+r5PqqPzyIE8YENTDkgRf6V1kQLMDZciUmwqltpgOpKSLVp07ovDV/I1033vdQbkiS8uJ7u5R2m
o3Y3yMpmKMkLU33uiHtn12RiOx7ynvCBN+GAgG9jsZr3NHa9DuwA4lI4P+eemQXZzy+C4HYi3lkh
9TMNFGB4aoJXybzkgLoAzy0RCJcELWwXpubAU+G+Hp21sVfBs/VB6NZweJpxDaoVd2M8JVxRJO3i
cChZPBEg3eYuT9llIEPDLHxHIEQtMAnVLef6LxpO6HgeqQr01vslk2ch5kKti+IQjm8oSeWRDN/1
OSD5usdqTkzrS219yxL4OeRLFtjlIv5OXBSQbKdaX6faH/ZV65WJzz4/4rqCDujVCaYisag3B0Vy
uo8FjZxcNiUZG+w5SPuSbmydcuwvbzW3dtRhgrV/BChx51Mpd8y7L6pWAh6VBrv/BD/g7LZf292a
Lrv0xaAXsjkgo7ppp0paZLySw4+bWx87Sl335vL65m0i/H/Y0rD7Ov3gd8FIcH/JrpOljKRN3h1S
KDhTxO9Oq0bB+cSyMpKVKcxLC7QzY9ojeU4qR3a6RJlW0szysBFmc/lvl04cse0KL4iUAXf/6Fmr
+aB+EdIsexPesxNnE+ayAyXf3egAazHo/rYLOxUvTTNHpNzER6iV+E+lYN33CcGxE93DqKKFy53y
0AdkTTjNm2EMWNmgifc+hhV3txLQ1+LKj6KgKU7BykMq97zwbXRwOnC/WcqDfdOUN2wTaQQRVvYU
fziD6ijnocDR/fAjv15Y0wCsjOJ7k9p/Cm+eybLjrpqvFz3tAdvAdNv4yAQpU6CXkvS/QeXxW77n
7GCJT8msDuau49wKWRvLGVQjeAr+PaJB5k+Q3Jps+f3FMJ5j4oHWDHp7dUrc+QjtGV0bg8neNBWt
H5716DBU8GaERqowJciTHL2aLvEZGkcq5Ysr6YubqVo+sHETmPjNaICNn/8qmSTmYcYe/wUIgDwG
GYgCwzgAIVST/dohw3QoI6J8A2AJ8PGyRtUCXFLUsAoeVWIcdbj1os0IZ5HGixeyWGO+gZqW9QRw
nDuXQmMttvi6/U9fODLyYvSH8oA6OCm7k7yVGCnY8WJ5D9voIojzosXoOhv51vqFqn9L9L7NKwhj
VSUi0eDY7CtSNGPYjEWvtR44a5Qr1ybZTUgTe3sL+36VgMzrD2fwxwCSKdYdpTfH6OSfSAjXnB/0
Dl442+yuNtUeNDONSoxEeGonz1GFLK18d9BoiTrxiKvqJL6mqnJQSsgs0e8pIPPFqX9sXeB0kb80
AtVRcMd+xd5nXvbwOh/CP99kpWBb3W8v70KYlJ6x/WePVk4g+a4RY//ymzTedJ7KMw2/Aq/vBayT
2uiQt2wapECl2HlDZvQZDMLF1egRk4lWscj6ylK0ds/aOMbzQkVN+PThuXnMdpMd5g9DBD9ngXaU
QFDyGRw6B37jcYLlJ1UjplAzaisftFAfbkM/NcYbNOfCPJJe+Fr8RPijlDgGZeWtbrqxhv7DB36g
dLZf8hf5ivrepYuH1Zp9Ic56j+c3CmiYSFC6ijl9evE99O+WYsyRLapifs5ywIkNtLVtJhe+C2IC
v38+2py0IdpsZuCVCskdAS690jqx2h+FRyuhS38fXM3IisT0s8psRxrDLQL/1tNup6n2jgoKJUtP
Rpc/qE0R6dCqelo7ARMpCzhhmNwjREzvkH3y4tzn8eTAn5mD2c/RzUNxprMDxtx5boQUsHAGFZsM
XQdbBl9WQJlC2s5ZgJt2PdGe00Cyg097+Oh2Iumtu7O1/WIF8hAWVb4BG+z2e8jOk3yHFz+/9TAb
R64a6oGp6bfEMGJl9POs0Jo3NG1Qn3sGPjluISiqtA7kIJXGvu+MqEKB72KNDbrEJkApuej3Z4+X
5gsQI8z/9Inj7hDgNiW1LMR3BFCe/Z0plIsNP1RKjnHMl3h1hXq4r2nVondjtQBe2ghX/Y3kY9GV
o5AHtRixU6sQZeEUfUqnd6IP9qyUEXE8ixdNCeTGA72zCYJhLjBOfKeJXwaKqhcLBZnVFmJpfdTF
fUO7Lttdv9zia8YUPJPnpBlmNmOu2TRQU2ymijeAE0RnnegLt7xEJl2BoQlKPDqasmry7UWKSdS2
oP9Okn5z0SQuh9uw8Vq6rQCeFK9ElDfgqIfjKAYxKV8qXeTF3t0SvzGvemUT/a9t5gDWwpzvJVk5
9BQBl76aFbjajEaId91tYAv0wDq38dGo/9QWR7E/8P86CYiK340YmlDMwHJbYRm713KxePH5k2fm
ViVFWyEtRgPeMEp4wCLlQ9p7A5duIoqpkfpdTJ1/yS1EsD4nRsg2xE6le4cZLQkmOwZy7Iiz0SW8
JMI/Hp38XoGnFa6BnBpOSIjNYLLGO9UYaoRjgGW8FpmZFKjXCq1c+X7QM7Zggn+txkn31dxnNtjN
/oLKwFCxs8bfLIBigcAuzvZOZuMFFD21as9SXj3so2fRdLwgqGuoEnaS8v6qKuyzsDg4OTlf91aG
hU6qFrOm9a7JLiZ0UpWAwCgW+wMYmuCTt1CN87PGdQYtrrNbQma3Rh0FhA/Xzs3k3vgeB3MyaatT
ixGH7TlflltAFGHRWOajwaVzh7TBiqDL5svbgCpqkU/sAGkgSsuMeq76RgAzCcLlKulP14DMg8Zp
uClYf9xUZMYGxEeZ24wfYGL5gXuOXeVzkZ0mP30m9l5qvpehn8I/QirrdSpboKpgsKMqa7RwQ+nF
hSvSciVkXDTEYRWb40rjzMrZu9i/VaDhLRk1gRWXhBojsr4CX7hA+D6aLWlWyOjaEmJAtaJpLGjA
TINDH/0ulHlU0DY5HIGvtIgrjTJRyUqD1KUmYisQ7iymoamWavjpr51f3f0oZh8clzgrPoeueM+n
BML3JPDmq13HpO6W3T9buJDmV3xTkDAt3ncB0tDj1SvXC2n5/wBbXmIEq1XD8dJpFIypwKcKAiEu
cmxvXyNm2pjbRLtYlSjKTFZRWyFLoXAS+YBidbsnJ/YOBKSfs7wJve7jSbgjtr+MstoKkOxrVWjY
uGL7LXRpC7Z3KkV1YZZor++hzsdveRkoMU89bcDNGgSz7yi/4InGjeOcc5/TdmKDSVJSBcc35/YF
rYgvzd6iq10IwFDER62Jbo6SpR+8BEvCYbdc+3nNq7L3H5SWOMQBfF3gQw6cOH+lbmtUXl8TysCe
A5xy5w7v9d2AihyPi4/mFBhxser2G7uYXIOXPbAyI5n3RCAwVAU+zOwco5vCkdjmJ2L/QcHbqYZT
R8THAS/bEyXT4CYwxFItzZLWfvY1Rl3IvRHw8LcB3Rj60/nvhwRYJaaaFUI61NDGR7lNQWkziyMl
QVIAS97VvPD5Mxj36NGTazCJezPqD5SqbPHH7OmvEThmRhPtSDr5B6hY68L/XbYzFP4ptb33jtsY
Qj3QxEY8Ahos+MiiD3Ig30jR6MUiUG7lzymNi+jAjWh5k3bAk5D5dcQR926YsticNHh3saoCDffC
itFmczBXl1+aMooM3Y7I0MaaigaEYz5XpLh3TvMl7DTw001pRdqL0x5jfO7SY2jDK7jR/s7ApDR0
PIUYn6CWNVDCtqOepQ8lELueJBmeQPmBfr4gUQEsZWSOchcpcyep8QM8JG4XVF2KpSb25pHi+V7R
eotmj8Ai6IEJRn9nSjRxIAFjMyqyCVX56xwblPc7n8ZNhZh4dBsYMA5WL+76iruOl//RQiw8gb90
8x+B1lUx+RgPI4hHmJuk/kDpzzPJxum91EbBmPCMvs6yf0kcCIxietPnbjlZifrocFIBvWhWu9fG
eL1KNdkBbLVRSjgr9emJvgws2L0l2SNYxiyA1U/wtC8Y4aRzhmWuG63B2kBH6HA7r+Gha+HwT4qE
LHhDflsE7UrCcxOw3e3TbeB2duYWZ6zNcJuimcUYDPnsnud/LaVkWYiDH/5MsUB7hXU2mg++YAs+
ugNGXizcQ5tdPSEKXchk+5FVimf9oIYjVTwOIE6xvPbaJ5L2omH/RI9wNN/8iogSaR1oJZ4rRDcP
qoyTM+TcdXFWKvd0tHOrymEpt1WpZTQZiwccxMJ0jq18IsRj0FY3MfXefQ2H/LY+Lm4ovhYzNgaN
ZgW/jYi1mQckvd+u7/dgmd9Ff6l3Nsq4mApBuQLVNG85ZPMOjFpw0xr3duZSaTzLvuNXfGbyraMO
DvIk9neZBNozBcYg/rn4QQZmxuOI4gIfZw4zLX/mnDWPc43cekG4wrcKvtM50HmxeGwuL1LBWxDw
fjakjAd2QPxK+6tpflmARdxvj1mBwVB5VVxQxkajbK7aUJMh3vyKnOMc9iI0phCUbPojBD+HzuJz
p/47cqdsjz7ZdXrBtaw53fQdF0DxUq5POnKCcFOe1HZVumWJDV4s6Y7mBVPB6Bvh213pKLmKzpZz
YWqTKwgREzUBJhvv60q7RqVWEZjozcuU+Hiaw5iC/AVOS8nLdpSKHZT8dorVlUVMc++HOFaUT5z8
hx/qvHglVb543Nj4YAdZnJqMTynsii80wSBC+J3++zsDY16c8ZI66z+6vpzCIfd5Yls9dzm12FS3
7C9IdpXMfWYhYSW/XRkEx52FaN7mhL4HLBGDFmjl59c6ykyn287QccpHyfU/DwgjplFGP4AvNFOP
6kbNmrmEwd3xLPv8DZxDMT+mY30QIw0Owjuii3pUl7Wa8RKvCg7Svhk6fK30qPlm0ackAl3N7svy
hifj+9n29lsL0DtHUbFg8ZbMZ2D0GOF3KeYa0m2qtUjJICOOpvX7gz2KBeiAW8BU2Dj45pQSOPqD
bmBW7h+t7Nhx1p4tJEBe/Ff+poqewbPmevFJS2aFK/UCtMQsJkyLoZnCmynYxmQ0jnponntUZ1X1
cTwoUERUloQQX08HMA3N3eCrtxRUEhz/fE3BjR7+XFdqycWGRgnrXbySSPRz3M4Oi8oy0c94w0Lr
iZV8vA1gTI+EX/NOxqhNKBcYxTCU+0ebWx0ylb59TEl/2UJLt7VjHdSGODbPOSM1BpLUaVd7Qbeb
1eGhxxvVzNaqNzFDH7W7wRf4OUAfQJFyhwppPC45HjGONt/HsKniLiIKRdiqXCagxLb/dqV3PKUo
FJgFTeDz1/21GPB9mlkVZNIVz4As+Nrq5KGDGI8ErscQIiNSmUcO1xYVGougQnltU/a/NM/J8Ng+
d2TIGkuB+V7LpxRe22E6nrn8AiwW4GTMPlb5Tgg4o6VtJspdQH+7B5pCDI8L2C6KtCwU2P6o3v50
ZajCZ0T+A8NjH8Ns/mguJZ9wjUw4Wv9+VWe35jS3aI26m8lj4NH1G/FoLfFU7sTjqBEWqcRET5B2
Pl+1KTqOxLjQsfgCcffyy5N3jWLXGzr1wJBkyNQ7KE32tGwgGemgAEQa3QylQDL5IrU+irK7ZJ8b
9l6QIiIwEILJZ6qpbgXXJFujkF9ooBP6bzMLDTInjwtY2Kh7WFFyLJPurKT265P6yyyyQpjedG3O
WJXquE89o9pFe1S0D9tZqFO2T3hb/3jGCdd1aFGv1IgfcOUJReQ3eiNrugCXgZG+uTUvS3PSiVio
S6TAiMAwO4jEj+mDnN44C3VFrT/8MEeNUov3I4i7huDZFv/28TJGpP7Km93aBkhdHogqQ5YfS8Pa
qbUbrJ6XGsFhEVnSBBPDiVU8xGKQ4Eul8czEk7uaazV9082g+nqrDj/FMmjiMP2dcc8nkty0L3qB
QuI5WGqIlfGY5BHzwgAXie7UDUxJtEHuKAa5WDJKAYtbB9o82bLSzQcHSuvX2JJPIdcwtcc7hKXC
TEuw6ajieWceNoVFb3vNhQPvETjXWcv3mEYdgZEFOhB3m2R/iWSd4tTrQ/NeWT9rGSXv69Mmbk3c
6yhsgWrGZ4ToW2nYBEZEk1uGUddgVyoJUYdaPaUGacbLvBSUtfMpdaAQjRX+wS9UmQr3nujaZOcr
LStlioIJUIcCAdJTX9LzctIP+vxDLZFvqczZHVSgNhf4m5fBg4WzZ6UkVya1fGkjGKHNcwA+3ErF
UJHmuqhHnBP4oYjmeE+HX6H7iNnt56ytWwXzc8xw+8Tls7s+iD9RTsompvAkXb3KviGGjxx6lDrW
S6unsPPZpjfbLYPiW7POH7/wBtWBJFDGzWcg0/tzyQ0KDqwlbRlbSpM4N5kXmBJENOYkCku4jYf/
33D22BxP+0rYxON3LIm6LbSL3LAr8ZH90xa8zIHFEeEQh5mpoJzSW/5GiT4oS86RZ0B7eTst7/+q
bzMacxyZCy6bnjSYhLQxHBSMoba0S/8d8CGOXGe9aL3f22OZgifzP6zFDEbbGDZmSzq0a1lrM9QI
/dxTAj99Y++hAOR8i9gVVLoSOaVZC8W3lJ3g5Aj7D+VdxqeNpiMrFQ9HjFfFs5ADGDcQsWVPdYTl
c4glZfesbCUjh2P12Jd1IVh6iVvrkKPTofDyctl3xPlSJJMwd2aKPK2xvzQmXB8VYg5E+PIw9tOL
NIiAtJPOCi5AI7bkU0QfED3C7hQOyRLZxi7YP32PLReKGKjA5G57iWsAU2InZQ5m5gPQZaPwxURD
PjzwNi3OemAHTArSGtUYXGfIz+MFw1jGQ60KVJ0rYTauMiDagmZTqU7X/IyrpJU8gy/KXxznSbO5
ftHsVvKSKXHZ7oCQqh+QyX7Ni2w6l5Stv3i2MtfEzGLfjLq0cT39SYcPTFPmGVlDGJpm3xAspNcd
9m4XX+vsg97jUlgQAo9P0GXhtGT+1/wU3bKuVYT0o/Ek9+69W1FesfPVDY8QNL4v8wgup/ZzIRb7
qV3yAPed0r6+FMpHFuuDtDARnXIFRKFZE5U79u3jnH+evwZSdZWiBg6PTbi6ZicIVaYNjpAaKb+x
a1gDxHcmfys2j7t22cHIktX/raoe8l9ZaIhwD7r3RcNFgZ74C1HGrZQG2/0v8kiZ8nYYyHt+Fqdz
Ym7pUVQSa5u52vpnFtcWtEm8geAsipePY1ohz+efwFQ+LMTtl/fQsv+gF2a2+ixPxSGjEJ7ln5sF
0xig3IxdRgXzjDn5R/eBqBWxRvJhaarBLObTQEdvqFC4D3Pj+dJIuL2etGIGC6kttf1TXNc4SXBX
BFK8GLBrTG03hIUFHqulZdxkjWaN1GQ8BEBNSPlgMv46Y3Kwj3yHp75H5URSA6A/+/luktRD0dDN
SGnh093/blXMG/iFYmPBBUCLyiD6YNCW2EkMpypvi3zXEAEGkNTZZxcKiu2nvTwXf+GCQYQnelS4
Ib0nDkMWZhi1dwBDUxrAS8MoM598S/K3LYQ4r25aYRAP9dAIOt+EPRIOMxgBdlwXL1S1TEFVMQF0
DylHH+GDaPFt0BtttCy//BDWop1I2tuDDTdH8iZdAz+gICiK+faU0cSDwPQCSRXQerKMfAVFUYvy
xdgF2yHFqbNvSlpr0+k3T9ZBBeZIN7kUGXJjGnTf0NxBhVeE3G06ciCBELhPPNlCtLv+Ncy4DlHb
E/p+iGf284Fpdllu7AbsYbmfdn4OFb/goE2CJ0QAb8qlPHDgvd5gi3h1wTDYqVSSd/zJM3J1pUzA
yX/Fsd3Wf+8y63hnKwOGJgr4U4mcWlbo+mkIQ4UVt/38Npfwz0jDsa4cs/DfGZDuFiuUmqvael9Q
/dlE7E6H+rToSKjqw1PAqzbM1uXO/PjOceK/Lwwqo9oqG4/Ashr7CcMW+DYPeb2zrMUHByZk2kml
4lUxr+wSQHBAmYGVp7eiewSoNBCliSOVqPEuz0PDvKuETEm9p/GzZfVir6zbrVrffcRJh+qd4FNX
MKbQGxoS9+nl5f+DXyOLe6GcsxAnMxISvURxytfxaEUZGcyfrzuJazfiRjG1pAC0A2hPjoF/AEKG
uITAjGiAC6ybaIOVPvYqzeiwMLA5FUlJUHzJVtwkMUPttvwkgue0bSgg7wbOM+Py9s/HHDaLVd5N
Jv3w5Wn/vNKuSMP2eu7lZcpNIz1xB/VBwHN9zg5xfv92KKrROcNMQEgymzIcoomLd02HAOcx1m8M
ycFMwgzZ1w/Gw+2Ppbm0029tvqGFWTS8AmpRNJtvdW1FsLXz1G8xY6ucr+wT6rht6bqbqByROh+o
ljrRwCgAD6hQYGrg1fhcFrb9eFyogfq7FDFRGtTmLNqcp8CqBIaAd9f6EjVZgIDaCWEO8brg1yTs
7s7YiEhxSmz18POUQPcGJx4SWoq1RVMyVp7l0cVRc20jszcgyIDvzF2DgCuVe828avfAbVRZvbcW
kWH+tWAdCtyfIXN2JfRiBkqLkXergeJL6pp6UI+hwou6pjhMDl6pDv+bRs/hg1IWVSwPT1T+XmR0
vQd0vSljsIgpCrpT/5pdVqT48dmtm6XWV/S7ZfEWDShvfFXQhFpjijSo4iimkYf8U6ynOBz3R7nX
g5PVI8eR18m53OXMgBRj49S8iyKcmnEwJ/qDUqWhV3oNRx2Z92T7FB6Qlc2jt3M0vJ+fM5yr4QVW
8dgwu5Pi3OJKgxXAikFCePUbW89ogK4SRaEdbZ+SUwHv8dDeaKYJo+5PWq3kStKQzZ7400T0J3P+
bfkoqQm4HMllGOkGnJ9aoInurY+mTOenCjDiKHkMUI6MCPhFdNuK3oIE7vIys2Ij9gHwerVMR/sU
xnRNx9ymH+8sEID0+f3nMGRycnGB8uzX3iUjjyJKyWXoWtHHrgIfmPs3Sq/+A2OGH4reqdAaZymT
UobIVmi1xo57IgLSx3bkLl0SaBtN7QQ395dFT1WTwunGh/xnsa+XPhZ0XQGgMzuaL4/gU66DsLCE
KyvjscNSjEwwMWOC5+vGUxtZupaq6Ftl1+ALFxqNdGyt85I2DN4z6jqOCzC7zU4QUbka2yP2Y3HQ
djGXqmBlYaq+dAlSTNYe5bpHi3aOAyszpZs9y8cmkwLMuYEWN1ecY0D/YRitK57PE/eCrCZZF/Hz
yzPJ+ZsS3LY5s+yYzN895Relvyv1g0OWy+1ZrhXEEZTbzddrHGByDogWxT5y8rBiYBPiuNNCDpZK
d94ITnomAgRIETCIeLrpYCMBxuZ5KP9GP2jJ14DoHDdWw5SXoknW3FjF8awkKw3YuAFpjBHCa/Lr
RyOLZLX9dv9bmitTkRQjUhOdP4qaYg4w8GkTjP3lFFv56xtYqSAVsKuGiD5e8UdlVE97c9ArggJ7
g+mvsESrPVlMzRwg+gLbBB7+P27w+6Dhd0CLSLbBmrpw4UMW2tJcM7FnZdicM8BC2YeborSQSg1M
/wSdNcVd0T0xnCY9ApW5cq6FBlg1oG6wf5tEzHjAfQpbvV4hFUaCkhi79M1h07Qqlmth7YOaNF+E
ttbrntdz/2ShkSClOVoNZRt8lGtvqii+na0nEU08ZvcLapsWhvg09VNLSQHoF6vAp2mo2qdw+eVw
QX8fJ7T7Lsr7JlUrvs9g4Yx2vNbajja51uEAiM9PNVEWkGlLZlmMYW5jg984YlThgKHn0s5VZ9q7
om9MIKE27L9G6GVA/NI1VUJQ1OzDkR5Gl3yu1VMp9tH6AWqbYblyvpUmEPnJbDZaH0CFJpc6FpFR
aWvm7Qh291KKanBMDbFfaVft9NIrcYsz3sUuJ9lyjI4t+WP54J9nbF5e9zT5RJs1cGzToElIDx1E
YTVpwS0l36BERHEX/H8a6XPoiTwkkrKVrGcs2bwMo0JGQUsFIeMj1SNBAstJqkDMH3oKJi6LUnk6
AmZXgYM/DsHkRicvE/OlxnPyHiKO/cWPiUYFiYqMGKIfFlHhjV3ft6ECxCpgk9HazHzZRZvc5u3i
PFIKB1VuTBfy9ufhkbDqDZqtNqHQDmIRgmL7CXunWyyWPSOh82l3uRqp2S9gqFl6829y6xYPKA9B
cJtTwOU5z57RTzASGPfElSRJXfMzpPrCTiISMePyONjbo+S9mo6lr6pMW64WXzU+12DLwALSguE+
LKL5tMcuj+mU9qpGa3sKnxY8l1EFiG1OfgyHo9vTifhMqvhmN0jJAnL7pcKaM1kVvoAE10+HMaAB
n3jOeG4IDagkYKwyvXwTy1cNViUzc1GcJ7ER/tU/O7Dfy3jeBLOQsXH8sPr1Q1QdjPgq8gKHt35B
fc7NkHVI03rTo2qrMk7xAXH49NqzK7lI+Lu/eMMtdjD/yW4b1T2C1u5yJbCh25Jvo7f9EaSaFDIO
v2298c0O2ImX/jIbpAsFHOQSRE1bWfeenpQggwsbD/HrjBt1M3FDg8f5UyRUKf2DoirO3uFzhpxa
iPqp/xH9KLWoKvFZG/4HcNCv25yEsWhqhUbvBYE7uZqpDIBxuQ0PE0G0c3tPCoswLF2Ca94yLdYu
F6pgdYa2HSemPw6txYCR8rGKLGk7qJbTJZ+Ew2aEFrbK1G4lnIIAOCKWapQpw/EXTamo4ELZBKpw
qOCV3bUZ2V3X/vWRmeIuidPpx2IMpJA3dccjoLxNjGtjhOKlM/1hExy+IxY6mXdVqqdichjSEAVo
Pt+iYgxKQ+O0LqRUlLDDtQ73VZ4LvE0aArnG5d71/4+6uYHMMfgWIkW85tuUlLzN46jK9ZrJNaYY
UPy8KLRhxvWjszt+GLUL/B7rvqJ5G6OfQt4mJTohK1jhn9f45V037CjOr46pScvvuxEZ/S+Yq5Mx
+3OeknQbDjvvm8+KAjb8SxzUYWPf20ALfnqZmc+5Du2jtv11hJ1BpCly4+bbQv/3J5eLQO7TqcJa
HbNrYvwywfZwXTL9sQmSXya7Dim+6/DRkTL+6V0ZRPT14DEN64UuUNNgIjVA/jSi4jFqIcmaobhd
1TguQ9dRfNX2Ju3UkvkSt3N9AbPMIdU+ZFexeN35m6JRGmTCH9rkawnrWBA4bEHgBVqk7q6v0gH7
SzyCYP+RANKV+zQgLieICUnM1NBQBjKPtlUUxh03HFEugD67a1RjqwZaknj7igrfEmBohXBjsDq9
b0F4TXHvojzwi37FmiZaJF+JdQhSzYWqqMLX0FkKAukSzs4Lv4gGs59ft9loNC0Kbz97vJTctjus
CWUb018FXiSLt5bf22NN0LBtagwkfpDPXO3rvKV+k9BIer03nRygOFpoUtlJ/WoY56+SGJjS7ZlU
NBkv5wCJQBjVXMLFyCNL15HYkHY2TAX8fniC9yxiQgAHbp7PdF9WipHbq3pUmegYUNycUDxU36gc
lrE28Ps1wTlD+xRMBiTC+/UsXZn98qjPNqP9rg5wVNS9xJhU12jSBNOiO5AXC3FvtznhoYm+TOfn
LUJBa6R18OW33bKXXtdhr1IM+Jg2fYIvOnxHfKuDOIKMezmgM7C+gKYOOGbEQB16Axc59motn3ME
oTkLvgurO0sdELxpP8myhPpZErIudd792pqy/95YM7+1WO9kBTmmKqmAMJcdvIAtrjBLFVXYDhkF
hNvYjiSWAZ87TfSs/o166D5oYjk/ZjuLbU3p7f97pz3A8/nfOXG+7m2LZlnLGGVNred97mYXGrHK
rDeK6O3RknatFDSAcEe8zVzCGfNijOi25io+HstreJgz/465HoYTfFeqy+O1nSNL8LxXzzfGuOls
IS4/M1L9WYNnOnUNuFw16iFxYPVNNneItkqTKVpzY04m3gwtnXJv8TUNHatp9QGUPPx5RX3oUMW0
Lv3vAQIca0AidiO9yR2Z6B7MwoVPztcMRMr8u1jzESTO6R5A9f6l09twpwVZDrIlMcA7Jzetda2S
RaZ8ALcpSt48cEgla5tawle3au6j8lUlSE4CED2kmMioCLQPhL24Pddzr11NfV7Ty4/EdizQ21Hb
NDFB21mwh2paGjnGUwMB2a+pH/ktTMAmsixHaLNU5kEujy3h82PEegppP+3YYofufKDWNZ03tpOp
acLaWMNd3JOWZQskxEKaO/pDp8PJfVjCnT2X5TSC3GlX3n3w0eVSCbQAu7l4gPkenzptJOXpmzIR
aP1Hvbb/7GPje0p7SAPMA1bh+VE3a4JeGxVrB+FSYWgJ+HEG1s5BYeCNH9IR18ojX9FkmOK3MMDS
pbvZbO8QL8cNSPkbfL2E/LKhqfBctz/jk8sCXif8HnXZDxbpW2tvq/Xs6hpGhcTj30kPXvn3wKec
acRJo0gdBq6jfz8DNTMHES5trvb+RekUq9/l+BSPt/uJLeoxDAZjDH4qn0BPgnvfVB0p9IjX4lw8
g48Yx07q7Logdo2DV8486E6yG0Oz+xmqcp8zQ8ys0NSS7iX+UUMr3uiKjqgZVe15uRjl6WTnGN1p
hHnt7zIqEsL5A0uaJIsjzTqqPRdNhfuOreK4oiRLs4kGsVC+n9bc0LrSyZ71JEO9xg4aw2LGaKVw
abgm5vON3IrVf0gChvHo3rGYts5HZ3Sx2nhgXrWnWXeEJ5Jmg+JWUFUUBz671hRPLJWL9YeIXSLM
rbGihtbU2yuZ4liL9+rgEEqEIxnYY8Y6Y5BvnYFj0Sc8DzzF+QpGTwobEVWfL/5vB/kiVswsnWrw
66Yxc2wubsCpTtRsYuVnamUfD5wut9s3tkbqzv/zwmtwOGNUTuxR2/7HPlpIjRpkAfBvP0yPmj6j
vq48KTxWB6+ZjHkGT02ccbpTupB06TWyhnhMreA3BSxpMUtgCLDRdMPY0OFqr+8Q5kKdSUUNdRBi
MutEmpCZ4SOb93xwUSokM3YYuYUptee7n25B6oJnp7iXnt7+FriG5yelbdWeE0WZLUC26cS1x9UH
CsUVSR+wmRYBGqgI/GTubluh/aKtmUgxgs9OJ9mNskgBsdXTiLJFQ2K9DbPZk+87Zjz8e8r5xGm6
sg7my1ij7NmRof1DPIEA0kMl0ku7SxRMa739lojK0cshMsOVHORRwZXI+SNmkMn01MU7lOJKNU3d
rKIDL0XbqAOw+MTq8trUnGo8E2skOTLwWXdJFN1SUVpNWvYC4Hbexmi8rzi5/F+NWIpfjmF+IsYX
c/ZaErmdOC8XxEri2Gax+6owTLOt38LAh2jWb7Rfqu55b67h1b+VYT4o+s6SY6ax7E9cM5NNOojC
SzXbRRNcMfEnqJJyBLmm2wlC5FaeA+sWmM6VP8I7ooaGHd+hGePr6GoiUjV2MDIXcTdy+b3r1WJc
lbuIV1646fkyCaEQLjjVFD8Eplh2Gy00Td3edjfg3nKPF/L15SSFokmy3K53dGn+UnaXs8FU06K4
eHrDQF7X5rLKh468D7E1+6H3LOC1uKyMh/YUa2xbh4yr0g9mX3tYFMbMZPH1dk+4z6nYlfdcbWoA
wVxp4pgVAvusp9BJhNjWxXKOxvn/9BK/w8t7J3dFqrzSWwvyZJypNi8U72QDKWuTTuFBaA2ep/DJ
DTicYlWYUEVpZ5+boR0GNk1XvYs27b7RwxDu99xKNaGzQnPcFcTcYgJO7zvSEJk/W8b4Xg6FZlXA
u0YKR0zFbbSlcqbv4cTmrrLhfz/ysfyzsl2LEpndY9fFpHAHnSe5vCW+bNiadbmeC+DmNJ5NWmPs
SQo7SQj6vwKaDi99ozxivUqqZqB+PNyBMcSc3AMoEk0UFItNi0wXoOw2JMzZxoVTZnrlZamIXPXB
cSWTN9rXonSJyDBeoDTPOWu7/QMoec1x2C5Vm7nk+bj1KynPQhX/FbbqZ/m5cDlH+no4xFVcU0f/
zX4iFSdb8qdtimqwvB7TnKYMFUbH27Vwiy0736QkzBaXKa3SefhgUu8IqzxMD7iNczZ+6iFjxLOz
zhqCydPAj+4LzVoG94PocOE0qXo2vh/8+i4gg/1XLn9HnWXcwjbL2CMit9musU3SSf4Nr/w7ri3i
xgsS6Q1D49/gGp5AxzcyBKOpY6S6gBnMQc0TKjRxpsjnwwo8Z4PhgM3vLl/FbffXJ5tzvzO42c29
Gbk6qOX0oid3FuaunnZHqzLKbGtN6u5caY3uNkQNdQqZfPm/A5RkS0PyX1GkbrT2bGvg70gw7Qi5
80b1cmwlzHVEezr7xBitTXjgyISR5QN2ISvJkEWTWqON3VZOSrp+kJ5oD1SyNgfeBR3V5dD8b7hc
7100njZ1rY5rNuTHVkQ4StGpiavukViSR2bUZdybZetBGaHEg8fHW6sU8k7LrQ+/ciql1mpyDznC
wTrE2CL/Lu1aSiCV0ibagUySZ4/3IcbOYW+DR5TsDY1UQCOjfUslxxA/7WmeWwwMxtpg0DWvAOh2
AOfUqKOKCaXeLxqkHJYLbIfxC3yivtAFXiiropfAqAXtBnCvyhMwtbJaNRKZkefSTxVUrUq0ehOw
UjdgKkdjhtLPzquwzR4WSNYWR+aO9lqQ0Tr8BaUuncDXRKiXg47ImyJqPQFCaz+RQIe9DF2evjvc
FBNozROX7FUFUBjy86TPlQwk01/3UQSMXuumfSOUc/mD0vAFzORIA0OH5ImNeUSi9xz+VVL85kzM
kRJtna07b3i40l6/vb8wKWv2NNiNUyFfcygg9pQ74780ZLRGwxMngSNH2abkeWcgF9IR0zI7YZD7
FRoMXQkRsgfn0eU2XOZ/L0CqHWfgqtXALUVgYNwmw+EXgDGbXHojzkKVS0t9IDl9V67/j4BVtYc5
OhIekpFNduoeBCrePjaCZ0cCqmEtEewDTpnbVEtVGhp+yA6xUDcTVqmDJCSnIqCV5YsVzUdgHeaM
/ms9aWw+w2bX6PcqygHcBT+fkR1T8aq8XTyiGTQZFCvMziw26IEHeSxvn4xZU9RsnbjmhoNXrR9o
NpApy2htZSU0eHrSNc0jktzhb6QA7zuA+qieYYj7HGHZtDQ5YT6JFJS2bzcf1HT1R9am2gZck0Bm
EF1hTvmxtQUmysYGRtWww8XvqbSQIXuV2pznZEGwBoemYEOHOwxW8Ab9QiKPgEi0F4uQXXBb2oSx
XOJT1DeWjRwzlUsiwN7/iX5ApXzgJqJ7SrlxwZd3Pku39TlvMg0T2qH3hisn4gYwfnOktRhKVc8I
26Tg2hnhLNCGBM0mLkPomuhhIaVaPfpwoRI8G7J+hVyZ4+Rwcgg+2JoakTmUZ3fBlg+D5ObWEiWu
Z6i2JlV4GXYwNKzPLD3XNlxscnULzVI0561NBvqKaR+uDIXZq9pAg03yHKm5Emh7RrSWCMJ+5H0G
KkbGK67lcOioeJb+FDSDJO+f8o5xkPCJrVrg+YHK89341eDuO8Nb3Akvz1zu51OXQmh/5fRe6kNN
4Wc+cXiqdVrjZaajutnKSffJNq4QTkvtc3Sk8LzWkPRVLN2dElh9ryZp8IC/WI493lxvKvNXbKl8
wn2DWuDzTaqWOUV4b8W6C7b9R6VuWN5Upvqmbg2pD3drpZGg5RiKXvAlRh6duTdJV/6TdlWqei3X
HweLQFu4MTk5jG0XMeeebi3pX78ejnPqc3QhCFhWgIfOUlG+q5XHKpjw7HHzvSyO3VBSXehXsNFY
a9NjPTS+umD0eOyhcoCkLucexLvKKptJuBnFr1P+bAkPQHJGuyEhYqcLP/TRtPFeQv3VTyRrg+DX
+45Q9OaKuCUKwJc3MMaAKkbkY6c3SSgCmHpW1PJb6jlz7CL8lvMJ3M9LY9pSeoAwW45B/gxK+fT4
6CtBhXqhDamMxniytoTUpd6aemB9hUff8iin8dBgoOTcx/fNiBQdRGaCOIZ5/ypjkmcoe/CkU09W
p+N2SCfMPrxSI5ki1UGEr9XzoR6SIT1mHdRpnSCrQSdOiL4IDq6zo691HSDeLwGrVdZZC5Y2QTSS
jVuIkXW4QGeMqWLhd3Ze2VSaEjahbR6e43CG5m1N+FDvyalx3OMSxjXIkx6Or6MfO+nMJMhS0gTs
JNWZxK7/keQ7rD0kZ3lL9tnF+7B8fVNNaBrUTvJ/TcHpfLNhlSy5Tg+d6Ol19Vrmliw1EvAYioVB
gfmcxyVVOlah1Oga1CxWl6efDsKNTCaLUezIuxVRmy+dG/r5rhuhpo1AGKA7q+4TCvYBLPUHkPOL
wktjDvlWMfF5Xp5flmRi3vinkMy/ZGwoFI0zo0R+ctiwbOLDYRXOTOxh/QCKBGN9QY0ayVkqF3vk
lO7Sz/keGvlzDWMnLelzwT10AGdv3KKeSntDAGdJHLr6MhvGMv3poP+LAqolD8G6YPp679aplu91
x0nknciRA7pobIOcQFiXzP4nYvLMJJY6ZJI4T5vfUw0iULqDv6GVCuQ9ydEeYO/FBZKXnB6DTo85
5nAT1OoQsuEl0LFhtnHxqOMKOfC1TFM+kw3XiftzUXppHBl5+8SEsEyAnsq8G9897VXBPM/cw0d0
VEFuBSG/ps2Yl8zzkXBiTk0wAGNT9tals9vtcCndPs+apR73fjMV9nMdHKGLbwMToCPxkPdG7sFo
9eFLfeiZS04GHhuMLvLoIEGRh3XtHhdpgdBK3hkLbNVK5uw6cLkcH9arAI9gxI4yY61rIIc4bB+d
O2oEqtVcMpl27tYGNCyszGUmsLy0gVYgkd8PwoXFhJ86zMWNm1Ay3qIMrCVwVZrnTP6TFPK02RQg
EoR2t/pMnl8VytfqpB7gg5Vtz06/iPHz82i6OjRRKdH7t7EAYq92t/W5f9ASrsgGM8ni/TSinVu4
p6BrROLip2ipKf3sa0lAHDoh95rqf5aqxv815iGF3WBNFIkISMDj+kixYPQmuuTwFJr0nPuT0PG/
hJSIBT3ZHBX3sE2CPD3PaurSPVzViDUxYQKZy38MF/6+CcqI/p/awN0tI2XwjkbArvVtBHfSu4F3
CCS+aUaB3SbWIN0CKUxgdE6PRK4vEarW8rkf7uwDB7mikM/oCw+9MdpQT0avAUnAoSxlYC2w3Vaz
at5OMcNx8IHC14UuvcVIf8ZADsoykb2aZ1BKz6nwcaOsP0lXXw/CgG9MWEIXEngKHECdILA+PP7L
EJudRvyJ30SZSFm2R5qS8TG5/4MR13cwFKvrmjQUDkDroe4zMcjUhWkxt7W2GkvcHfW0TcHc9DP/
nrfJRKCA4To/FFshEWvbtTNYxymoLNmVdAYQ1Zg+5qjYB/OmNUie8Tt1G1dtFM4peCz9RF1gmvFC
kaImDUtZ4TeUOn9BVH9aTUFNZbIduVx4XBGrtczo7a2nFMKrexh6g3Hb6aQRSVAEMmwbowksX72T
fxoXrQMUGIlHxjofVVQrOv6lrdvbVQ/wBVK3sXtZuKOlwBIVTcWIRPJmlmK3znGGzhzaGHKqExFg
UAykisLeYyXBznDQ2H+EK/+NdC2LrcACOqiyzv0fbsoqaMn7ht4R5SKQaLH/kIQc7JDjKCHB+MTi
jIJOh/khWEtZfWhENrSZkXv4svrEr9hOGHKJ4IOz8kyoMNXdyS3JXOqvvUXpsj3omn+8ykXGTMjZ
2qmt75i/aQtPxyvScEIfHeAIl5C48x7LlBctPCP11t+wgDX/uibE7T3RW7OXI2EZMVzidgy/Wvjy
jvT66uZJ1Y1W19CoFx50LxyT4G1qGnmn1eEX4ixEtmOTekVLkFl1mATNDw1ONYj5JSZP6rREzOoX
1IvCEaFg27C8Hb9UpHYKoY1BIbqD5T6AaLR2CgFFGu5NLP+VggS6rlKzv3tCuNFB/vaMi33Ru2ZL
S8V+HEApPdPvGUzRtV8rkThsUlMIsb2qJxa6mTe4RSBW7sQRgLfywLKoPOOKb5VsIri3H5x2OIjs
CkClxmduW/eDMx+jA4nBODSiY/Sl2zNwWuFOYkwVrDZhqAg0Qf84SRJKl2nljBQlgNmAaBYFVegL
lRL/p7mIbe0BSh0Y83rKtt41YOb69iqBkHFNc/DUCzfh08BGs9qgTO1WxcQD5TUNkMwTNbeYoEv1
97KFm3CcxKDJDkWl61TXdge1DOrV86zAevk/zx47itGNWbomZpl6NH9wJbJ/t/0aCpLyUiwwJb3a
o8h06/HHzfYvhNa1Z71MLJSj5mCATfb+yZjx2SdMqTpxlloGYu8AUUgswXMN8PFER4RH7ZoyPOad
CeWGVjyuZJarrLJ4HV1yotWBivwQkO7SKHECMRr6weOsPjRFPzC0D0HfKdeHXfHLoaZ8RXmZEwfE
ZMJSjrxn4/BYMaW1gUb2v6mL2EqNJEcrWXziyU0qUS8nUYtCwyhWHPZGoXN3Gf9V40zTT0j/8cec
Fm567L7XSNlpchGdyMDGQBWrWoolanLmcvB4Vt35gwdVUM/aUFKNhGBqcrYmsaG0dEeICWnhWG0T
5R3U5Yid0Gjs3sQB7O/wpi6KCIGarvGqQPxQtpAFhK+k0oAreecoXWbEvk4fwD+dtWaIganaNZzM
hznEpLwHaJ6OkNALFF3uMEZdMkmbY4Hp+/ktSvc5D8gOFoeUZi6ya6P+vp0FEV1ArEv7tdL73+qd
TsGSaDXNSlTVWQtexyThDweieEPwznWnJRd0hDALoz3WUh0Fkln10zf4LX0AEOE0kJMn1+KybpRw
Xu25uguxySRG2TVVnWEMup6b8HC6qfU3rj+wJWMb4Ejc4Jh9iTvqz5lxAF7FWMOgTOYtk2npdH3e
mhEHrgwbm4miq3VPK8NtitBkgX9tifUwViZ+iv/IknBWVUR9dtEg3lOBPb/vITmCcO3Rsqx+36Rq
vOuxxqqVhtdaospRQH0C6CP8hGP4LbuLILJbosFFg6w0yQcllZdTcRk9lv2S0okcK+1SIeSjSTDO
1EjSFN5gqJGBturEivp/jHKr8tfWprY2BTiWSOOly90ClJd5q4Nis3lniI/0MXKD7VlUNQRgyjtz
n1R6vyD94xQRhvT0CiNwp5KlNiSK7S+Yi9vL+P0Ha4A7uoXCex/+TYXZAtot9e2BeYemIn8VIJ/P
My/1HZhkZj6BHgkO/nHBLzqAkY2AXeRCuYVal4TyWxMEEYqyxH65aXRpOx4gNGooeLmJ2G4GASfI
v7GZPZuLCeJSFsDzbCXYR8onhcSU/GKKFuZQe/Kaez7j1bEVyiitWHTY6GLSBFqsseQeg7GwGeh9
WtC2nbrr7asOTD1+O2HqM3u6AEltN9bgrRIw6U1RDsag1oXRYCg2wUxJI4z84Dxw5SGRPlEjOQ3M
+k37vmcGfwxy3N57gLzwF/xvYy5+UdwX6fIWeyf7YQYnMAIGzyo8eU35rW3leIGRMVOZOOkzrkS/
4Sm+0ayrRjKfR3LI0obf7no3/vWd9ikiNLOq3iMJh0QFTjgy0XTH5/WrY70LdgGBrnWkthBP/424
uW3Zz9K7ZbKGqeeJirGGwPjEUlMiJnZfFVvUVpHI7a6nwvmWaABwiGF5SN/u3LHT5y6RJVBydgCl
n68jif3tF9fWlMEpXq5o4YQ6SZ4bi0PbC8LeszZFgGHY/Jq9yC3so/0736H4PCG4+guU0Dh5HBFn
W82+mDIdbFHzbj2QyzXf95vrfX5OoJ5VD9JeqMeHzwuANLKiCxcKkKPqnYlAyd0Thzkd7q1iqfFM
4ytCv0ejF2O+tMe18PxGKRD246RbcZAa2BJPCvdlV3/AliVHnxMsel4wYGXfDyfbF+0slciNZ+xi
jCcGknMKpDVptHibCCQdA4NzgPeRB7VkVrotYwThBD7QqlyLf2EHemyNa/RqqQOKs1zZaoEclZ1j
fdN8IB1YYKB0C4Vrc5croMz86JPh7SbvMiHWxVu2wyE6EJs9VMT+y0Ni5jQWX0X9AM44ijj+yQv+
u9dHQi5X3rt34qGF/h3huklrglPIp6Gk6nhK58rLb6JT1w48+bPhxOe11p/otdFeoryRaW0pzkMx
OOpQbV8W0q1LLr0jhiXjCNq0hhwOWVxdBgjmhJcuTjc0+UAovTv+ItL3ia17BvI0XX7jw7ebGWT2
gJghHSktGTKxNds4d62Y8Y65PP6OZz5N53tI6OZ+A/iDGqUaXmOzqEc9EAUEJGqGArvg4eW7+uuZ
MQDgsaT0TsfoRql721s0NzuM+Dhc//SwMBJeQtZ1XxD5BNc47jU3ExCEVnB6sFfkM0coF6Xf6o4R
gi6zOVnYLIZ6iLWrSHqLWVXEDttDRB9hFSXyzIWwg5OM7jVV25csq76uzi4C9XWsKsmmAA/WCzHB
eZ01sn4LKuE0rvJTs58lVOBnfHBy663RUGSKEXUY2bXiRPDzoY88JRqRnRf9HbbgxWSXZuytumV4
WYsVd1D5G84A9fqSZdzfzHAYGpAt86sGakFBVmj68Togz6SAmXOpQMV1wKN3d37wZe7GBvCBqqzJ
XNqa7U/YGpfmz0EM4pV+QeuvwyzVV5KdHqtfDFrdhw4kI3meJKlHMszFyW4NSQSkKwLcEGpJTW45
pw9/ag/K8sDHXCmFbBGczc81AycTL/tSZVksmiv2F/U/Tn0QQe12CDBULuehqSsqAFYNAbKXlnN3
TdRFK03eiGtg6IaJp7Nr06iOd4CE2qj27WtkYgqPcX5saeHKJwZl4a5ZP1h6EDAZr4WKsvTRcc+/
hPBS1gL1/aG/rMUXVkiIC1b2FuaKU3SJcwsgDg2G02FDsWEHyf2JBj3pgUjOrN6K3gAIK6L6Lm25
TsaiwJ9K/MNFRjdqj3CKR0i6skCdim7TMiV6G4qM7bT5n/1rysM/KXZT1Plm+13WQEzVMuHmeJUH
7IREhqFmyH9xAPJMdMB7UbUhGtgy9afIpriafKONj9l9yXOx6tHNLAVHykCUSsGVUgT4hIgYp0Zf
RlY+tZJtlIqaDyP8aEBu2Y+yu2Nh1NDLfkbyrIakBDCip07JUJ3SGQJoFgwRGJsvv9Ji8y0bnYVy
FLpTl/OjPe8XEF13UXJXVXAKd7PjEwuCELBVVciVZ8ZT87POduQuCgPpqHim05P+lU5th4bulydR
ZAdFiZtOgz7zC6SVZM1JcN++MxFwtUW3hIBsGasdBvEuM5xCTSDvhjyVDSW4Npv366+80aS/tCIh
3zKmNoKUlaSNC4QeWsRbWYMwHy0oseJpeUWXBQVPB5mBJkiPyxO2oEQEWf/7rKNs0YEzx81PDoaC
amCHJ4R1l0g03ex6ZIxggrPPprUc0nyY4JynP12VHVMrVkDyYoaw6vG9Qs+7vZz2vnC1qmmvYLmn
x1gMCpMcUwBvbfYLcKcE31Ac+tUF+jJA0lb5WclkRnEoXWXT1FniMlhnEje/pSQq71cqoS2T6kzd
Gba5w6zGLW1DQ476oZR2qd6rPNZ9IJUD85WufDVj2LReR2Kzps0xCDYQBt3YplYflZXtdSOuI5oo
E5Guw5jg20cdozAe5ANXY1GFGMtJehDoDzS2E0TtEFjlo5AZu4YzLzWoaop23Bw09htc+byvMSub
O74Kxy0JarNFAN94ck1H49G5/S9aZyTt6oI7vuTMbXKirDVFB29QC84Q3G3SRsMPDi5a/vkiqPRb
uRdZrHQ3Q0sFNrFE7aIdb92EW+xO7tnkklvtQZFFJaMOwYqMEnvvzMzRSiUghi01FWwT7EKXN05O
OmxFR8tPGnDXHxgPHNoZcl7ILOMwxghqEdv/eliBsca0LErz4x+GL4v2SoxS5iXNlVNGi309Hi2+
7ua60FSEMuBqRv6HqD36bIBWcmF8up9vM2Fu3hRsUEzHc06UhXNCJgrFYaWBwrk3Lrd6g+JwdT9u
cmeQZg9+QU/hj2d8+COG8csVGTXcfaB4SWBukqooNSYr0zhmap+YErTpsUVEmbK+nkyY862WlK5r
ZF+bRnGQDyeUszryrnd/m8SmJDOunXgt18SB+LxBrYJcXZyayB9Nk8pqE5kQRR7fPSlQ+43BtarP
AQhlFWmUy9jHrfMMC9cepH3EnuCiimA/PF6+KgNsNmuv/i3TmqjKGKzcBqPiM01yFJxIingK77AB
qiHCD5+eomjDZtA6kDVNTZa7+qXPp1nKaxEt/7qvYRpwOA7Rc5d2AWa5Q2zxyBJKbHVDtRfN276X
htjpPdFY/l2XoNlQTr4U6YdQ0ud5uDkR2S+wPQhHRsodpjPGc3vnAKSyda//qbjLTSFoTXLX+qBT
5VtMvQi3/OzJVzrnmdaqOdJpTesn3MGnxlwj52OdSU3DYGAzIvZ/c5xfCBkIV5kDSJ2oOoDhw6/R
VhhdSGt8WBfFq8Osi5QL2FIkJ+9rbhlCFEyw9Ub5ytginr1UZQAaHczqMPqayineYi+WjTgEm+rz
liUQSalW2PBhcbfSs5jizG85iM0LXZHukrd+u1DY9iD9OmrCOJiY/SRcqFDEupHYLbBEyt0pjuhg
fU6VdcpCYzC+YuuN4nKDa0V5noUdlsyQmSM58g42lG+LoqsI6Ke1FtS+E+g2+Sew/FdxbW4GFtnS
4nqk4X1FiUXS3s3R1OZEGhpnWyqxUh800DhGkkirwLIuHrsaM5u+HBUWbibuAT77xogmDThW1zDS
+gZ1id7r/h+BCaUTK0Qk9Y0XyAVr+LSnx72VXK/ceEBLgvHT+UNR8beWLg0bfa/ms6cDbiujAm40
jryQ+zfED7ELe3pFbrlGjexCNPpR4NxKf2kpq89KCOau9/4wpk5NYXR6YQoHl3N3L68CCOuEdXt/
qB3tpRC5E4bEXywu5asYLrm+HeLIWlEWifMS+usoXlpMjnFHgcdNCAquIFzif5H59oYAAYaG+IY+
hQZG3CxANeF8r5P/Kc6woX/3QlOXrF8pgK3U/nk2OGaGB+f9995MgemATdQOAUzgYS5gKWIO7cMu
ljwtfE6pjIAEbP0/WNfxK2wZ/AQ3YhtqKrtPXhsyIYXjaMIiaWiUJEE2F76FY5HSTDNn2r8qLjOG
XDtm88ukkBucNGNk8Rt/V8l2apC7W6az6qxTnI/TG9cgz1QVeqZWWpNAuXz8eAhc1DwktOhAu0UH
usJAWfkQnhLCaMY23u1gkWWQyfS2gsp9dkrgdRNROYOXWS8p8U7GmiK5Zc5NyHe7yrVK2vwHXDgP
xh+izjcC3qHtgNxsXvNo9nonRJsf0s3wLB2xzwMADxpejhoBAd7Gc8dd8ghqEG1/GdgcEhJ+QH4G
sEZEpGiTIxxSrhNACvBPX6k/296CoiP0yXq1mIYJz+5OFynp0YekyAuXDWXPTmEhsPynMKBTpTml
dstkQvJn1SHZMvIz0v729BRirPMVmV5zH47yt4Hy1tAJCqncfJ02RQSJ/eaGd8rwhctNQU9bBKX/
Nbi7lE341WUQflYz3VW6vzd0SsA6Y53vdcFMXuWEkuU7CyZ4STDCvMN8HeoFAt60YEYmE4YYFwac
OYMpuFkCBedtuoQ71zAvFlbv6hwTfowWJgB3gXkoyQICDl6WiKAwdxd6FNrbrgi88mJF3oaZ5dh7
qmRQ4x5r3I1QfyWrE7MQAmHwfdwPU+eVL0I2aKjg3z2DsNUPNDsqgsch6UOsBo1rhYaJoGq1d3nn
sz8rep4UGvb3R/ril32MqAy2KojD961qlRTwkgHokim7RQOJsjacuzJDgMEjzGk8IBfBO1zemlAW
ENhE3AB6+B82ufY5GtBEanaw3wya4J98q+1d/j65fp8h53EzEZs5aYb0sq1E3GgCcl8m58R1fn3x
Uqtnzblw2kDAhIRbqEsQ6SNE9nmPmQCKwOdzoQ8iqaE6LlRmJB2wwE6FXoAsElURKDZGVf53Sjcf
IL+XNCmRe0BIZNVZzePXQE7Ew0N9Gbprup/K3jrgrv8ewmv/RsZ/h9wbbDqth40m2mT0IQsD0Asq
phFwFSs2vMJ/kMQz29DK1QPzKVrnTSZjv5bK2IQ9/3jJiuU8KFrI+Wo4Gih7CUKQb/m9lU4DrIoQ
MM1E0D4YKw+PCbEGIkkDOUcD3CXf/L+bV6UOdFLtMTu0eEgxIxkRsR8p/M8zcOX5bHYKAhel5lVW
J0wvAsgS8QUscJrakbPlXQvWYd0jAbLBLRVERlzuJyAIP8IuiiDBolxSLcPs7fSV2YAyJIqtpzta
CMCXdCJlhp3xOXbjzazQmhVhJyH2OJU6YFSImQ4xBCisyn9LhINQiuaUBTfF4ji/1jnkKBR8pw+c
nKxAhOZFlrBR9R/wn0wOFNc6k3I+PMiH5qt1DgFCxoXpMeKuR7UY7wAh+/jGsKhB8Ko9HVxfTEf3
AE9fSdcO5txSaeTEIGsW+8u6bXoDQjVxJFPR6qkN2xTIbBncxBBTl8IIika5HNiT4bwS9c4XaqBj
9Mx+k24JqOpnCnZ8zZjF1PzYshkZrR9KAIWEorxW+XzcdowpiSHxT22w8bMMsDjci1xTJhnXYuMk
Fwsrfr7gZnsUam8vVQQSa6sr+rnc909SDnk7SE4GtczUpKJZbRgWexT7dFGmyvRPZ6nLECcXSwXU
hJbLTeQa4TlmTxispFW1c32ZnOWYaWh4MQamxv6xiUgyI1XfOwDxvu+kabIrtuNHqrv4II6vzDfr
yJqtVzV7fo2jhTkDT6CNMB2h147u5n7te36shjy8dLKiPcWgWxrzpNvGg9BpYsl+7FFXm8ZLAKMx
y4ekxLjAp4BdO/DVBfUniuLliB38mdexdpO0oQcBjxczoIDdPqrE/2ONPxButi9YbwEaSHA/nIdm
Dp52Gp34b7yvdKn6tqwFBLOSPZkWe0I5DSfnpVb2KeaWM3qst5bWtyaWpKqls6MRt/rsrPWmzFmA
suS+m2WgJi9k3JOdoXCQr/X6P7DqdV7Hj61eGd+320/7YPtgcOHNJonpxUUg9XIheYQihPkJobE+
IJV2u8kSqCa1fd9OkbFGt8khCBwyUFhQ1PCnRjPXzyYkeoyEA8SB+ovn49dtT45SA1SytG14j2J6
ddQUQk3h5qyZVDIUi5N38cAMHun2EdbT32f5VpP9oxq7bwrLRI3n2fuAHXDnKCWVn7RcwCQ7RcbN
hGgsg2z8rWcbRoOZ0wAdPdnMiW9fC8XewTAGPzXsYWffS6plJb0Y21d8Wyl9gOgzYAGLC3aFapH5
aGoYxxeiq7N/aCb0tWbKu4TWnnUvOjEaMQO0S0GXupWtIveLt9ZgnO+uXu8A4uc+okg+b37kNlNY
SBlonbCLsXOwXi8meOH38Ac8s/ENJ2Qibp1vBF/jP32b7zl45GA3KUReSgRx7eiQ4LkLSAscW4aO
yZb7RivPFpR3XWJ0u9PVeID3Sqt8F7GYO0JBPsC8C8XdReftIX7s8dGimjNk0psbnVLVz0Qe26na
uAxF6KlD5n0WD69IKAQQ/VPfLjeVKMcFDrbXIksxe/k9aiexpB1yZB31PQfVUx+sidcSOUfAoxOB
ClwknCZ+0vgDn2ZysNAZjC2upW322IWfiW4lSXYZ3xaWF7Hmgo70kg2ilP0alkhKc2fkXHzEtRs/
ctnAuvcp6qpPyHAaYLSH1TKics10i++5wcTUjtXbziH18Z/foFTY7ot3R4mdrl7bThhhER0SWk75
LWFldp2ubjVMKgoYHV9kD1tL9fzi8co+/Jmsi0TU8uBnD9edAdXejYgDdangjXRYrgIJMUd8YqyJ
HSAvTitLcxfXz6+JJYbJj+aQf8dW93a3wfGu2sr6oTince07JDLaMzLH5WDfzadwTSIQkfyOF+pn
OtR3Tojy8lqoOavULddsF19pGXh9y+TI3V/4pMoarfRnLysSpyowHCgrSkIWcjzyHhbtGfLG/b8U
oeI9T8KfpsW88/B6TXZur3h4NGKCi/5IsQeYGWaQR9zDuGmJ0egLkMACuP2hPfoyVtPd6HKpd5cG
pu8oJzKFabUoKpM/XCf1vAstr1UwKmKVlSf1pnpPaGurE9uvnIGFZ8RzD8KcVamD9XFYZ+xTHLi4
oDVwqrkEGUiHkudmZReOq3pA0e/N49TWd+yhcvtVc3lDjGJ6eRWZNVPB0vYuIFNldEbnNC9p0eP1
psL5gPuEME/dRRWz90OiVSHo3TKgDI1mEsytUxZNZezTfSJgAET4BgV0RLsmTkxhU4PeLEqTtdtU
xN98erCgJewAR2ErG8vlyPJUcGLjKd/P+wZScPfqhPD56HNR41A0E3xKd9CpRaPUFzDNvJJMrBTl
blw8w5zEMquvRjPN3RC6eHczxLyZhOOihmuIMfpEsSiX71etPPJ6rzG55fBehe3X5jqePW2UGgHp
VXSW8zB/llOBWfJ5iyZ6ZTySxWpxKnfJjYE2F72vsApRnup/qOaVzxOdt6HExYfNZ5XClypyMVXl
7zim6ftKibCyXohDWmUlMtWkng843muT/xN12JMTjv5O1uAlaU6QBQtBnP6ZIPQ4ABMnYpq0V4IE
yPDDNcfbaTbWbjT9KDTLXBp189fKWk+NWljSzxzfk6ry5CeO7pPPfS1QSecKEu8WnvKl7shHlZLx
LUqBdmkSJGV9rIOQrSNJ/HOYybkL+LZ0WurwJ0tOWQL2KmRW068UoeGrFTfZQkKxBz4IvWFQ4ExV
tjgmn1mNATMMrmsoyQIcAVh7GY9a6lc8g1ByNK2XcfxruwWYLs4oSCMTZH29KeYpXaFR9phuCUxv
uWuf3tYgABjUNmDvVNnIduBEiPoJSLlwML3QK/wOc8QvN9qyGVoIA6PWantQEyad2gZQjHztqkU3
6k+bo+rXTvgDeKKKwS0j33Q7PDn1liT1uhZu7r7HYpUZ1N2js0Ht8SebBsYFEG9RP6wW/uwBP7Nx
fW9p193myY6zaoPrPTfSrEH77YgiOVRFSoDCQZQ6nujPjRD9Yncc1nwzKzke1DPSV2OJZvStAmt7
TkI0nFuS+ga4E4NA0C85t9xlhKbG7IprR46iifv8mZSSfgzXUmYiLoP6OQkthSwVkVydv9hAeIh/
ehRaCaynuemlcw4lby9zA8Cu7ypiNvawYQeBTDzED1M+PzS68mVomnkNeHvKf1Lg6gKFn5IHh9/n
W/Np2/hD7JNljOCKYMjeZ5y1ApoTQvtwrqPSBd6WcJ9LUyoC0xzd02lAdoZwavMnI/yWQk2Tx885
2E0YIY0ZUdBCf/cUHeBDnyNgH4yWfFPW1osksoWttwTwt4zCTjy8+t5ebDf5KBTPCyPKnAFo9Oc/
Vt70sdMlHl25wnHgCwaZCfmf4US3UdnjA9w1pkpFqgMBg3bVTSfOhvlCjM48GGBSqweu/OoZbE2R
yqfMk1/XZV5f/QtHJLZ0CTQ4LcsOMT1vcb7mlueCPQtQ7i/c9g5NyV2oLwOj+1JSQwZnLK1smgsz
HwKrvFDMNyu10viPX8w532q4JtNJXI3AD+4vLvrpGu9NrmZqZX+VRD0pQMRUd37KWs1dMxfhkFiX
Hcm1cCfonXa3/ahlq1T61I3M5CgKS04//pIRXpdW5FwYgYt1iRBJ/K1pIhYccdukGGB4QoM9bxmx
lg5Ldvn5O4Hkq4TaIMZDdrcklij/8a3EIYMWJp8mNOJYAl1qgAy/vI/2+rJZyCoGut9LT47jFdlB
9VGGqu1iDvTnZRoOYdOOMrKB3LidP4LiK0vcwwBbOKlVmaO40oQ4Ss4wMAyODB7oEOHv66I5vIzg
SO2mDWaTdebfWtk4msSLpfgaiYsDUH1B3oVWEFDUtrKKKO7XdN2ulnynxsf2hyb9JIe4l8ZbUNtM
rUaJ/T7NLjFuRKe/ZuarSZVF+9gkQB927C1BJ5HPdrFZlHdzJXmSF1RBMB8bf0X8Sj1UKhnGLoff
BtVUFRX9UTVMFv+ooURkyN9jACEtt0eWI5lw4FXgvsZ5qg2uMC3h0z8+RZY7c6Gv1x0AzBZp0bzJ
1wnQ5TIh+E7MZouQdECmOiK5U055Ue8NlzwwCZMVHpb8ZQbAssm9iLYTX+rRcwre+f81r4skexeF
LFihxzSy1bS2+/akr2ggMoeA3/I1JwAeq5BW7Hrv1YnFsdHMiQ7el0cPjmXD2UNrSnlYXlU7GETA
XO+Q6E3nYkumaNEmtPeqQ3Ina2ykLGJ+hK/mUrb2pPwv/4EDg6VrNhUdw3yz86yT+vLyrxOJVWEw
IPySV2OH9vCzA0aMHbE1j9x7qKmiyCsNZmc3exEjVhUdxzKIoj5Gb0ZJwJUh/XoZ7l1cJ0O8wS2n
9wfrNyXFIxBhiO99MDmh8CDPYQqhVPo1gth7IP91cPWgfsjUBdVhgdsvIal3ViCCttly8ePb/SOm
7ZjVshemqF12X6/JYyNaiu1rA2sz+/YQ0CwGwtsyMfBfWPWQ72J4BTBEAjQRvRokuFHyW7GYR2sZ
yhTMKJI1Y56ruTAunCVEo2tndvrO9obCOYQotvm5xgY8djsRUlkCmn1KgmuTJmJes1gGfnhoB8sG
1T1O8KV7aJSUeivng+b/tHna09YF6POae+7KrJV3RDfPX+wTSmm7zkIx+kWXkezzDi4u/LxrznVq
vhEpTHc/Z4faAeQvbLUNKHDqknf1uSVswd7vFT5DKborCAmqvqdaUN57H3EWgbhqFIE+WhdM8fur
u3K1qIiOKKLJTV5bcT9nPFdeyNXDZcJUN1FwmjgXA4qK/XwR5WXNcLEsr8aYkAXXvejEbWXoMfTr
VxSVzbaRFwsuKnQnk5alDr3+2OXKbvLQCmapdrrfyXQ9IeTvsBSQWFQVnfVEzG7n4p8J/0WjPtkr
gYk+9l6saGkEhpf6Zhg6dLK5UjBoZtwCWq/G1hJTSNIU1+q7Soh5tLR8ffaUuyNRhM43hB7kxY7O
AxG6k0eB++sCzPiYvF6UjvDfpvCJJazSf355xnk/QRqc0CWf++NOvoZG7llaNQLT2sKDLpi5KYvR
CVxBJWIUwodu8SFEw8MNSgSZVopqejaQgyr6YATpVe3Bra3KPbrUqiSSF7ZuHs3Ru7DMeXZ/DgFV
28TMIwqvVXuoeQeuarZU8ynwV9fLYz0Ha1zl1QHV0ndLvqIKgGUnau3jvci9GW5mfw72neesAAnE
q7jjSVNK43o96or421nW4HQdfmmHVHcJi24l75cBnJUU7gWRFzja5De6JE3sTl6g31/N/j8v8Lot
3mxLHaDbzVo7Agzk5CVGJxh2d254Z01sITkFCDMx83R78v5L3IoZoeGdb2UrtIwm+WTK6dOsWIGz
puEu2L2mQWIRZpFcY3Go2gxRK6vgw6Pq9PkEJnBeXeRqGsGvQngEh04WE/G8bMAC56HsoPeHbARN
UsMdFVvDoQ+LzruNLbsEK280Hz58S1OFF8L3jzP6E2PSE/J0ZSMI7Eyms5UBDAb/qriGduq7LihF
m7EqcePVQL7twLnXkTitQ0FKwu7SoB56Ko+GDSV2qNmgMu51B2P89A+WgdJMIXq+vFBthk/AZOgb
nHSM0d/Y6lngMd8ctBrTVcrZiKz38VAKhbzuSZLeeM0zuh28Ws0tauqlVxQFCI4bg5cmM0no1pza
z0goEa6GzW00ghUMcTpbiISibEcp/b/rl42HpnqzwbUvQALgPPhq1bkgHu3bMF6BnzD4z08RaX8G
i6n24+wnnARmtP7Fa+QNnjl82WRSGljOCgJTFBjP/gMSGt9mTadbw5l1X+xAey5J27DrZ5aVyk1p
0npL2i54uz4fG67DPouzWB09nqwdBNk6ZUtuF3ZadjSUu7hO7FQUZloskwZlwQI3ALP8BNntouI3
a0TLsh+OIAHfiXq7WD7YxiU8+LiVwYA0yEddA9ztdl4D1PrhEwxR0Y3gD/0wNmKtpKO4bIhotgOq
sNZnKW3Hu6FFUPhA4sp9lgQ80ngJfBoY0b5iWErzp/CyoGsiV7+bRTgV0kHzB+lYI4ucS0PbUR+P
Y5v4Gz8bWUMtOU/zYJM0mFjbyx+2K9iSIQTtWk2phtR/Id8z5B6onePfKu9PwjTGt8BDD8ALx66E
Ic3yC4MTjlm4vtOxAGkHJdOaIUhrf2OBXH/tZnmrAY3gmr/TKQskjwUmNxGBbT+eV/FKh163D209
15MiO7ELw2wS5yyfv32xN21Bg0pmpcglqXYy2gGPfs8nJXAyoBdT994NWb/LEGFkhdeC8n7+hGZF
yqNw7yS/m0ym+1qV7e7vZH6gLC/59RLX/7OgrIgZGDfCYmdqg9DVccTb5VLOzlZGT6OJygWSzcEO
PZJEwmHBlh4bUOaTyhQC+rUbWpwnL8W2qo39YdJ9GNZn4OQFealllWsZMRpf0A2/Y1je3DeekW5y
BxuUAnLv5k9P4pOxVC2RhZrp9Mt4kkv7E9g1vTNuWLDlrdk7/Oi4gBT2oeod3Ht6NPKW34NDCzkb
DhLkhD6oyFhzuhDQJ9JrjTqI/XdAreC832j6UTXr8/Ivk6UBzij7hALKI9kahzwz6EHPCc3japck
ehMHcSeSENOYxDi1BZAJjY+a4eHIt+e1HgmOe0yHjERxfQKw5lCfmQB2GtBPOyxd0xCFINEs2sJ0
AndUwX4hHoqd1hC4AgMsTZo4qdEhpLo13A1tChP880G9w6BQYvi87dM+rM9C5C0hNyCP1xdXXVRc
+6etsd6221YKbFxSB6VCP4qxCTkEIy+p0+fRMsGSVD1XQG65Kinp2US3kQnCNmaxZ6aweu+i9uhC
rFT3pW/5MCMbvPj4ZPWsxt1MO7E+cYwfkcmkUzK10LqUlLvhs0wn3sYW06EDleBiqnJZZAobdczF
18YQaaZ8LtgDJaGb5dLK4i8gaM+wNSCpvLOiiXFDM7DbTwTY3/eMRpBvOolkdVy6zngPUrj+gjDE
9mLtXlVdvpcPgkw5fyek185IHJrSPU+CpGh+2wcXvMwjALEL4olkZg2n4bSjEml3dn/qkSE+CpUk
lGsCnlW1uJu/v3O3R4VjqIXBglhFH6HCmT34tgABREFN1M6Z9Mzjzhx2EbKk82C3rTCI4BMdQeTx
SgdGcPGpbhSoK4Z6r4OdmkAx9Ju+taMScS0XbfFSunKiD10xTKdOB1pvn8SYlsiyrkVw3UEJjpI+
Wlv4LDV9cUTNCOW5SU0pwFfZbMNc98quGL2DVXT+G+m5MLAor2hhNsQrnfHy99d71IWi8mTt+0SI
EQx/BGdnFGt8QILqnsEn8NK27DOIU2rFE0MM1gZ33bhNJ8w0IWYFkQEM/cxk6N1xmL0sKbxmmr77
/EzS8zWewGPaQBuJgdlF02rFXXXABXl/7+p/fRB5mJiUz5Klq2XhOeXNhEwUqDfkuozL9goGW6Xj
mLOm0RZidrYkJ2YFc1BLVi45sBN3vgpaI9rhsQDW06PG9+R5wIo62b3nuZHwTKClNOhRh0YV7bEV
b7gKNSRGaHa3eaWG3xIF87Fg5CmX/MneGdHv7UxWgib6XjOSlcIuBba3Ur2rEjt7oExBPXfti86C
h1pSDIKbbelLaPVrK1HOwMvUijBCx/D7vtl1TGjzb0BU7rGKkSQjOBZ/GCo4WIUjjX+6P1JHuzHW
ntMwWNp4DRo4JD0+PJXLhp1vZjLTtXSiJHi/sgjdaRDq/ogk+aDxw8iY/dkEDoyu31K1lOmzg7VI
1I0N7yRqChsUxBBJIGz8PyBc+brpUxVsbHnrC8fz5SbgQQQNVAGiXYX5APQppY64sRNssUgv1+HL
uLMuoup8WwoBLSEsUsvlVRJn4JeUSoczq3bHrMTvZmfZ6KQ8c7WxdtdYToQx1VVUrGlDGedRbnnZ
V8kTCgxFSGhERR9ueqdV1uAy9DpRBmYmM39uFJcFqW/flPPp0lplbY9GFVlk+l4GlNmr/48+UMiR
U8ZgNYb8SNc1hsXMfWvEX4rM5rsgyde1DTz1gfom2Yv/wVdugn8yNvSxFJQcYZNDbBkEgzGDG5Zr
QDXtM4EvlDNwy8FZ+FUvBno/H4xjC7+2Gxektk8f/d5FePvHYE5qT6V79HYkYpfViD7wJQizOr8+
/JZYf7rdDaH3UBJJ3MU3WxgbtcvPuUB+GRnowzU29w62/EB25jN8NWu6UFGVW4PTH6evcaivtXpi
7F+zztOInHVZ6qtIwEYvt6wbX0PH1KqN6jNB8Sg3hsWcm5RTBF/kQxqv1QVblgwZHgg0ElLj/Jzd
3fQpbsH7tSTIsLwIs1MCrLEMRTdqZ+azIeUb8LwgsGqJIwWDPKXuc26ES54m3dMIR6f2/0XQwJjL
dwPFvNLPYw962wPiK1hX4j4Nud4GhU1IsJe9DIpQGwQ8RBw7GD5eG/YS9iGT5gr3e2ysOXW2UUeI
MLV+rbF8hlEpCNUnQ5lglXBybcX2+VM+O5u5x37coesIxSb4Nm8nupC00u9g+aMY3u72AgfWCu+I
J3iJr4tzRfvfRlin7f/wlc/ZfuzofFVrRI9q14Gqnaa0ppukO7O76P4WlEKKZMW2fEGGLeTdIx+G
zwYz/QPyUWRq0jWdfYm2iOS+WLZ/sVZWPHRInJPB8XfJT8KELku9ORFaHPy2P+Ak4VP4BOFIaBbA
lyGUO6F1AKTf1odRu2E9vBURU9onm8Ayg5A032+aQ2QyuD3VKTvHgPD7E4ABJCj8wity2PPzROkp
etlDVZq8GDatflqI0oZINnYPpf6Kq2TZngyUU5BSIwtUfdTtP2KTDTq+3n1duBIfoGohMXb33Il8
Tg9VRKoc8QHGHJDLz70sEqUwfBni5EScovGZz5M/CFnCalO1HYzYbHT8A5RrgNRDE+57+QGAOZ0u
puFGdh/2Hvi5D6oWFxww6dTg60usPqOuJGzwW07x4H4QL3poqtXhFIdl/qJApUMfhKKQAVqj63dC
0ryGn5HbgHbe3b2EYHH2ZiI29rhYZyi1SfaaphdwRsrtoe1mlogWK/yMVkf/4lY3hEoF6ymKd0rY
cAl4swx1W354qg3Qw5ZKqUxPn6taWIc+mCFXKhhvRlX12rP85t5q2fijxseeTnZVK3D3pbbhkKQZ
4ABOSNWO3GpME6oqX94FtlCS9gaF4l/lXYkPRknbnw+nccfkKq4ANhERmD/s3YwlWNK3z69/26Sr
q5nCuubIcx8vgHut7v6o9F6HkzgLFkcWT0MJcQPlOPuLVCDC5BPPQiKPjPh3U7ggL8eb08qtEAGv
i5as2/vy1HDqbnhg3qbvkkuagGRaNYUF2bF6BiKmPH7dlp/K5q6/q2ecMa30DiocfIN+/7V8L+Rd
EQ4TV89YDNvdQic57Di5dWN6ZtzqAKoF6NKPsiJaWyjY9Ga47YD8oB93DE9aBHOsspHz6oRp45qz
fkLSn5CCpdlNB2Pq0bdXszUI4N1iaFfjzEZ61S5XshrNo4SwcYTH6ml38M4DNVtEAm5YyWspvlUN
aaMipZelG++WMcLtaF9ILgOXfjQZ4+bVhfXKx/b2aAp56sZgMO0TGYDOtKm5sD8CzAaHmGwuyQlU
a26XJJ2034zVf+vCgzfXPGSgy++gS9jmFkh59n+0N95sKyPMD3koRofU6gRMVO3hP3VLz3pKa7Ba
V0AcKXWdfBygrzIXFBxM2mMVBHPK2c6lP+dJmhgnKjPKnNiQKTWAf+E0g7Vi0LYutayNPtnhTcNG
RtAvytXBzO3oYvHlPhhqjaNEHSNmYVd9JQ29nIDmvQftbLB0QhbYkze2+huO/suvD5yFfaI8SY0E
yUN/5ZWn8ZL7Q7nuqYEcUWc23R3EUdo2i6rchFqCbDyzn/mzYClJZJx1VLii5Cq1W3kx6aBiEIEX
Q78N+0azYvhOwH2xswGpSMCHL1rewODeezCGn42j/NOdGJJPA38kmCTjNOXMvMmCHDrjE/kD6fXe
+WRbp9DFmLTZfq3TsJGTlADfRodC5gGHd4KC8q+bNTACZeNT2mUSoihh0rFNrtewCqKO2N1g1WWi
DpzahDLT8vZDBmjWOLlStDowfAKOSFRdK0ZuuchuYSVR8wccV7SltHePjORWaYUckhaEQ7j9JiJE
/BuhfG4/LheVrstfGNtcs2fc8hMsnp1icCKH+kpKRar+jlvM9i86RWsGBCVUDPOmR67Tm6LVedN2
bj3YA0VFGqNzHPg4enATeieEVxxYt0cDwlV2Yo93r3zWZ/8Fi+tNeasPJSlq/z+ky6DYLx1gJMW+
fitXkSdAHynsJlokZqwZ0Ac4HTiNRizfEdss+vvx2IqpbA0h1wjgz/LZ2Uddr8EMw9qmIP/+B1A+
yXI8e8bi7woySm2+dE0fl9O173cmCw4TDMnKAlYPG+P7/EIO69fdyI3I3C6bVlcgJehA2cFYLYkd
SIhsu5NkGEqOYp3KCBrpEHt0icAqOnC5+KFpPYUY57eq928gInogAh5+RixRlMaF+szOyVaiCwbI
Z8VRELhbceCqeO19a0ObQF04Rw85M/ZyNDBH1t1nCdIQSWN5KXysPc3x0ehIIij4A2ijMw1X9KGg
CTs2bmnPSZSncqqJczMNzFfc5l3ReoTOnbNilV2LQIWq3dncSEHMGaGCjzUvh9YYNDs5IfldhRE/
gnkLXFrJBP9BGdhxLeS3WNXyQt7+9UUawmS2tXiJl6CbUAvy3NI1DrB3Dv4rYMaTbfXnY4McSIa2
bdsPqBCDeuqHC90FG0G31pAERx0OLwCmBgJMJK0hSZls0+AzYQlqbhYr9a1Tc6qDGP9eYnlK2l2T
GtMwdEdAGSHIzbT8qJu0DB575dmD591i1bVcT5Q97N8wHhvq2yGdD0TwsX/T03kk9qud15seoim8
NPjfC/62WSq/0PT0Js1q7axjfgU/XSBzMR9DW2L+l2SOkV8ctl6qS1tsGa42VK1DuYTGrmsCHDUN
hR2D8hsKbrSs856OeIftVFzEnC27aVzX14AqUNdCVCeGYFSayL/edum/Q+vlwyGBMhxTZCBdw7w4
kZn2QKd/V4n28rWnkGH6cufKP3X4RIEC1670REWXBPDUEbgf/T1g9+3okJIGAYcT4nwWNBBWUcNU
Wz09hV0lhi3TOKk4MTDwtFaveB+O6rwHYpipUvau5VS4sSJZgPnmnTaHeySGQcLy5FcFjHv+xq3w
rgtpMmzxEtsquGkEi3MBrCEui7OiAb8GuAw0s1aBBd2NGQnRbiJzjDg59QNiXTg4b88bWQhQq12M
ifMA2RaGfRpSgGS6SVLBlBeWJSXE6mEH4xd2i/oPmp7Or7rEkN5Aw46f+Ged7VMOmMwxGy9wIdJU
nctW8/uTTS1faqChBAeSn+Cuihr9NF/Gl3EwVJjZ9mUVUKI6fO5umf8E1sKSLBqPCF3/HdDCRCKD
rYI2IPlnEYu0b3ZdAAK1wDAqxwecs01sLRKw8FTVfRpiID3K8JNMl7FIOVWhpi7Fz6ZmeRVxtimF
mzr5sh6sYJjr6aVXaeh7eXU4WX/UnNo+QVfdWfqDIepbAQKKGV+aZlOVcmXi6l+XroFiylHOEPbm
OuwrOoseBlHkNYnfWSQBJvNQnPsHliEgeNpocv0oqaiD7GJlEVovQNVjvtgYosjO9Wifv9zgAnLL
kKCyfBxt5lUWAvbitY7/8IrMiVajpnKeRrvMj+rIPOLkafkb1DiN1/l3szswLaSzNp/ys9HH6jCQ
Cc0J2nOq05wcFmOioTwGh6A/JB2orskFdXKu8nnQUF3V6HbHB55pkH9OHfZT8SGqzGL6PIe7Xo+0
wD4yg0FjDHwvu0KjtC59bowxuo/Q22x1MtEQSt7z/mHaXug5S4thcz+IP4KybfZfa+9VMygCDdeZ
m5rvaLM3d+IfvfvC4IiO3dlCxlNBlvBENydQpgR5CMKuuWR6THvSyEEbIUb9a3AAhhQigxzN/tBv
wtMbihWJix7PPfZx/vK6aplHnxgp0a5PURf2j5BqiD2OSr4S6Q4etdypJ7a4UeUWAyIKiX7itedv
9JcTyQuwmyvzT4pi41aYvWNE+nGCD/RlWagM1GStw/3sIUhqPcCQ06LAqNBzZDMBBXXyjMNFTdIp
RMZOL+bdFFLHx62c/F2srOgiFWa6l9RX130VvRqO7BCIX9UiJAqYLuz8A0yOGbnA9P06wJYjRh9l
OTQvw1S7b34byRfeXV57748vHCNQi5KnvFzsfHK+ljLsnJGpDzRZZlqz3B055t2QoABp+3t1EwQx
yvMzjvBbV/U9LFu5tLeiP+w44+LIYMn9CTdKBbMSfY8N9ViEdS4yuW6OVFd6YAWwEBGGlGMKB0FR
AgyHhtEWLLehvT3cA3tw7quyi/AA8cVJlILRCh2ftDDsDGyuXEjT7CW9GSox2z8VidT+at7ZSLY/
dJUMdc/jgg7Fs1iPUXedDn6soqVvwAxiS2J0Y/0Z8dkbu9L7R/qOZsPJBms/umQ38pyyo0Mxiakn
TPT828CZTRsXEOzi13X+j8UM7NfZVBMXNRYfZqRhCrA6RtxQ9ZLKXfI1se06FolXhghDA9bJxZtR
ocfHT1NMK7j7gecDSGKn97o2fo13e4rOtLWydrx6I+fPkrdtnZjKzCXbllLWgTZ7k92DOlw4+dqo
h+ti851Pp2XPglIpNeIpJnik7IZsx3ZU2tFnR2q2YqwrMg7EjwePBndjdJEMUU8yKa12nNPX6JA5
TZVJpsseUOknCyR1h9FWTiOg/5MhFX9zJS1xg1yhSVV8p801UiyNmAozThmoKHU7Cnd9SkAwxoP0
0098SPRIXG/g7NibAczKDH8a7fc+Ecyt/MObpyvHSXZQpm6gmSIWK0L/dEy4ix34hPI5qkuseKpl
sNB0/+uMzMtC+VCsNCgWxMoshTYujNilnn87cA7W+cn3K6hjC5roFau9PszPN+gNTq+ypseTnthc
ZZmpkrvu0QmBizsbF0UV1Be6tWiLW8Z2XQbpkSrsbxQ2Pp6SQ4cJg009rPyS+QQIxts6Y/TVx4WL
/zZZ4KslKaXAIEYjSneLgntrp818HYLoRfUBgRm2BzvQIxQ53WzdOUc6E9Xwe70DqI9OY1+ovizK
UtjU2kZtenCES0+XIOIu7BlbA5jZEwWwALaHT8Fo8RHU25AqTFkyzY54OWftHEV2NTaTBIDAmNBP
//bU3lBXHTH4brhR40OVIx0vzNKrOIuOrMw3sD4YRl/BHLCqI1xEkmFD32c0wBA3iLFgSqJ9SLLw
WwymZ/WPb+yqEiuSpGTS4MHD+ae+AzWvMOuOK4h5PCGBVJV8tsFKhwYWc+AwXcGzzmY1daEWTZOb
UvCl921krqu054j63YUSWAMcfHZnSyLD+xw9MF8dtSnbOUmgnsFxvz2q+LIQplFOVPo8/Ss3p5F7
qgFZYI5M7QtxxjN/LwcZlCsqAoHf7P31axQSLWXYDRRxemygT3IM6Vr787CD1STQjYrf6+bvoBkn
q+KhPrL213QCMQgUXPGy37JG+f64+5f5jkMlMmm6WoR9LkIdhhHmhdkd5gctaTLG76NTuNT41LAe
7myo6YzYW4eAYi5wUO+trRY5Alm1E9fb5obm9ZovYyRzZLWFB/w+k+Hp4C3+zYblOUxmKaKgJ82C
w0/YdAExh1bswupv6HqjiWvgAFHZZ+r6ZATsxbBtmdNmjqNjL+CXL47QAUOzqQEv9vhchu3R1OxY
EbdtHTkoMu5U1wlp2pY6+dWXAogjjfwCylRtWR7CKI7RlWH1LTbkT9JI/jtd/ZAHh+qvgrO9e3KA
Vb+AP85aHmijRhHnZXXr+39jOmJzMgXtnaZ0yANDinIxm1nz4FnHOMTQgKohuluh4UHGG/GNdtnd
qglvfSChqv04nMXvi0wCbbSJeMw9enew4EkfGoJy0lYFneNZB4RU6TFR/ZXkF0viySrtmciDgB2m
ctm3ybI0BoUTpMWZf/t8UOXLUQt4TF7bq5qJBiH8NcOeBdukGzMhPGNcYDO/fhQDElwCOJLNsWJv
gZzIYoHSJfk0HSU89Z5J8C5+qyqsy7SOnmZohlPBvwUSwtHGtggMYDWjqW/eVNdDqxw+2C6qPijV
Lt4cP/7ddytXLVvnbSM6sA0ifAYwALcz99/qAYpQbIGRYriNE3iY0eEw8dqBeb3HX/ihhI4A/sjP
7zA55kc/x6blsMzBXhSI2l2rF/ot0/cygrW9qkBCGjYW8qooPqW+uL3HeYIshXJBGC8EoyeZUz9y
VeQg8asao/WDq1FwnoiI4q1E1cHiNoxq4tyk4HOHSgAUT3iXTrD+C7d7mtiH//B8BrfdXgQ7OilM
z2ca3ACnlPUrZn4EzDaEqlru6B/sJ8i3ztPGL/NzyhkZVMVuYvfcVBSaKDHNF2OIXNEzBJuMgLkW
SlO4rVXxzFx9jAguVaNH3j5L6l5LAx430XI5rLu7Pp+honNnKtFIDKBpvE5JskvBhtKW2tULrFRr
U51oZVT3AY89fq4TPWvlK4gL4CsoUDLqZPqGfGq52Ig33Rs63tSckiTFMZ7y79OVwVfTLdiJ7cWb
Jua/pEizyvoKQFZh5j9f8uwqV+uyozTycyNov0h9tza97+RLIk1JXdLmzIRaZyz9Rh32xsSo27UB
mWUh8Oah0rbLHckxd9VxgEiFsWdvqbVQ/Ztcez+/VzyoSKf6ZYFdEO2LdwhDHVvCzrqQj+7w5042
3UbXGsxmE6aO+sI68yK3itRmS+LjQqfoCbazks4DOmudbd3NCXLCFnp6SnKH+CY+qT0W6DCkRo12
3GlW7oUEQw0AOiml6balaBQkus78jVMaydfiUwPJPf9jVW4niAQCMwn6QiscKDRtHDX+GlSczgPv
mwBwHpB47rxaOIJmKQIGObJxe8tpbfPWlAsmrJuoLvxdAGwBHovONxSV0nNpbvt53H5Dc7vlEtSo
Hk9ieGRjOIhmIrdjHh0mwdYU9e/uTvS954qQ8Qn1RWcBY6c5nUCmJ3ivt6CioEwCxmo+2oKKu0fD
NOuxfTLwXG8Y0CVXJ2keJXSIBnVOMzM260CjNLo2rDwejRY//K1A3dr1m1psgSmQHM0IvIywX5GO
njptRFDUCMKs2x8zkWl1wCroHU7sSgVScyI+BF4/GZwgqjyHT/fK/dsfGw6pptKMiotQ4jlOBW4k
qCt7d/CHgB1IsuxkMv2tQqYz6uXOEgOIe6ngqlrbh5CPRh9xuiofa98676kOmGTzMdWT3ZXiXe/q
asSvaapKDFVRpS9qJF1+Q4/XrLzjhEi1jS5wE/isfcb2CCxxUlF2KwdcNcksH9TPhOgjLabhuOcn
NhbxKMhx0P5aIIUCJMnq4K/7zqLDTUMED7G5iXzIMN2KvHyUSGgpPA5uVOf3FUrOKysnJBsQFzSF
8lSQluAN6neeLDEWGcFsR/aI/qVCdSw3ByigjYyhh+hkWDOXaHrNFeT564ZutpAo2YlTM0dnTGBS
q2zM06TfXI1N0V47uqk177lY2DQa1Eo8lJWV0md0o9YwM2yMt2yXcIemhr9eaDg3YL67DKAHk3Ed
QSK8WyDjWeB/k//NGYq8uJ5BPHROTyXoOPBIFpWowiXyXnB+VUMWDS00Kt3PISP3csGsU/sLAWaE
iMJ1J/qDb7xOLtXen821MwoMlVmsbvg5M/0plRHXz0JEKcmaNO99vTCZFHNBJtST+FPBTmiri6UN
59tZJYbJUE0WK+CVDya5TUJj6O4wgG3h7a1aZCT8Z+BVwyXJ3EOSlYEfjngX+rLiHTTQCvYxEPuo
vY4tNKndPZffPo24NA24/clRDjjefvmvFF++G023+5Oqj1sGLhaDMw1IN8WDVoDXtN9CpwVbx5ar
3/xJ6+w9WxKGm7bkhzxCTAKjgh1enp3AJEf3zWY2v3QC4XsqWDjHRg50g9i9k38hyQZzTxlXxQor
xOs9AA7jNqIwOYjHD8DvtbBitrB86XZTcxzhljzvfgrD3Ogx6QPd+tBHH6kmC9dGwDQEMc7/Exka
EHD/uTmKdYkJNGlWY9GQ8Eq7MhZrQaZjAI5wsbJEIXwLXOmHDrw3u1RutVzU+e7Tvpmdwtk46gVH
+g3xQozEnk+vCpgutyTJW7qZUPbP6PxnGO+ACJRot2Sb/KXQNFe8Afp7iWAOrQ5aqPsqVvMRkq2X
B68qbQ+K5SQh49NA3z7QjOH0rYyvrQAZTRU2sxClOpYysSnp71QmIjC/HcuOkv+nURsu0ZS7mtt/
HQg2vpEbItGlQ7BIPIQMHNwWdUP/Z6d5uzoMJ9RlGKIBcQUS+k1vCpRXslYq95r+3fJYxu4AP++M
sfnANPNt3z9OFxsr8Bphn/34oUj2lJ07kEXWm6RZ2Tt7uiJea3XLVVBIMp5Itg4NQPxI1AdvSbmN
DE8NpcI2TkIDqjyLlktKyYXA2NwRQZLj9nMYlLU55lTdGoSPMIEQ99XVbJkSPrSJ1BoO99w5/vzh
GTz3iLh+NVW2dDCuXJmaPrOCm5P7V8sYYdz15fWDX0RT7uXL29SabbB2OxtYtSDIcUK5GpTRXhr8
cDJiv9Leyg874lm2vZKFQN76phmSZh6a6LQ8e9xysRIw2z/W41Q5OKY7PdcjG1hYxOZOIaFKPg2K
0mfBORpl85smDe40BbYoK8S90PuogxcP/qJ/RlqS9Peph4VFxp+irc921G+x8+mEvd1+00njDqiw
j1W88cfskp9NPZJcxKSpYyQGzNcS6nkuAsTmRZUxoALI51xUEpLmdk5wNZ0JWaygHfKublicS0xf
cRvWZyIUqjAP9A/o8mg4NehiJVDflnE9/Mr6lqSElXBHc760W4K0m6yLuAhEsP54oPLjO0uNgUbG
S9zzkrorZQs86lwzbgMJpgbkhAJ4IK3ZNaUrTHEqP0kypPhaES79Dl0VhRTX02DREDEzWQivrGuj
gpktZGK281xcAzqW3z8ZkDeEXmwR0nc7HYPNqYw56dHnzTqXeml9Gi/L6+fp/i1+so38KnYM8oyX
nQtI0u17249HfhmvbDoXCZvurZF9qz27QUjhhbuRA8ac+GsOpjw8CdlErvKP1GaK1WwHvvO6nm3E
WKQgnb4Moae0P4nIh4nW/Dpg8T43XnomjVk4q8X/Tqy4/jKRXE1payn8pmEqvV9RDSuoKiKDaoAD
8Mk7REKkQn7tsLQOgx0AYXhFH1+bqIIf1wwWHsbLbXRQV1kaFdfcG/jdX4kxwuczeYH/gsAGNFf6
SXZBETedFEerwQUdK2yEH4Qksdpu7zGGpDhp8su8fYP0yiuyVdoL21SPxLWeDevWPwH2qOWMwpdy
I5Ml7YwXGWgnCcgEaypubkQ+9B3z9jovFfT03C5vE8C66xjIJsxwWsBp7TgfEo5v/URX9nBVFtl0
SrdaYcKR/i/qa8ZRD5ei3Y3XjpHXXedXftrr+REuh8CPI5N0NwYNbQYctBHWAFJNZczs+KqKn54t
DmsXfK9ViWorBSaqsjkqlTudwzGHS8m7xZerKnFHD7QS5oYoeA6V0cIt9hNOWcLG/a6Cmtab53En
AA6RBSg0hswwK2TwBXW4+u27T+YggvB4OLrIHdcv1+2hX9tynA7dUKj/tPGY1Pa07wgRmgqTpP+O
+GjGzwtIzo9duU62LUOBZ3n43RQoD89hQstvPBMnV3pW8Qsr630LMHDHjJXEkqU2sdHAb0QM3Pb7
sNJfarWwTtcUBvDAbxZztIj234NLHDFymGueJOZNv8DlM5+wVIscEOi3rzcXo0RVJzAwkVwOVYO5
f18wM720HwCxgn3J5I2znHwh6+tC55mPdmjdHGz82iXGIn3aDZQI2xEG/dYM09TkfPzQFl3d5eja
TuohLpFAHxre/uhWi/m+lI0cu8DBAV1P7BFta7j7SiR6A/8sPLCCiRtTmEO8syKF+xmt7++OOByp
1g691b810i2YUNI0Anaz8MMY0AKx6DxdKa+262WTHKm5cR5vgs2g67s/HRV5gtlRaR9yllB8+64i
GjVDeqIj5WBc+Y7fxfW3Q6rF7Ycy5j+BZ8p+S6sP3OkgOcqZQDv2V9Zd8bMVB1u+W1h3nlEVFrvn
WqhOhU0g9QcZR+ruTYe1ybMTzEmyhZLFsrpfBgwP/O9jRf6pQ7FBuI2I9/27cwWVHhxn7v/B0lWm
tasnljC2MGd2/q+vVzgxh/HFM7HrUh2d6bKAcBu0+03LfxZ4FfVHkdfmIqdRzY4cl+hkndGmGwy/
HNqwMl/ZdjumAcCjGhK82LpVjlSoPKwMHjnWfobGjMPU5chqzlaqRtfdMoS/p878FJCnuOH1BzsV
4OAoV5WatISbMMb6fh04jfe11w4q3CoeRjbF8B33HFTz/tLibYlK2+XqJ/rsFrDk1eXb4oUum0jQ
RvoLs+ICM7pwblc6+oXIwz9NFX1SzQGX6QMxfF5YVwSmkOcd3o1wqrJB+2IkoMagFmUsx9plEXU+
40gu8ZfLNhhBVa71dE+a2nlp6SVuticJR5kX7Oc2ob4Wgf1BUxHFdYhmhiq5C9bYq13ncYO6KJOo
0dsBn5UgCN9i+6UJwu6JP5Uo52wmy1i6/7kU946bamu8w78M3I5sf6/PiPdrpjvKBWpDwM8B4Gbj
c4srzL7IAdGNsb13XD0JGR9WqQJLKeLuKAV9ZYSHQ8g0waa4qJzKn2pzh7QJ2tm39jfKI5xq12af
FyHeTM+DNa1n53FB2qeXhJ4hRUqw8hQh9QuCz+A/Nz69TrZv+Sl1M57sQrSYQ8b483M0MOfyjvzI
Luv8dIMTWLnEA1AARLaZWlRqBJX5/9Q6e39p3BWjtNUWyq/eSUX6z5anrnVkOXp7SitkLaIHXwGh
xU8ID+eiVRdWMwR4qjDNdq7PEuOC+Dr9kvPKyO8HDxfwdMZLefjFryxmYHfK6arzjnSbrcxkC417
dqjxWr8DocBRP+kRBiTW08uAPX8vJAET7v03MuY3HCHodT2RASAgaJGrNsUXn+k9GyoE/Kom9nv3
SKOipgBDEJOGpB909sEoEuFoV5OrW9ThoDm3Alf0zUKNiIyfA/4zdjUWWs28seNZPlHyFOPKgN6I
WbQo5qFZ9UywPn6T89BS/o+4fa19Bxkb1U7Ku7+x8v30uksxyk4pCYVld00Jd2XTTRUXOB9gNm7V
xEdI3n7r4yLooyhStivdWpeiPfdbRNrpFKJzwTwywRCUSwuGBPi200yhQJ9VF72xWcrUcoVjMfWe
Rf+1i2/YwggIT/Konlb/PAh9IYPTdSwiceF/j2absaS40D/rbsRHFlMYyZuLS8UhF+muhcOwPZOe
dRXcuF5scbs+NpnIeevHD6uimDg+2jwocAdFe2zZ/p/eK8pMIt+1f2yiSTVtQYXrq6rc5JQvb4uZ
/gc6hgUDaQ7r4RyjU6UzJD/etTx9ieW3Y2YRAq0t1zh4pr8KIwuEO0qt5rZhx/JbcU0T2ZyqfyLP
khogB2bUJHaS2ffKeOl6deQnTI6nYIn7+Q6EwbAKwJXF+hm4z2CJJBd9TtBqRQYVuJpBDS14XDL/
7YkT7qlrK4vn8GFxZmF7bfl3w0JGOYuBhHX61j3hBVGYdvT7FVCqhRK4g+il4mInojm1qOqOhsoJ
e35Kbd3B9bWd3F83fZyso3rYP3aECFykY6DSl1mSBBvQbsNsQkgbrz05l6o4vHPjMFbgLAo1xXMQ
F3edfwq+ajZIhwseSEv9zFrjoOzTO+gJ8mLcnwUuNf2ml4Ts5pM7HAAfBb6YvaKByN0x/GGvtQMy
nJ1rDurZsRgMNm8060ZIExpWPHunNmA6xICfr0Q1J3YOr84Wu3fwd6zm5JWSbMbYz3phS5yH9iy9
f7akpEb5UYxg1Hcstq4sz+Blz66nJhHm1Jxx3wfCBjcETmySuXO5wQQPWwZ3TV3RgWKcSUGLQIB4
IwBsoYtMqfN8uzV4rdPhbGuN+uSsSKsOL3A+fmBjhLzMW5syqQVCZjvlF/OuZTLgyWzARvaAje5+
ltai7t/oF7ISY6feODv1veoHvBm33RjH3/z53xIB/E1jo3aIk0Q/5RAS9TbNFYg4T1sW3i6P1C3j
666LhwXhNbHTL9HNT0JGnYGFMGuYdv/1EwjAvg/mmVV5VpfWeVJkM/egSWZvMjsGZeiUUWl80z2x
fLHo0sNaT8Na0sHSLt4nQDhmNMAFRQlxOiohPRU2PqtNj4coDKyY540K9XGSRhR1syk5+XNhzoPc
NXUJgrxZkT1e2Lv6hnhUL4tiUKl1pA42YqZsANGiUUI2+oENRElOXkTQmKx168YkMCq+AhdJOmIZ
5RcnV/wnlTkjxhDVCvIrEvBQ1+hIagpXJ3TMUpYDO92b5xEtJXoQaSAOIfY72pLUXwglVwwHJUR5
FYmBEnDF58vU9McA4DAHtu6vI+Ki+WoEQ80kQMPCu89ZzjAZZpQZTWsvnib6wmS1WeK2sVAcAXk3
4jE9qNdy7LYbi1/T0ZB6RvDeSUqCgZXTX9UTNcChxJMtxNhDy6X4uYlkRSFY/W3AsI+6QkFRA8em
y2K67LEHE2kiFNd4dO6hqiV8OCFiI/uMoTkP4GMK9LCTL4jt1gVfJ3cCWFLXDyRTul4X3xk4CBSu
1Egq9MpjuwQCJFFPu5X7HcjYOMe06AMR8Q1NCgf3LktND7snIk3lklwxyzZcyaeUOrCASQNg0tMY
KkoEqhvuSoMYyK69xiD9pA9V322u3Lio/IsGlBLPdQuUJLZzp+ju6poZzkNG7U/xu6wNkbct+eC2
LP2sQCrwkIYFiGsJPHnpIt707CiAf3zn0eeuCcaGhC3UyMlKzJr+D6cpFARh9bRPhIJ2uTnbYbIz
vJDs35G5hcZsR1FBNONxSUjocF3SsxPQNE2M2C4jYwGmL4Ex+0EXfrxOdxg+7tmxwe+fmW12/fFN
JFHcWETljNS3aUrjcxmrswZ6Q30jV+YeQAni0tZeWGVvxnb4r0qFxyyfovYiL/6FXEz2WlBkwYIy
CC+cCj23rPHcLht2ZvSiUbdEg6MQafuvuVtpfmuWmSdm9ZJX9bljbHR2P1lATNsr0djaJextoHSA
G6pAxXMAajqWSNnaRBDBd7AlzeHmYaApNEd+rZjTRJ2uyRd+ePbJaViHUgZ3oR4K0Aj6fptzBDHr
FDtcfraeySrqbr1h/o5jf+t+lDTPjAPUf3wbLZcRQZb+jhZAEHhzhnkVrNbsd0wzGCCbB7hvMPuk
3HvxyFtbn83aFdpHDi1YJ2SSkR6lhxl7bmMZ+e4MyF0D54sMQdcHqOC/PN6YUxRyi+vkzsChclxe
8LyOHjDENaTbVGlZqN58ftJo9Cp3fLkpgK2/94XE25qW3cNPE/wJa2KKvpsNYQN1+sala+AJI/EU
wtKuZWiXK2e6pVYeWlCafuBvoQHbnfKgrDLL7vNbvn4JeAkuPWLNNSeDddp207DCZ+IfeH2xIOoU
LYz9bE9V1Zo7Nq6L6w1oPR4VPmHPiVf6GmNvMwQSn1qVw4ofrXPP8N9h36cevyCqIoRnixOZNpmK
g72fhYIbPvIeCh7q7ZlHviyiRwGFsTIZolU2d0VQVGwMLAIdtqCI4yWn9OVJVMZzBzrOhpCTlxjx
E3IcxS9GnbP78VWDEygxpAvOSLp4e43LyvFQa4PPbOinEGoku3PypcbWJMWizsx7WE2Ieue7k8wy
2FpMh/wI/8mL1U++v69kUb3xiXrazYoqOImkgaMC+wd8bsuC391WYPuNuraWeUuKEV/wRsvdWHRx
AFhuAO06BRtArt7+foPuYlH8lfBiTN0hUNDppdkpjL0OaBGhi1nHEiaAT+ts2oWldzpx7OO+6Rp0
9/Aa1Q3KZOdB+Za6REVzNvU69EyYQX4d+FaIRNXua6On4SvTWP9txPK+7EJtDcbiB8Sq7mTLtT9S
Ciy3IJki0efFjkNLx/SS30Sv6a+Jh4WwWcSmiIKSr+2ktr4sLIUDD7nm8ZqZRtSrtWQPzOHuKp84
stWbCTBWAEwl3nyoP6PdX9wdnYBLKe7Yg50FzRwtlwm4BH8W0miihCCeLiZqUQpbHv7WzsQKBkEZ
r/iuoPhw8lCn59YwrkI9CF2jlQO/KNRqNyDT4QBDN6u4RZtpI9DwwAG4yj8x0LR1fBlRxWTheIR2
eId0TOovUJfVV9MlC2Jl8FTj5jR6qlBnKO102eq1V1LDAvxvbSdXHtPiTzWn0vwP50JFSHJi44P8
77z4Z3htIVv4Hvp+Q/GNchaTIKh2rWLFaK4sE3LFTlS97WtXn0b51Y6y466usRA9pUys6dfeMLdQ
OiQ6heEPf8HQ2jFBbm6CCNVKaWu3uMKopvyqjCHXxyjonPXpF7Gslw5SEJMIEiBEs35w+RdNywaK
NUaRIv07CzYsk4iDB5sMgbM566royT6stWy/8dx5dTfBnN/F8jzHLHBYrJJZuG2W4M3TKvlwW97C
vibc+6uGvDPT0B/3BWvpA8HleyfeoLXAbh0s1gIEsHGSojK09auNcRBvHdx010TtDculPeIb6uPo
MNDvYmqkLDk3dMMeIqAPfBPh35cBRaKcGX5Z9ZKQ7G0MfCm5NKeXD0Irz3xpcA5MSUxfRJ0VZlKo
BkU/WjmusPO9rUCyTliMlAdAvocm9Wfh8ddEnegYwpyEIfpx/272d5Bf6mxIlCSAtlFBHiidF9Uj
hG85jwNzS0vDKhCKLmhFnO8ZItxrf0smH17r1onXyiLMzGOPUPddj8JNg5LR81MMATgR3NDP1O/L
lCCPgpKFp2kSojVvAt4lt2pvAWSgcotCx2trUZD1Z7k4Tl58q8xvjqVfHU1ndNtz0iMSsvpjxaxl
baBeSub9Xwlwaxt5ut4cQZSUoa1CwpkHE/dbgHAlAQ44hiIqD9CE/sVUCILL49bHmsnz1AEsKGXK
GFDLgRa8XkCEhJRpuwrmxCpBx6L7n2G93KXMznuI94rYFAD6SV/jmD41XSzoGtAo0zCnpjRvGrMs
hg1Z/PdL4UjppIXxMWQxb1FD2fN03UMPpDKDPk6xzME6NPkf8M60bMJ+QiW07w80b1EBOIcEyynr
PdiKURYMHywcVHT+1dhAAoLBiT5FK8IOQN0uF7yQjvaBs28sJfxBgs4SNASR44VzFYldSg1Q0+eB
TTTfRL6rB/fUJxZKj5askC2HyOBAwPDmAGi3OLXTVlbaJ/uK6vV+72hQ+kBt9ihHdJZPrIc9c/x/
AtbKoDHKc3pa/Gysqc1igCrSXnmRehM+kTDYC3FPPi5kawlHikbCHJqSPTLeIARuCInwbgbX0Utj
wfi5bCLe0k6Nr2xnjui5NkbeNNr89dPHuOCLYmp7AaryDUp6qzhzvCJaHWku04WAfLz61spQeiLA
0j9TjUCbrGpMszzJKUOg1Hcz2HP7cPMLxrgkEysbOcQeHOn3PLJ7+PAAzenDloi9RhPeR+MA0w8f
wk56l5mgHXZ0H5L/i3vOgNZWp3Y3mp7T0sleZSHT3NIkym6df7sWnymhrjrnsB7uxO2CAVw3efHL
ePH3PBk8+qolXRn2uOCSHNj9iOg7PYvbdJW8FSDtiPwe9hPtA1+2SHbW8ZBLI9CNKwAmt6F0UcDl
xk9986kGb912qskeKoGuWMqTuIaqDW8I4y+vcfAUfOh9MjIwPX1uBXMnNnmRVpcJJ9YoumgRlQ98
xYSg3V2mJZIxWueZS8FVgysxelMDdxoddF8f/96Bk5AeAUE+w19WwkYdS43C0q3asnozqLMBMjuq
MsfoSGE4P+S5IMtYF4AlD54LwavvDSLgHH192mmYoftWWCNJNi6Zh5T6is6XseAEIi6RW8kbHxw5
n9vT6jjF6GyFlFllfiOFBnw7PX55oyv/i92qktg+S7rqm/xVIQShw+RX25YD2ktgKxf8oTkO79qH
PRpMSXRIkXPfsOv9ZTw7xiMMCgZ7LC82S4omHyfGcmi4UTDfGQ0W1r0rZ18MM3DF0sNtoG2WTxOg
HyIJOz7rTYLQRTP2bidh/J0HyyyD12xsqmLFjTF85IQtcLZG1/J3YZT1hAMpGxrXT6pUbx3LAybd
4wTuYscioTBuPR5LrUB9MCI/PRIxd9rGvMtEa5VqtZMqZixHvCOB/GsfmybGOBSvLfFfzytyKG/U
R52vttvKoNlTbiYcg8zxQqeLIUkTIUPSVcY79VD2FkCkUvnsWJg4RhzccQEy0Ynji67GS0FxHz/x
C1omlic8bEff7BT2ufRWYZSdFkT+fVeSqFNtOeBIG7OmWwGLNwhSoQXUD4z5nSWDV1RYXG+9XqP+
/ib23msaCZjRcvs7t26Ys8haPHzlNE0FPI3TyGfuvl4HWHnHiqYIekobeXxKSH2qMyr5L45E58bK
TO/e86cKl30A7oUWVHs7Z6r5J379t0iVd9D45o48feBKND/KCT4wd45h73sFhNlQGBHRxYn/5+9a
kDR24DEv/wtUNXHAQsGf/IY3NhEpBDkMKMDdTvhfi2ZQ8SXXu3DCGbfHWeErM1Y000pNGDTrE8FX
+X/F5ie5rm/b+DK4Wx7rloN2f5vSll3gSlcT5Yxo1lotca+37nA35+hEdHMzoXeQ89qUm5B7hTuT
kFv6zF8Scob7+cHgdIDsNJsoFXkUl8vNZdAf9YvA94ECrjQm03+kqEu1+T85waDPjmL9Xq3EyM56
dqDNrLt32Hcc8XpP9QKjQjoo0k9l1FQe8V1lrGn3Bm+ghjRk0ZRUrO82rQyCvWQEnrQNDanqw1sE
f5ff5STyTz40+YgKpSzV+6oY7fguMD5jIu8Iwh4oN81ZeJQOp9vwdqFZNmZSsXo68ZwQ9wxEZlCl
qRviniqxutMt/tVYe47KpugJsNzph/dYQbmdChFvNMmy3hwu2lChSPlUsoK8itwZviHp3Ci/XcrQ
yq0VezUCY49DATyak/pNe5TGkMP17l/FXNDSyubahkP6O1MlO2490rlVQB3aBHsf1rCFG0EygHBa
fWl3ZMCbvE7KHEyH+vtZEV9BVlHFUc/8w5qiPG9iL8PaHwiz7QDOaclJkHyHxaVonWoQbcBlk9+a
sz15ZK+fXeiq/KQ7uK7okTw7hPNA/9VzDPIT+l6G/z7a1e3CNTc1Cgq4FPHXpVG3q7z850TlX+km
cJO30tOhJKbuijJxEF7LjD5jxyVK4tf20uk2x+j7yINdw2qYZZFKNVXmaQLnLOdZG4qfg7SD1etS
X4ZA5mUylp0DYmSVNaoHWrnqfj5dz18j+j2GlJKL2K6zVsAhJ31+lSR5fhXkToX4ZAG3M970f2fW
dnHr8fbFg/pNLHkG3H6QZHsLHRwV2D6oU3BiGvtGExi7PJzMJ2oab1RKl04GUSW+twqzb3DaOB+2
9T9rrtFXovm8qp48xTeuTRAn6i25Cz6AfA/I6YBVfl0+tqi+jNu6S9bUU6SFS/z1hhGUd1nv52Bn
WXHJX1vBC1K/4q1y+7/b/OEa2guG+U7ABHTesszPRiO+IOgnwhEB5NPIKphD7MOWoa8kpDDSqt6Q
mBP3/GVsLgpa2QRr4XI8SCYdRAVAvW8P8rX0b/htvWR7frquRUYeJtvBaKcsOz3IrlqPt0j+tUVc
mNKvJCtNLh+HIa5sUqLVE0u8MwnSACLvgDFGAGLQ2E0gHc5VZ+mo6W4Rva47r2Cs0+zlh+hdrO0+
6+nZpBpCd+YDENBAHqTTzdzzVcrI8C75PPA6XfTuiANaLqWjPe2U03IAEJPbEWAmi+J2GXXvosgf
5bF4eQ/5gMq9KemAKutifARadRZk9sYPslgQjF9oUjNm+e/Y9epYKSq68rwJfwVKy5JPwi5be2sq
Po1NAKUVwTWT1h+FTT9nd83LHLdcczr7fZ+QfNWlY7Er9W48n3L2A1VoT2wjHFPgtLVUPHUnMwOF
FVGZcctTzVCGEqhMxuXUznFMmG6GlGxHt1FDDfphynkujNrFe71RQkDO4paLdMtIrCB0LFhB4kqo
R3xod5iqXlNckcHYODaIoB9cDG7L0rjagPilYFtmjwKfAlAzSf3CDKrc5gjSh31fg5JrWKA+iLt3
Z8Vp8nXi7x5wZBhL9c4ttjoYyax4b9a+ZM525NkwXNLm2EfhFBqaxepOpv0XYV46xncdSam1Nlc4
8bRNRITUFR+rSPNErEGtNEQcHa6IMROkxlbkKcO53CBe8RoB9NuCUr/UVDKtya29Q3kOSy9Xq0bj
DErxZ1VCGDbXIj80GfLDtvxldNtiWteCViVbdNpZ4z5UuGNHhaWNf4rPEjUyuNgZpUGpcguStCWc
JvjNiQHHfZ2nu1yC05V13NwCgk/quX/3ou+rmeE2pK05vWIgWaN5WFZ7nxIERM7Kg4LDZv08Otxt
OqjesSBHnkCXeTb4qjTCOLvLuwl/LGbBavrH0f/AvMe/jGdZL/cgXOnPR5LaG3sOmftV3BSNhysu
p7d0JmocVyOGaAS6oUH5ubuem3K+xuZMzl1yjdCiiuOo3wWyB/47cdA+9lbFRgXdXvLpa7RCDOpo
WnCpSPJNIa5GJErZdzPtrto0zgxd6XSKvip8RUfQqSYl4bLBohnU2E/JG/+FhDJPwn62l1Vx7C7D
uGQV9DmNTdIEqtjjBxrSulLeaKi0cYJat2mTh/NFrtmMRFbg0bINw9A1E1PeHhCpgdW0y+uSLedW
qWKX7Bn/WRgsQP61adntSGWYvMve6K6wajF36yeZBINmX+62Z+3wJ59/FInWWHX9/jEjv70WtiN1
dLyecaVt+MlceToBI8ZaFQKV25kpwN/fHlzL4DbHJdJlPKscuq+UGdXOCCrmvjSUpe05eeZYe/4h
Hd7FfU0baEx8gmGk8I1PoMZ5KbUhD3uQwa+GyBddgmLbm+9sYZ2TTz/pRaW3RK4bMvpJqkrWEW+T
QsZHA5HGUiMv9hJP4pegr2jtVDfEDdkC8vOgRsrzxPtK++N2eENvjZL+/xPyv1K+ng4Nf0vtlH0a
FwB2xyqKmB1hSJ6KK4xH3cC7Je3QEei7iTJeKDnvutcn6HFU4ViSHocARg0rXydkUc4vqPn9uH7q
iGjvwGiYOEDvYT/Lgj7B5uweNhRnw9rpQ0kWqmQ+y5+QtBs4IE7AZqFZZsLY5hkV51XsA4w8y8+0
+KkDlwhRT0gA9lcLCktKqOVLq7//lkNxxwi6v/w19Qf9bdPKocn9vhHQJD67ImzbTnuujQPcWPlN
lSz8RYf1UaMvXDlVCQdCjH+Pn5QoBG0pq0xKp2QHUERY510XZGbCv+GrIapq56bxJHobNo2e0UNj
UOQPl09fYo+8OpOySneYQvorCcFUDL9/Tx/fdRJqhuzbm6G+x1G1/cBFLUFy78wou1D+dqq7lUKa
IGqHTqKyyczQxAc2AQSAUQ32mdrA2PcPE5wh9mqMybWjVaLIwUMtpdKblDwJS+8vFLiWl6g1UjYN
P7Kltvbny3k2Ufe94eveL3lkxH4OOUXo8tNXSxYrfzJisbb/Mjzi23Nyay1TV8KErzw/+7XsSr0r
yhwp30GTMqoO1Ljspv2yONvhDz0sGfCYMINR8a/lSGPjBw9t0lwQK2Stvn7F5ZRnLbyTYwPO+M2F
7hGvzZKGzYg88LAmNVWEhdPhVCwSq+b4a8hgyPfzRei7KlDiZIVbv4OPnN/iFKwntGNxIIiVvC3s
PHqxzYc3dw6TEZxFXL4bpY6CXwFRHXa55amSOj/flnyeRiKLdZzdW+uF9ptFe2MXPCneb4GQgotn
l+JMmpzyxnRGYHPGEdqDJAavCbYv4MexsXNXbypq7QmuPiD2kdt3LN8GmzyI60+t23l3+Gah1b6m
9OLtkZMo+C7CDdu8tuVh7maEJyAfHgg9knzYT94y9VhCuWxpq9lvcqdxJVLs/wYbfAqzV9Gifvim
AnpEWGIqTDs5dlyWp409BFcaSO2XaThObh5xjvytIRSiidiBwq7ctKAzJJRtVytSzEt0x0WvNphJ
Y9izt5a9wjU9r3sS8scIewiR5s6FdmNMR59ybTg3bqh0tmxYTNrdaDDsnUSsD9FBvITUXNS/clzF
DQuRf9QLaR+EKHK8k0dDtZaJ9teLYLnaht8Mrl7FJY0NCsNdQDiIkSkEPflhBquTFnkOE0HdWshL
S5HaKEATMli7LKDji391dDUfrkdzYZ+0PetXJ9qeKp2J+y1o8qaUUFM7k2HPYn5x5jRRPK5nuOrt
PD8PEs97bSoccQV+TIwTIMFhfVRI9dhkDsFL1q8tvj4uHSdguZi5b1RhXLJWxr9ly9HPuzpSpdCj
uhv0EKGcX62bLmOjweq6S+RyV47hpiHZl1zLNay9vqPwGxJl+az+GmtI7oEOlWkSegrcU1YtakCv
td1Vv9sxKTk6jALpQw2Vdl8ZvJyyfXfkOlu1MfdPhnlfWGuy0G4ZsiQWSWW0sG4fs1AfmM9jFDui
iXpL906cz4AGIW1mjv6woT066TZHb2nNa9bFps/B7ZZTSPQ2ZWpbS/cob06OLOX25Z2FwkPtKTMj
j2BOH7ZF5pOZ1IlJBpmhMRysCSYO35ZX/jBSDCnqV5uAAMCnkyKBQ8gk701NRIQyUW0eLuRSza5c
0arlKbhhAK0w43Rs6e6MO1WhFWHvQMnR2PqQrxaxsyo64T38gwbNKyCucB+CAWTQKLxAtsyJ2WwT
DS/d83ylqF6jsOXqKvD+IEzCJBFLpi9GM43AXC+4hlzBqw/OLvOQWRwAnx5gl1TXqEWvad4XcrH4
WXeRfsYargpPnmKJ3bYrpDv17GZasDhr03lTopv4Rcfv9kOvAXIfa3kP/LGgcV7DPIC6PRNYEypp
0jdvSaLI5oGTfEOfKjsZDWgFzioy9jfMeJpiRVGay4n1lwDmeqU8pozyuKb6z5W8f2TTjqUBzqnC
sNZVHHn5nGwqkH0RuaxGBPoLQpy72Jjz9TZoIC85qcH4x2m6Fnwu43s+x/kjKCb0CIZn2mge4YU2
KrORR/anZipxhXwYXQ+4yxEk4jtnK2xOcipbzJweFw1Gw4TFMYZZ1DtVoIXcFiZQZUkSPCCge1mo
HikeRU6y6Ke+Ttm1OSmbHzVtVlpQMNmKVQp0dPbrQb2UbxBZmFWFtOZPPg343/dFlLak/DVJnTcB
rJzfGTUpPgXe138MSRylSqorR2x3WgdRAWzDKs6xn8yDY1AUHQ1yRIWdb7Pes514aPJf1P0kmj+l
WwuHVfyIs8qg5hYq7v8XY3d3wodNcr9VXCwCoZ4t/9ozeVCQHDj/kZ9oP6mzSeRuHoNdZggL1jzM
5vfTglAjPrmaCDiOiSPrQnJQ6u/kfhmLDhOrFdFml1CV0GtupFWGhpR6S6aPhjJdJILhY8onIQHi
ArlcGlNqJ5qiN1b4e3OUODd9BXKKGb1fljkn0crFZdBmyNsxn8vsBSfmcbpGgnpnz/e59KxZ/uZp
8eswTBteYw6J3kS+avkUvt9q0lA5/zCQ8gyPyAks4qugkgnI+xhhaUsSK9Jm4vVfJUJfyis/5hM9
9bdnLX2Y5AVt7fkknOgVaBBq8dIJJh6T/fob9Z96ZJskaisALKYJObtjTtIQgR9bK+5WAOqUdyWV
k1iL0AdFg5QI0o44028AGojkoxyrbMDlOB2Gs+2DgVkc07t6NbU7JWf5dgJLfOpHU1I2/EZnC6co
kfyMiVINnDZagnyt1YMeYVON8yaW9ELqlIVopNIPRT83wbbqMH2asNK+3lZHog1mDgksuUKqA1c0
0yLftJLdr6thL7cdVZtZ94RbXCmLTdkfiOQqBKWPuGQ6GTYrXA4k2Doyno8Ai/VHTh/X8/eKWtnE
Fp2vR85+w9M7+agOLpJkYkT/NXD03b2AKpKGH86xAG3kdSFqTOv5Ms0xF2d+KfW5ZW5jW3DgLWsC
0ezrpa2WXGUYgmq+ix2uCf7erq7s69wAwlT257ltM7AteZMpuZ6rUVdkJiYVw6yHzBIIWV8i/pSA
E+UzCM74Tx2Tv8rxdUfzgFX/gmxFql/My93aQ+Kpxxw1cwwWebkix0M7eD0A/I7Boc5N6z3wAUAF
aKLbLi0BcwZftKe/2NeD6nB8AI0PUN1EGRPgbcjTQEhcWALJbXLDUG473rMAWeOZkquSyrRaFLdm
BG/JTDywtZlYcn4mAIDHNDaRBfrLQJMl27GMg15v+41SERcV3gA7xbnHdbWYvHXnocdacCYGUmZK
qd76H0mH/JT7yMcQYjgMAkgzLEXQRpL7eo3BTesHdqtGDtmMhhJaZdbeq/RDnE+X6oiG4uOVQfDO
UKNOGSqN9mBGcm6qhpVRrQ0a5UUFXh2VCDJSbBtg7KoPS60fae4q9J2lYXNzSBskMV4WxYcpXLGN
im1qkiOdi/MU2J3V1W/iL4MikJKV6aphbndBSDl9bdSGFhsIWCAkyq44JcQVlhldsULG5Av55bTA
e1LyET614wOp7K/UR7FrOdw7XU9IwZmrAxpvMoja10ONiwf9H7DohGA8nw0ayR7TBQNv8CHq7BYi
C0sk40wq/ubf1MUuO3L2eO3N5UcChz5z2Z10Gwvd4/1we59ssY03W9LxFYRqxPTLSCaDKCy/1SaA
iyHCHBbcTbs7KxAdkJvkn4MpHD1Vujljh0WrUtKffQTX/EZ34xIUcr0/qtRy4FHFzRF63tCu6m+9
PWqudwvxBXqEv5c/sInf3Fu8Tt2pBS7MxZ+sTOJL71uKfPYT9XsUtyM3wC8FTuKfPbyKhnlBlPr9
RnGxi1vwRbUhAvLV67uKnpGYqzcYq9MePcOGQRjM8z/C2ZA1YKKjDZg8CB6uRyzJXgmo0yaHnaEo
UVTsVP4tv2kdGou0cuIuX0kaisvzHEgCcHTF8Tg5Ff/numJ53XTNUU5VuvgfNaCulka7rDrKmbow
8rdwnHJSo8Ii1XuJicIpb7BBEy63SNNqIzDoYpd6DtaiVflYJh6AN3O0fJN/cPk0tVMJCXf7mHQQ
eoGg5uV9PxSWhduIUGmV/uYFGsHLMCaqPlAQmAj1xVYRkzjFL3uVVJbIKCGtVdj0hez+1CDlBGbY
ZzOLKXLlz1ORyrhEHZnrODryBIk/solhZ3LnOqx5I9QTN19Lyfs97bgp+Pf4Uehv8UR0DJ7XQOzu
6I4NFeQyZFfQmr1DDllMHnef+vIXfPNNHaxGFRwks6Q3ulVKSYB4mf0bswbzdd1fznb8AnLVHQUG
bcSRIPEIUEPYuwkWIkqNY/t03KKqUiXYZU8zxiLw451FO2BqnW82Qjz8TFxw4bS9l2YEN3LvmNaG
r2/StbeyG/oHcRh5dgdAoQfn0ipE0TkgL3amlnp+DXEDgT8k37i8d74+3leDMOEoaMul15Y5x9JC
6Q3sxgvasyrypTTSbunoc14JflWYedV8DM7AgmVY89g3Mwiqa8n/pdq/av23BQJkYZtyxePTx+bn
EN3arL80zIMXGVwVyHtWPQm9O1y6uCLjcmaERFifNj2UnGXLYI2cR4SWuoO45vXO52wD+3aNvOAd
uPp6haO+yHh5dUeU/I7SKsNRqnkUizanblg2rsnDGZ4MvR52kDGZR0tUTT2GvjjYoSuwO/idWaX2
6yRWhvcMeYKMi3MwmSDso4E83sE4YtHUe7BRp6GRaWlbFamWxKQXBqRy3y1E/YDVfge2xnwcVGsB
PAOfVaAsBw289iGcpBZciKJ4Phd7SqtTqhKCoQ2tU2T9Uih6HJaD70BeHcoYOiJdP8V/QaSP+jMW
/Clz8GXKKvcEfhmSkHTZqqm0jW0TXNQD65hezGkAGWsGUZc8mG23u1rAk292yhs9jyGqcXIlKQlS
4QA47VqV1LPTsLjk/ouNZCm37gMrPZidHMQm1Chc4iWjJWj+j2heUDhRbLpkd98bijkSMlcL02ns
o/FEG7kUE8FWnLZtlKkfGu3wa/Wc4jJSuqGO97SOU94qee4huAG0HDECM6ZE8iLAqAOHuuvbjP+A
n0x/aEb4FuH1dUZd55DEULQUvUKeEwMRMI3tCTmvM6d648RW6lt/nGoRWl8Vt460TF3RxsoyttyT
2i5liFiJ5g5dHy3EyaJ7QekMQpTgy1Rh0KcF0ujtgKzbyLuBxog497EPlGYy77GMltmB1QCjdMIa
A2MFKhWuOUl1TJRmmx3fO6whfWB/XgL6oJH+FW4qEPGKOAdGUJUONO1yheCEMUWSv7qd+orCJXVf
BeuSh6Jz/SnkAa2TSaEq+KiHUjaWqY4k/dLW/rSsFJqzZr93x8wDmCBPS7GakDhp5Lp1kZbPWF1J
sr755BSsHnQfMVt9970HbfnxVdSk45eolNwEENOTsaOIB+ae3gk9YMyqTly3IXNpaUGKLDupP3Wm
HCk618r7Ly1qlyEBegB6Wx8ZswWYUxORtfVLebv5vIgQSmFyHDKaAe6DR/lE+QErimbD40qT7XCr
/ybGSg+Pa1gpnJNlqsBricXo/ZQFKSYsAcCXcbfqmROiJN/59NfKtkeASv21iIYVcsH1/nija98B
UQB1pZ4lebwhYdFrJQxRaAKNaG7mEdwUUc+Yb1PbhYidLNWZ3+eZK2JyLkr4W8JZ7Gx0cFhwnOmQ
QZKuGmUl2U+kdUrEPF231uboEn5TDyiN3rU3ME/VmMwspnk1ahmLRIkXaf8A37JEXsum/bsjpsVM
jMTDByzxkhiqR45YHMBxyIKODaVjgtDGHXhg8p7t9yt4tFoh8SPNa5wBRUUQiJF6soIeQhY/83sH
vZbcQqIOD1NjR2iIhlP8+aM3pAVI6tB0pWvzmOAi8BKfZkJNUVIMncP/1mpzGe1p3bIO7xtXuWFC
gKu572/hB4xT0aMFp+fri68G9Bpg+wI7MS05vIrjRTR1C524EjGgkz6oAVxxWqVX5nX24uM0rakl
AMQ3NrDwvxuP7+8pnJldG6zWUmgRlG6m9pUMc4gIaG5o+z/C3xasN/P+g3KooVHiTKjtiBhPTfFJ
BiL/zIePREA9cLy5zZL4znFkaGUtVZyGNO+GLUjsfn30HCDIiMSBEiqxAxfRenx/j1LuC/N6nxhv
AqKFbSDXnb1j78cUZFBFoKf2Wa9pcIYaXhhJjw1UjPITHhGSZl0NFAPJalxAjeWH/AfG4uqLPL+W
1pG+MFuRe8baxZjAiT4k/k7pzoRJfWZLY4hz7nDRryG2blEcRXoNgZDMOYtpbC97dhZoKwe4a9o5
ZW/yRY1ut/1VL/ncg3nOIIOmk9trJQJ0EjPlGGOfDkkPz/XZUfT6rDVisefoe6ksacppSkqms190
1KjrM/A+MEHTEIAXpbRiciDjNhcUSJ8BbacZI1DJvf/iV6Entq4GZ3HQe/4a/xc1BSRh/jUSwNp/
mvdzmPHO36AoIfB4oU3VXw7u4OBxyRLTUh2gyDb7LZ1g8isEdvfSCQmKZRcZ11x85iofHjtstSr9
O9bsDK4Y5mhbGAM82ZQWa0EmV7fu4digi0VZDTzuKz5KCMGX0kfjxvFTpxcZTKV8wgHriCUS4WH/
T/ExmPOgoGUPiGyPIy+D+/HzebhagcB2oEIw5+cOBz5ST2UyqNfsocvi3OOByiuAnKBzHOnEWTCf
RxzFX9cQwcWHZ089mM+YLCuunwP1weNfxOIHEE4Xw3+5N77HPrT/bxvgMcoOhUpgajiuzf6zFJr5
oJuAApHhnekCvpmFWa+uwX5J/ihCQkMhi5C3MievgZiXnl0/BUCyrHrtRIBX3xKFjRUtdv2j1UkZ
3ML+3aWG5tQpKIKqvmQX5HMXmcMG4Rm3DhXLNW+iFxO1B3CB88lsoGctL8674ZJAyE9XyBvo8jOc
fkQB/NuAHfrkJfBm1J/t30yUO5wdh83BbvcqviCLfz5h+O4Kf6FhDrmJibaVxPk6SQ0nDPk00VxJ
aW/uYQ5tRpQNc7WfqvWGPj3z7BMP+0FGWHmRZzMd620Daok+k0hsdSxjD5+XJFa1NAR8yySaT94e
ZeTaCCNx0eqil4OGWxGsuv5auZ2NO7K1AA0cY7Yafr2uF7WCd+DobkqesOFkx1GNnZR0nuGd8jWa
TSPulLcIjt7M5URIIXz+wsf+Bfm+Z+jPke2w+0cmB6gCIoXoMg0tBMi78F2g8yseRBiXqHQfy8EZ
nQkZurw72OKkmQtC8meCaoGHB0x6Ufn0s/KjHawkqRlTzeu/tcpGVGCTZInGYE2kRzmYY/oNkcvh
VozKqC2N93NRtkj2McEq+t8llJbvp3/DWCez5ZLMdsa27r44/EbmKRtka4srZEL49sQIbheN9uK3
XFhD/h3Zg5N7E4rzF1oBRvCACOGvZAepbwwvl6ziXfWMRUQtkaU7OJ41JeT6APGewN73E00b3QCE
UbM6avNCDVye7SED5M7IQTM1Nbw1EvyLbfBMw1uXhJgml5BUwQ2v56P1phl8wPR6rkLLuPSaDJ2O
GuMl61w5Qyx5D65PhQloF9s6nLxatn6mlWWwZoxlSavgeOPCQeh2CJaD+3bZJYEODQx+rl/BG80k
bZP6RqUP3tgvSzthnDqaN/T4inzkCYYjnoHpN+HNJmwCB4cbS9cxHbYRPoMHZ/gTISaPP7F9j2Ux
b8rLoOnRQNfCplWPlmrAe995EC8nv/5GTNt1/u/WEKl0FXGZ6nIe4JuBE/INgkgVDh1uEqsDPqTO
mKbabfR1WDhS2+SUguSHvQ+5Kg+lr8T11PGBAt8qfR6LuQRp/WaRQre0aPo7HCxJfKKVE/DBTvbv
q+sIKWN3HCUSpzNpB9+O2A+yMz0PzaLHyPtRJ3h9IerDZZ54wWUqyRA2AiUPC9OqmMoAdnIBzA0m
ML5L9FVTI5fN34lhQXQCSSmJCSHUjIx0exiXojY1JQEmdMO90OMm/rCQ0OaSuA1bBSRMhz0oDbwv
kFSvh19ayWDYr5Dkzjxw29KT+77MNTu/+SwEOMpXqL4zGrqlWz0eySQNQf/a5eYJsBUX04WYDeWx
NIPzkEM7LORIaReu2Xr+P4s72tG0ibBjCcUFXPJVtqEg8lXQdNLQYEDRqnZ/EpnohR1sRXab44am
fUNQxqFWP3AsoLMrqMo4OkIuUIY9wqPLM9wts+k9NuUQ/7htSNEJd9NYBjHG8wWicQc0jhSe6vz3
fJ+0WVx1UkZy8eUG3uoYMUqIAoZsEKjk+kjygHMYEocVsZcA/sGFzUIUXgSRN/vt6tdug5Iuo04q
0cYNWSc7qxagh6gyTppBPOzQn65pfBlGCa9rA8G5k0rNmq982SuyDelXSronZj8AHdrR1h8cKVwu
HW5RR9OLADfJhWiWBn1W+NHWuNE0b+od5LNlJenf8ZmiL+LyR7ItlhLjQKaJBh7w9pclnpuoJFmJ
bc4vhxvJ8a4MjBg8JN8/zwr/V/I0ykDMLME4BO9KgCuTgXTnlJ1jU2WzUo4dnyY72+z8U/K75WVY
AzD3+JHkUYYfCJUEUAnZXsDbmP+YDgSLbkDDuPiBjz2+RQiDSv6TwhmcigbFacBQUPet4FhtlWYk
WeLcuQPXjbxWVLmOWAUQcKxodgftvP1ab6c5SdXzGAnL5asPl8EheLuUNzpWLRP2tmQ1w3HdvMvj
bLmcgY7xtz22klbbqJD6I06JppVVFCRLsZgd1UXIoscPKv1Gg/SlP8VhbXhXk2EEM3QUZsxHgUtC
5cc3iJfwRxYFCtPg3A4qAZofwLKYmzgkqcVA69mp8C6gv+Wnff9+bznKQv5FDNhpN7SUqgHI6HxY
sKMteSu2ZGEcV2bs+QJ0AyQdgYAoOnFI9eNZ3uZ45dSawhefSeiT2CvpSRL4Ma9qkAocOsaAszLq
csIJeKvj1rSwMsU+I8qBOUxIm9EIKVE3Nlai4oLwNmQ+euyegwOebGhtoPwWsvU7I+LVgS96JznD
lJ6A4/AnQyOMMM0jJUADffiXRTKJdKAFQO8YcurojM5CuJNBxxfaM1l6Mq1G8SaEnQU92SSrhdtJ
CLSHBAjqbv569pK7L5w55co20H1N5wI3quYufhHob+shHE8rvSsPc5H6Ecm6Y33djQQ3y5cFBgVx
cfdGkQrPeFRi3Hn1/YlFoTEysY84svzq4c/zMZ3KfhhDjB4xm9cZwlTXCm4NFFJ2nZrMWRRJCVIv
HxQLR58vi3bwNDZoxFlycSY0T1VZykSnbeuNxlPAcHM6psPsWjapL+RwFrcIVOFNXtXHr3f9uC6b
wr+vP2sX4hURxOjed4Q9qOZ17z/aXHiebJrotfZBh655rJCllXwrVGngmGyCpenanSVyaitRId8i
x81DbncVqI+lrC4SXkjfufyKAKVmmaf4mEnZ2pjMl87ba+UmVfGv+q6FcZk6x+zTTq3NE8B1NeK5
AEACPbThRxrfBBoBJP0XMueQAUgcVagfhn0aW3jzyxOjrx84FcVpuNxzCcTN+ouYntKNhQbEbMvQ
eGeJXNf42PuvssCZCHzEu2VUExOhTBMH7IQJKV1u2oZLRFYEggyjcIuwNfsIzVbStVgu6EQlx7nl
1QiATNvRFr+4TZL+rPCLQl4Pvdn7gsgfSkcTSpCHUX97rDXAmowpzlaoO1cEa/Inrp1v7wEaL1pT
QCUapX1CTM5/RS8ErrYmnrzVKQmp1s95f+IL/huQEhWEXdB0FgqtxQKKk1EX3RalojSmpNH7tQfd
HOwe75maEaWXUigjdivG12rA6aIzAG/OCXdunztA0R6s3+5ZkCvRRnoL2k8A5IoIWqtRltQF6xNK
f1rJnKuqBBtTenfj+XOW+Q6pt1rUffXmVT70yq6ZCskktnAeyxI+mHQGSb/vZYYJRNqgNfv/r+FK
nPglNBGmJQlO0MwVmZrs5RRJO+kGz87zOxD7i5ZFn9nMcmDOF/tXOrwVeg4kMsc+EwR7qdCIvVb2
kTA1JC3EhXIDofpRK0Sx4YULYfkrkA54Qn5erYHBiTUJEQrEqqcyrh5HwTm0NOLNzYhnJ2rIp1wn
Vs3k6MjJMQKxE7Udx15qjb624Ih+dYqIcXV0SknfXAjepQwLnx9kzS7q2BAuRz4mBqdnuAqIHfQD
aEjRKD4I6kD/zivkM7wfrmLyogAAvPCaNoMYkIeg7sOgWpxGYVYLnuyPnYI/YqBLUSNj1SWw8n1+
+MPfAPyWr2hNZRYVSMcTupKgSOfTOFcG+QK0tPh7A0Z8aQxSz+Bu4ZJhu+6kWCWKjFazW8fxs3ZV
Vt4UtrOJeyRPyQlLHINPlIc4tK3S7aMhMrTpCWftTuPBleQFPSwF8M1H21yfnZsO12fcnSe6m9kG
ojBqmFY3FQG7tiVyDsviaIFQCSjMmh4Eg+GwGbKwaZKHDDtWlOG+rLqqV+m6R3TD7GTLS6ylmvr9
6GxyaUFxVoeoWJW6tCp1BnYqvmBdLte1t+l8LT1zUb1KEsDumswzGhv256TH0fpx+p0bJDu6yrFh
LnHmqg3f9ekzLwDJYYxGZ/Mbq+gRmTxX+U72NxlwqPhMHNgZRjvgQkC8ClfoaQ79D9XIX8vqQqoW
LYntGqbJ+4aTk7hzxOEr3DvKvm/3kw4BnHfgJOrbgk05K2Ts1lYZN2BRvnb0v2bpXZty/rS+Xfol
EOSC48cEJfE+ziUXfh6qkA/ozqmab2eokA+YK8prVBnfSOahtkvCQfGceYaielQNI03WjKTglqtQ
lHwGBSQFBz1iQzA6LtNlHrbdFC/pweorEzw2NDiloZiXjfjyRSrNkH6wwBzwiV2SuMsip3joadJD
Z15ItoEMBJ8leCrpfDOP/6ddy5+3ck/LjJFXFOa2mvc/YNLyrJXfweUU9EWiEH2el1yWYi3REUr1
Ts73OSYCAdz+2ocQozNwKeaJADTcVvkX+dEexs8SRo2O4QmH2tD1rAzSB/CGEFKZhotSqh1dmsAo
JhEDyA+OpvRarJsdhwm9sstdmKwduPDqv/XomVO4PSlviyltmrt/6P3SO+rMyMeafmA6/kt08WhS
YKFGXBKEUvBVkEHR5vFPE6gtjca1CC7LQ9EsThOnpctqKU3VVQdAikXtkd7OlevFROrjgw3kpDut
NqZdCDBro6iN0FN2+aSqNta9VIzf0bJqObkCLLbHjqd8KZdI1fK/Rso212VkDcL4Rk2Gobb1dQ8E
+PafawOUc9eLAJDgTlXd6QO24bGAIuWm1Y0XQ+bpLSltJeV4X8P1dV4z2Knh4DgiedswBMy0zL+H
k+ESKx07XaONAVGeQW9lF1G5kMceNK4U8a90r/3ylGMEkvK7aI6iORKkJOVN2532g+t3GhCVSfXt
fgT3z3y2JLpCzDMsfPuBULLIHMO/wQgaEGKY6103T97qy7bZFb5NP1TahzYOHfvaPMfoQ+wPqGo+
35Ms+g4E+MwjbmB2Li4vvzV7LpZ/1mq3N3lnu1loGbDm/fQKGvjKzmUnOqlE2Zl6xSVFUvZ/dQMg
z8jlCS9JP0EWsXNSxacW/PYn7Dkdtgc7lDNY9OmAH4jcgcHV3VB7JOuJntG/yHKqqpe+jNBrYItS
J8lBhGbtwlYh1+vcWYnkxs3YjCD/jlkhr8hAkVg9QMXV2h9wdj2292PE8cV8P9+HUnjOxc2MORRv
8Wu2N7crRVDhmNwX9d8xTYM0xvRPhBrpnxCejL9rZ63tRLUwPrJeaRf3LaGSJilCWC93F/LFUs+0
ItqmM/jwFRgd+obho7ms6sgvlVK37UpS2rzu3sB1ZcmcN5Q7LrF+yd86fp2U8HnD/FyuLhoccubT
Js2oVLYg64OpaQgjfadFpSJ89L6yI+Gn9yOPSCc5za0v3LxguVN0rLIYOm76NNhRSCYOO5onUlfh
B2x56J8VTBFZEs9d3nTIZW5+822cb7SaEIuqqe5XlZZabVPDm177ZFtJQZzA78kk/GUx0qFYUL2M
ufAHAincO1vTutXjoMxiveIMCCDroK4WevH6/gNyJpFqG0DLxDG/N8fNO81eOY8Lg+hZhzYLEUHR
0kdaTxoT9Ci0Sea2NvsvxHWy+FUptlrjdn9dlFJyUuQkhn0Cujl0ZqPk2ExLclz4bhS592iP63AL
ni5OZpMLouyq891VxB1b6muzZSydQSnDa6dPznQX1NSBS7I7G+cloz2r1jasfWDQb2rX4mOmqwLG
x7eloCBeRb8PLK6Xv4Fee087bvn4969CbkqMvlZqexj9d+ROtlNR/Q+bXOo3D5YxkhB1Xe+ru+C6
myLAp2l0EVsCUJiEItzz9mhWp2nZVeG/sIYeyqyu8BVaYVckamZZij5Ns08+CxQI5zsSq8QtQed5
sxLOLUMwCgYMSacbBH+U1AnDHpn3vT61S3X9bQhX/Kckj80r2jfgbhauKnMToehMRzNfC6hPoft6
3TJPUKuWdpVPQ5wdRI+a9AgiJCjCNrHrtJsGnSnw2m/J5xNmQ3Y5c6RhlSLSK2jqt7ux4ZEym7/I
4t2wPKkKnJrkqEZ7/QKLRq3TiNA7MZcnOjROVCGbn8rIrFGlq2xloBEakSE8ju3NbZ9T7oOZW1es
hO2/eWynqgAXVALPwgno89Mikx1lzhrdSyJ/C6TNUVcfat56ThSnCSHtaYTJjpWvbr5mlouwrr/Z
ZMej4O1K/Oh7FPmJO0iHNp7OwW7YTsQ+8PWnpgeHh23+3NwP5OqV+TZ/JU0BejJuhRhyhYbIhWpU
uoNDbgU0jYY1ky6qo/vgMBcuKn+nTL/DsyxkHRaiebw6dZF2ZOR2xwZ3rtVLatnb2ysxTcpXNR3g
KBlWFmjx1estdsA8cp/CsfnO/xUtrM2J3/nEKqLN1PEk/qDT4qH6bMemWTgM9UCpGaydJm0rEvbx
VFejcmbyv/1lUlp4LLIkhxL7HvhPjzWRcSeg6XYlxx8JhWwNKy5//kOmOWe4INAVYSGsadb2+7OQ
bsK70rGOHpOXw6BocLF2d4t0sV5S/MgJrndhDpD+KmuY686XgUEM/r8m4qXP9b2IPNC0zvEOtY5Y
17bDCKIyMjuNivUhc/mPHNgraYm9umVsJYL5g1t/D8TOsGPJ0Hc2jACJhPzwczfXJwsTduN0wdtz
5D1/gakUKRJnATV7dhlimcHzqVpechRXDyJkcG/JsezqULfe6sjLiia0PsoramjLlFyhlw9Ihpin
ArQ84ApRwVbP9Kn0M8u4mmfyjRFp8QklzLs7u/QQ/T7zv7xLVJHNfsvjJek0uXAhvEikcF90vmLD
c8VLuDE6WbQVczwkDhMPMhWBHG/PLwNLzw8rliEp+k3geRty5Jgb4w2QBQCmYKkO7DtOg+btUErm
iv0VQHwhgjrjqYA3LyOkiLUCTSNaZqIC1NYDU5JFQ97bMLt45xbZXLWEv9D8Lg7lZW9HEHMgKwgj
/CqHHs929MlZkGjm85fLEzItpTZ0qh7QBJNnPIq4jLTA2wIqYK/kXEFUq3gO1fEOurOK8MVmxQma
B5vzHkDe6FlLB/WEIP2aG0iA2aBmpfg8/HQKbJd3N0xYip0pHur302puVJJFIpnwiI6Are6WOw8K
GHCbRpFg09KATkR9DVeKjoVQ8m/EgFS4L/Tw4XYXMYdaxsd5+l40XdnSRzD2BPgAmUCtgJAgQMcD
oUZJdVFdOqSyCVmQR1xMsOhOzm5V9kiERjTrscZ21MsxHVvhtu23Qm1dcl/MYDGrG90JQaD0mpd1
7o841o98o3VwAVsMGs48396XERqyiHyKqVOR53e8MQHuX433yr9+U7yxUJUOwDaIFr/hpl0SFEBb
n4OLTcT+5dxMhvtZLeildqnuctBoIegbOVWxDaT1hdkb+iMs2E1/dHBA88zYKbAZ7jNcHdmhKsdn
YUFunXfjLmPQNd/ZzbeuTrk1etan+R0IcGEyRU0vYlyJnFR5uuUUil20WEmyuGIkM/DKhTAXpnPY
jrJjxXKQWcnccAmlByI1MIuYkAqPlDmTtpz1omocdP7jslwXBgJhkWd4QX8gOBee1xqUKjU0gVP0
BHplKgSQtikSi5hF0mXaJ7Hc0h76l3D99woJjAqVJsgQF+NkrPcbmULACE/qO9UYFYV8D+auKIsD
erq4Wyu1IZbBCaCobWPxeW6Yuxr9ijxNyPsNxk3JEogW80m+yD6n7kfXd445TMvUQ0ORqRocdtH2
ws1v3ZNnq8Ui4bl9euJBCWjauB5cScDzjvZ0v3qZ2kLw0jhgpwiLYkPOXyRqiVVQfdAHVkyBxWg+
Agu3aZKda6Tssts10Sk2vwxnVD8xFvfYBxLuABaQM7Ln9qDNVN1wJVvSt8XmN+s0rbkhDWZdqaqz
QB4wk8hU9EELnEA2g3CU7GsXWyTjjU+RYkg0rwkLiQkVTRSI05WxG2k7usiasrgtlc0JIpHguZvS
mrBw1aqk0O2jrQc99C9/U/Z9axlrd+GcDNW4gaU9iwsAB+M+jshCe583EYS15LS5mWJSCot7LmyF
DXrJ0J0M2isLNTLHtpnu8bVteGyv4Sb5NCq5HzJBJSH1oRY6oOSnsG0yg7ixM8JJRiv+nkES2NS+
C2wq2Tn3pc84cxyXP7fbo60c0C/RO7kUgAFKSaeGpKpHGPxt/qGqMvA0i5/2NgXZuIFknC6kVcY6
/vIu59cUekji/lO0hTaaJz9QsPnek7r4vVBmWijLTqqC/VYelyH4W+fu1OiFqClJPssD7fwIuLSj
lIS5U4IzunSB0liCxs4WooROsAcNPuyDjq60WtjNXctgUdSQfxl6aAwncUsh7AQPcsvC+3XsIVNN
YSyBkgXxDb3a+vENHeQ05P/pK06BQvJ93rGLXUGKrAqW8ddyoDP/a6Z5NZN06B1vdBOJQWFkLP4X
LRRlTv6dG/8zeZrsbP3rEU47dUhVusFirCCBs0uciXBrfJstNjWpRWMTdqcPHZMtX5mKbCKxkH3t
uGI9Lg8HShDQww6y72NT9m3VLGtnJUF/J+Y/sYLhdS+5y5lDwz4zM6HzflgnD66gauh+VKePjIBV
yLz6v1DOBwUuX8KlWeM2eRY1tX+hHTOn+1Q//Ts8gfzVEfrpN7rRhNC/1TqyUtf1Vzt1cGnQw1Jw
T3cbHL0AQAa+Yb9sdPXUURsF21It3sPOoVSxOOWoXOJhlDjys8P9X+ayLH12Y82cO1VWL+7vtFN7
W09OZl0iCVcAWcxFjMKJCKbt4WTPGCJPUCVTEb4/DwZR3S3vnogqO8T2AaZJmwrjqk9zi3QdVeKT
BJn//aDwN3AaGzYr+4FVMQndgRQ/CQkEheqVgzFLJ/lrzxCpD/H3a4jqUBW2pxGHTb8bIJ/xIPyi
2GJDH5m6NaqMtVn56eTOzMJ4T4caFSSP8DZ/VJrj0pJtm0KGSC2gsZwyAknqMLteX8Bc3iDjQIlY
YzPtkMPqI0CZf9/uAf2eFy0sCFw1CBbjeSb1BqzHGpURJjM9i+e0y6i/JH4mHGhMzQ/pquweaen4
mxeHhZPADCVcodxKsimHxN71q8cyKNFp3CQWFDSjOdJDxuShbfsc3FpKTw7e+LJLrA3/EXjLOZfT
eggDKX4dceV1DTQf2kUAYNkcCB6ngHDn9GWws5V6sTjOyne6J/tjI2tIOJpJSn3PwVDegYaDFM0g
uYj5/e0F8eNl64TojbUUirVbwrs7loilzIp2yQPBOn5hb13AxWMmljFwkhgaUMbn8q87HQuFkzmY
bedKSv2uehOCyu0nDwb6v8U5WA3Gx7HqI03ia9dNquhYyicNUKEXt1qYJZRqYG2DmnMJDHgPEb1X
VaY/kbOtQG8suZ7VXnhchtkTd/q8czQEHj5g5pgVqQPutwSC0/M+ZbUXOVIRU4PVMfTIgWDVwf/o
5xGeVVhekRGjvpb2PwOUZcOWQBiMuCVw0uXeiuSMpyTmcmDSQKM465Di4sopFmJg797Nu5KpopVI
j3ySg4EtuZhmu5RHjKdyzUKgAF+xAyrshGC11nrKaCO574msFHpdh7rudpIQw1/WEbFqBv/F+Y80
PD0Ns+4S/pjA287u6a1ewGJpwq447eI22WS0bAF9TqFTHQks5GNgGNBnxZKrYIiBruGkT/t75oPc
5Obaq9qO85TmHPlfJfrERruaiVmugQJ7vrew89XdkLIsYRFbkqZVOtpq/X4aEUzTPQSICcTWTikh
8lycjmb9kkuXFtDkMwW7kk696DZ0Jl5ylECA9G0n+XRiBFnjjWSnj2/MFH1IF6l8zbYH0hjU04JG
VYtOwOnLmgXEmmuGWi2jpzdAFDelNqzWFbRGR1GS/igRY84dhA9bZ1+mmrISDDIhUP6cvvhjwv4u
gc0yx+ZT1pA5D7cjAwxM1wMv0fbG9mBGiXVggQPrV9MskWXaLQPT4E6hupKTHCM3AHCibk/ye9HZ
qVH4ol+gnNSzlyRPBXa3C9/dFcg76xmHhTunPuQHdVL1/elx05VwlCZ2WxS9nfyUu02omIdurYnS
HwKKpMnMq6Ql5VPpF9tFoessA/EnjoVlkifZww9ApGRZ3fQOjtdwA7J8zkbuZI+r/DcGQfBxG5Dd
JCedhwY6KhVfvHcXDY4ZncN08YKZZYyq7fTiyNGN1SiGXj+BVf+kn2jZYg7A0OjtqsEMzzqxfcy1
jwrG5v6HYV6NMIqv8QSa1PCRUSvHmahyyk5U4eKSY6AAus2yTOQN5MC1DiwzKW8hCzZrt5bTzAbY
9QC5s9Zo8lma6+K7j06t7TqL6r45PxNqAQMV9Xu/G9BjUk0iNfJdvZoroumMUTIGWiZSJhN+Myfs
rz8H9LlbhSGGQRwK9jcIpv2GLZMI+SWYCQNAknBVe5bkzVIPiedjo7e98gBZXMJa9CEZGwUX1Rd0
lgaZDxm34mNRil4ewwznulbus+nyNCVkiMRECCSebuYt2/mkq/iVJ+AQyVt3AVGl3ofaWWbIIEMJ
ud+RaTycmQiYUcHcsY8VZXSH0OCRnX9o9if3dc8KkRtDgSTihWf1QrS2liKh+KFg2vJrqzPw9CcO
2NfpYtrGNaySBNh7kkfIJl3UVWIQCv+8jT/9mRWdE7CWLcUOQombk+mAGFSoVd4nZ0DDOk9ZXlZ0
OI1yPkvvSV1QMz0kyEfuorznuU7mU1YdCnUBiGVcyS2Ub44JsxlYhqs/DxYFRD6yH3tcivxGEdJb
Uzfk0P205sQ2QqKPc6i66mhq05uXako+PCCnXFXEq91OO+sFNOGwEznI5f2xUvWhrjaeDv084DWt
bulmWztGN6yPf9Y6LZpfWLQxXe5Qfiz4cv/in/3Xwr5xDln9ZgcI59gob4Utx5vzwDVE/NxBi3vh
Gkk0FiCvZmi117RcwHg8pZbEz+18ix81G7u1eW+oxws5mZYR4PlrkCOqb0K3VAbaLAliySqgkE5F
n8pDfZGCdEUQMcVYKAN1iyDQN122PPCj6llmh5OQXWFTo/I1v8Bu/XlerV923zUHz/fnZmomJHl8
bWjDZOmSqY3i2nlqJSxyxLHuCC5EBjD8bBwhxN/6Z642N39jb0T/1tUo1fkFjI0ootilMYQOaFwJ
pMad9Y74+QMdDGUSv69ODFqbF368HZl0KdLvdVsmvGGX35166KAC8VNgY6GO6GMxL+jABYkZnCzr
PYTjj90bwAMZcrEApVfD56OTw2gWDnXqdqYCnzp8dp1qbveOLtwCGFdUZmGUAmTZQixGfd5AkFA3
4o31VTrqW9XJPnndvhMpgnEsTCyGekz3uxtjLL2MLiJVauasE9zMED5yKt/5iDofCuzYlUjnTFtn
N5pPWDvUYCA1mtbRuUsImQpk+u7sDuvU2oG5dkzNvY8kKV8a5m4WzddNz8oh7iOL64t68rRk9SJb
LxSVdUwXgkdvcob2M7Dg0PJRzJsyBSU7sTb4bCDnkmkkBYscEihZq/m57QhR+yNzAkmEXm8vVNgV
g0k6PSjXUc8ub3NFe6TXSeXQeGxBfEB4Xjg35uKWgEai+qWpVnLbgagQ9RnRlVA9N/2ry6KJgVoP
GJU3KeOmugaoZCQYpwpGlQnBz2iMv5ejzB1bnU4tSRm7CbNXATgSQ+uiZRhfv8F8IdU6vftS4hx5
MtMQut7Spqz1AyXqJG2A2o3vZukkLXLXtgIjRS6b7JaLPNyzwKfnQ+JABsNahkNV+SE4wd2GN5mC
WxJCIkd+a2rLVFv27/6P+fE6WZ02P3u5pP+Hq2gRAgPZHSK4MtnJ2XtBiUKhz+F9ksp3C6rF8NZN
2fVJBdFBltoSDAlWgHFIcX2d96SNmrtXp9S89VaeBx2CYL4Sm8iyPNce5IqF86Ri27iGxDlxPcRj
A/dqcRybszcpFUNKajfQYWy6n9HS3CvFZ1B6pw6gAKE3ECqQeLWucBkxrQU6gluwWuutsAkPh3/G
rvM7tbRGYTi6eEQUeZgvGeGzyPoLMdE+Wo4t9tbh4+S4CU+qtcs8zYbwC7iGfggfog/qpHYSfJmt
KjWDfhJNzlQ+QjsKbgRF749Cwj8cVARmvJRXN4k4xMKpA1p067SaG2e1JaZePxfuqBW33pEfZzXU
erE4YyQ+O/E8hGsbR8QLXRdL6nytC98apHSWp/Dq3HydGxf7koHIfzDm9K7EQGsJhn8rlz5YFqAI
+AWHWBE95SDqrsPbppkJ+v0ZeGv9sr4R9oEyxMsYATBUwQpVz8MJwYAwYqQWbP59WRTLGKm0DEz/
9Fvb6/V5QtR8eB8inacCKiuXEVAKdw9jK/fDCNciUIIaxT9JJtkiF6QZrILo3UBSgB8yPRi2orDO
CvInCCvGVT4ek056zdUlh0s5Lv8nHALHgzUNwc8LsmocRyXOi5jz442i/YxOXElfuhoCF/Gvmwwn
LcArE2CvZr5O6OnJXQ2kWLg7koW7Vmau7fjSYrmKJVLQWPbhzfHtWFodQ9JKZINHYSQRsSBd/mYn
/E4VSs1gopVSl05KNr+I8C0669fsE7t3O5wOk49W4G64a30Ev6wwzYcHTTjt4JmpxfXXFb9LmNzb
vEMtov5iu9FZ7+yo/7f1l3sFsGvn7kYqTDvHSSrUdkpc2cGgjqXSOvG3/QEvZXwXbbqcQdxtCjUQ
/q+u4EedDq+V1cOKD+sWDNZ58L9vi2GLe16sJ3u7k37hNrQbeCPWmyJA7kBWX+w9iRaMynPIKIQ6
pwJXY+RRN0ryvqu/nGBr1aQoNZl2GP/NKFRRPAIMkEGpOxDSnTUAzzS779m89tFgChVLb5ZT2QIh
js4SxTTFitve2gZpsaQO+uik3F7mrf77L2myh6Gjo06hVOsoB3y+F6zntstU05mMcMsJU6p99mjC
GGwg+nF4xlU94fTibl65szaRy3OwvrMNJcCjYZoS5INNCYgCZOyey6ZqTdNzcWY3M0Pv463RT9yp
RuPQeU9tlkDhdYtOanZR7Hh3i/d9mUFpzScyQ/jgGO9k0GqQ90UVkeznFAjzoZN6RNof1EQGH3wg
gHbSlnjMdykzTgGj0tF8KjJiXI1xEBaA7YOakFesUV7i5wbj8eL4BZ8B5r/PVJqg8dppPoDsLl9q
bEz7KP1/nM5RIjRBQDWW/iZQCRI4HLRzwCX+m7Rn7N2Fv/HmF0RCTXb/UcTxC2ix24pN7snNv+8o
bpOdGAQhbbgPSVOR+BKKBoSO6ktmoSspD1K7qFE+IJ1SPvtnSqK4HXvlN0IC5rgdjRxn00NXdrF9
ShpIvzWEoDfu2OpBWWcc1ZWiZHg5xAwKlGiolDF2yRVag4N5UVYud+uN1roTX0UOQcdK1YQPDqXy
iLcTktwyzE9gbjwoGxKKcfzNdxGLUQqUHF9eiZWDg4zaehigKDKsn2Y78mi9lykAJ8XtRcuoTpMy
4DJM0ssstQt0AA4RYcP1TSIP99flqnxcS3HYcRJcgWDMtE50JJWto0PCLFMqXifSDlPysqUlroi2
9ysthqY9UrImlgcAsFsfeAQqXO+CYXE10XKqF1Q9Xfn8wA210WZqfdQE+5EVFzLWVx6QCE0FwT0h
D1//7aYr0dsVZwqMcs3WHEsiRVHmocrftgNDLxOSuNCAwDubh0FYO/SP+N8qMjcuL3PvEhjH6eRp
VFLDPf08IfrPWgLuZNGuFmIGIChBYeQlp/tArBrKqejd3O9MiQRomFJT/nGN8o3eWoZG0yAhhZ4O
cO5zHXCfj+Jbq7MkU57yBMG3ELWRN95YV/q/OspDQSNrQSNFqWN23wcl6PGDLgmuJlZsj8OcYVGj
ceMjhkcQLmzfkWOml4zqrEfO1ZVx2cK1PxU8u8BI9lCInq1yuKS7R11iKTijXrdmSCBnhgWv6aQJ
tmBWURX8vBPxqgYwywG1PUa2WpTv9O8ctxeZGgYGY8c6SNnDsCjTE2sYUhKbJ07N0hGtqF9K2Rqh
dw7xBkb8CTprUU/uQ+wwIrMzjl9oetN0DZYWyP4KjMKEoabfOfuRpB01//nvSm+/XOuxTxU4HT05
QY6L9Kf2N69IBsgdDuWkSCwq7wBmmy3xcA8vM+GUYWJgSXM3wooEhFirTIefeSqTgf7Xg8jZdeBQ
9lx/JrhG++cUB7icgpQbhxQtRPWg0Ebgdz5Nsxpyggq/p/3DwYaMMXgL9gNGsJrZe4J6fVOTVb7L
THGIs24kK0GxozGXVdyuBEwG0mNiW/Yc43/frReTlNa9JKPU9rIotT5sBCAjVYGAmGgWeRz3NU5/
aHetQ1fOWV9rE6ddt+5J2uMH9Si+SQm5G2za9Q7DhwFpL6Ychc9pUnLcJJqLlTHLdQ3a3xXK7CCW
b8RxJ994TgAlb+SKIzfVuMj0JwZp/CmDWwvy2Le0EdojJL/VzOvjp+aTkDhZ4WzsS4F0Wj68AxsE
xbYR7ba6E+hYu8os5A++fldWDHI3mbp/uRxy8+g4HOFq3k+CCKNAXBDPbj2VQh1H4IZtxyr8WRU4
yXhVXs10UEfei7Fdn+pOZXq8CQLB0Zbvca3aAqPen8jIWvses7yL8EojrnKSVFAc5FERGAmXXVFZ
LuN6khtAucXWsQBmShqGdt8kG8eh84QViB1udyHzTg1cLKJsY4GFJJJZ0Iuzpz4GA3yeVHkA47Hc
CgEtNqRnXl7gS2Hj3uu26NoJ0cZD3slUXq0GBQXMnTBdZvmzHotHrYfCUP51XI1ngouf8M9WksLA
J9MYNQFC1cQbHpg0g8rtYnlWVUtzQ3j9TV+ISQNZnNL6DL581kHNUs62TvnfoCAw4dq/CSsEANOx
TSA4BVslXigiupLbnTmqTo0NejDnjvJ5Orx1FXmCtMww1cUJiqyO2RwBfP0tVDQmcVGLJinNTaPw
hY/xZG9zwd0Jt4EaLd53VbigmfQuqQ2nzq1GhZZmwd9lTgYm60aN8XwtVFR5aoVSoeqo2g+E8n3y
OpfTfsx7z51HwhFfCmdcIQ/im8FWFEIvefll1/9aoXrIYmxn+tk24JYDUXwtjgumn+Xs2JlKVZQx
YxDZn2yFs8AZWalCA4dx7G/73eb7KvhjtQBBoOVqQQ8oyIItPKumKcEG4feUN18km8yxI+0OKMHw
y3OhHKmqKd6NsM7Bfyv2Sz9bp95ypw9tX2bVUjQpRveAvcIiT3I5+otgAWA55yp4g+oX2+BNUcH1
9RknRG1h9z+9o1jEbIg2vXi0DEck2EPwDHSmGHvw+dtUrz/gH+/9eoU1j9J5PMk9cMWDPUPIWfgm
kEnVTI9XR1AO/o1Gk/RICYtcREL2lJ42t7EoniUm9dNAIuty0WDq7rbKSsXIOdH0jUTYS3iQiLkS
cMVhLpVQ9vIChNY02+KMvv0wExqqjmsLVZvl3yl30YcVEJhKaXxhYMqHL2mlaEGF+sNNozLW13Af
ZXYbGieWl9uChVHvPc/W1HFVOFCeBcBnUtcbnj8BK6hfAHXgn3bDjN/oB3Ua3hVfYLi3RDGqcjx2
bKz+bMXbrJHbvw8FPB6m0NNiAjrVXNxcdPQqLxLWVXazA9W6Vctss4rhMrlAirvBmlHWkcKVkQ9s
I8zx+uXqOKmSPn/+Gjv0PA/0cZcJl6Gy8tuz+F7XWngZlPIFTroXQIu5k8WyJZ4V5BZ1nl+RMkCp
oA+q+npwiFHpZ8qnricw7cP8u2MrLMdZMCP/Ya8088BbeEE/ah2vKwuV7K1eZiMPWULseG+GO/zO
Yb0MVQlWNiOAL5yD7AMhaLdNidD6LpJQPBIoyvo6pabfzvQL4FonSeoQZShJqp+wVQ0z5w24H+lQ
DfMqS6ZtPKKnvXGtZmYBUI9rneALAZ7n4EMIg8G9isn54NuOrSmhviHwpBlyA7T3zsty3/fQDJRY
vm4spwu1h5Hx/pnGakFOputdfFfSE5xTStWRTekCviQUliiOZsVBIs57Hzg5UUeynpfRkqIDO+1q
g1kpExvqOz9DDPtzgHBvl9nDfBaOgRPC71T3iwjIkQu+v28nyEp4eHC+5xa76Q7Gjmx1/RF4/YKv
M06WibM5nFyDvUMmZfrgkAYsqqCWG2+Eixdn5nPNUebofMqliM+vuHtafhvIH25XE92onO2enf7u
VQVmZWtN4v0EYhXTo4JjLc9BUfnaB9rX1M77PEaROAKIL731wkIPlC/pdDxm/PTz+mCXXPMUouOh
HFc10Iveso/bX4i7R1Gv0mQA30VIIy7U3nmGqvieWeX6jMsRayfxyzIDtho4dWlkVv8oqEeNgbaN
VpqUbEYTAG3b09YN2ZJwaCmPpWL0DxEnaKa4tSEcdNgd8lFfeghtlYbxk/B0R01OYUdsAyEt3fjU
4zsbxk/lzA/7Y5DAGxkUK6aJB6skhNZQ1POFMIMo3Tszbk/XvW4QCnG8N2+eWt9MUtnz5v6O4bD7
SsZfIr/CxxjX47pPudViMBTQF9OnnviK4qonVALHqPx6UlH0UTUAw3FG5cT2UyKj63hk/ZXUpK+d
zjluzhs5CY/5SfhdviRGrQTGmxTJLaW9/nv8LXk07mRdPyqsc8f3S97mqugpmjS7jwRiHId+ptL2
+/LFkGrvFy3xzCHJubpgHBsMRw86RSp2pqsIKJPPwu+1F6FmeiygGVqx2vm9G7yZ7vNcz5brTvao
WfvCwziwlWLAgK/48qQf8PE9D42BlU1S/1qK7Ya+Zp7te6yNIvM+bq4fW0xhOrgiTHBPnN0Rwz54
ayVVuNw32VjXxj4cCFT7Lhopqq2KR1WSM01PM8b/7ACGFHQKVhEp5deXf8rnZnwiIVHVS33sxCw9
m6meIYyXPtCc+VsOPBscMQbAiq83ujchkODtbf/hMJgA9fwdm8sR6+9gD6VXh9wHxeFmX46muTSH
VvEFtSE+sy3dq5e503sJH1HN3GsHjcaYZyuYswOUKbF8fgZix3NjBGFZpNj+DQKAFgdjy60jAk11
ulXsohipOHeHfM9cLUemGOUEdPW5Ek5OrYI8vQnhQYzx0AaupZb96Z5CDLSqxgW7iJ6QzFzLrf2r
7tktax9YbLWdjJ8v1jfd2p/arnL7ZvT8vpm00Nj7czQylVGKkmuj9F0ENA39PTtZvvtff2ZDTeB7
EkmeHWyptDl819JKxRUM1TWzmzx5JIXdwFuXRJ72vsXT6GBSXOaq5np+ad/97xUqDG1V//hvrwFE
6KiX9x/f8AEj1sEUh130kg2S8lFb2RKZOl46rH9rvrzmGbvbVzIOZFOLCptkK8VgBCCY8oAcVeFz
Emu3TsrCKy/4c6POjg8C1ddWFNVpz4gvG9EWQRStIkDlhiYIHrXGK+AlTEHKdsAt7I0TBC/Zm3IL
ebYwYjhFuc+h8eQB6w8ZMbZzbnnrPDq0RpMAHkx0FdA++yE4Hz052hPQESk15Yl81xz4keAdy2CP
Qb1Lk0fwVwf3GQS19ggvjbsCHB9t46TdnxPJ0FMPxxZQKjmtMBMZ8z/c9bVJ/6+W9Y72q25R8usR
wLnmQAPkyfY9OlLoifYwtoIDvEWd1e/Hj7ex+wgWvLG5AG0xUhk0eAOFUF/1AkI/+TLzn6nlF3tR
HHlzpgQwzw7KrhghQ+NYTQmr28bN9U3L9vp1+bU2aWpsLRaL70mnl30qaQj2hEZMoAg/57F0sCA2
8OZ6uTMjFBB6sRxEnfJ8D+cuewi1unnU9mRwpJ7bvcwAitC9eKLy15zzuVlHcPhIa/aAFFqX4CjG
92HRkkwg+B2hraFVxPqvqkf7oW+N/ImdMyBjHcxEQr0cvo4ISz++GhUCC+JbBbrSeizwK7dxqd/v
GDUmXcCkArdd72cnTD/H5M4z34aghqJ7mHiljvxgACHdjzrwpFUStYtjIWQo7wdSfEQp97IEo68W
SgxVb/iUKp3IndZP0QZn8TJq5fEWZeXXbBsrwFAqtfgTO2tSE2zAbNBrE5PyM0xlEzFQO+vMVEwE
eGWNxjO7tBiRZh7Arhat/ZwEymJ1mpDNpXOrrG2Bc9LX0YGDQScdD+LSXUYuWMyvrwlBceBMol2/
9uLx3/urLcEjzB3PuIuQ3lGN6hl02BtiUJQywn01ZgXEllwqEjoBWgHOuC9IPYgsyj+9tns1Kmr6
2Hm4jVQWIsr5VHr+OfAX2G9ZPaMQ5ZV7DnoSovrvWRaE9ojJDTfz5TN4+z0/TdSmgxCX9Fx6Pmtf
17B5Q0TdVgO8S+8xOYVRmfNbolJg9XYkAwxiKhM1wP8aCCRAb/ntrdfKjxWeOgSSDNoIV2/A3aJ8
GSOAvOhdVig4Kqom95fCflnNAQ446YeBcvX0CbB8RJDy8FrXSin6nQpKkjr/3ID41zxr7XEqT95g
49U61l2zy711kBz+Zuy+6RT/tkZJTKmiv6Thmrf01YEDSqYTzp9I6QP9bmFzLHH3RbFC3cnj2+Xb
ASPb0tRUzYXypdlet/KB5OzOkSZstO5GbTalQk0Ru6PejaBM1BvXA/sngqeMDSHPiWhKWI42U5Mi
CoDJsVmBD7O6sSoqGCA/5WMuK2OslHYFo3Sc+S5PIj90LXh0jGN30p8TTojex6JW9GZ3t/pHm822
KdPWApQLuMr9BO3IThI9NVuRaX5bXvoLXRTwLCznv79d2eIR/J6K3mzjnjkztQKH7QasAXCVpsnt
rxSdJGOg1yk+YZHOXd7sTEbP5Ju7/X99UIN7uEzxjnRDgLCBFV4QneG2N9gXOZ7iKQtEurToH5E+
DJmQqm/YGGcfFpLSiBIaIP429YiveIfsq3BmbBZIwRsTZLgGGYKbfmpEfPHxm8GNjT/m9uKQEDeS
g7FXkDLFVbiqe3ZUdVMPWBZHNDz6eF4euCYKrqJHD0JYpbm/DEEElx8ADnlIBzhE6vM/LjfNYp5K
hAzhMsLkRQSsQKIBo9nn5C7KbvZiwzdKZp2SUnraRiEhPp7LEUd4F5OZYP0RLU5qCj1aifIoU1LW
Qxu53mkXlhaARasHBq+lQXWv3VpoSwS7EdbKnj6L1Itlh1+psLrAbQ1UyPVJlp7hfe6IHY/+qf3w
VT5ZHd8sNK+XaXvdiw+VBVoNOqJbBfFhx2jVG+8TEXukrOEoYOM45S0w/AGs7thdvhLVR9wFYB56
9TWPURSz3eNXYCJxNY9zXpXbweyqXQcOBb7Nrj3n/cZiC2lRKpYyp3UCw3Q33joPQVCEmDGIerfr
jJGQEItUM2yTzWb7otC9F7ndLqVyC+nF4zn5Z6IvtW1+Ti5jzFWv6RIpslaIkxnB2MmjHxviUHaK
kVght7WFkkTJ7VtncFg/GEk/g/qTEmwpGDdL7SREY3Lwa4AHto+xPueuTKg+pCtZeeWvTUT1SGPf
JGSxCpNuZBuoyVv7nnzqVN/cUGIpqsism+8y8oGo939UznPL55PLULPForUuWgoNxqkxIWvxflWB
qYMdm+i5gtFmUOHjMKwN9gXCPzFagaXxOtH58+9qFewMaYFzBzJvXuWQQimHcoZ0QPu0fj97cfPw
/wtxVkRud1HjT7w9f4kEh6NhmrcG6ZJpRJ9130OHrNIzuxpeIOASzYcJltHY6787LIk+plY0WS4F
Exk1k/WmahhpgSx4JB5hiv7CU2FQK42T2JV8rprzc3p/PPwDiQALtHpBIvZXWJjhn0S3Bd3KpSDB
EcS5Us2rDuym2KBOI4Gm3G3W81YZmNYYINNg7gQj8lhs08EcA7i7v95ktNECw+YSlbArc4TTt8ZM
OT4IeBD5v1meW4/YI2EaZ+fAkWE/D2YvhsAWliqiEgZSsr0I97kXSCQPNt/6wuJ2aG0zcp0RUDhK
M9xcmZROgOuh6CldbelGycg7oITqL0oSPrcHNO1z3Db2SINF+1GJbU1nLrDuJXNxAgB2ZLjzSQrD
bbxT5qvgbj/EVNFOnWZCGXMrUJ4OrW8bfXv2tV7V50WfEA3eiWuvf0SE06md4kSea7/Zc+uknmaC
UJREh9FOVAXsTSTeLjZM1DWK89nR2a/Bj0zvdNx41fRJQRBFf8cEk9QLPbnktMlTSVER2/th30eQ
hGpaQN/JQMyI02PthFaEw0hqby4ov8ogPPsYH7/cPQcFodMMhTcBsgUOtgJuaOJHl2o8Yicya+hD
QgpoGaX4pT3AdJiEw9rvD4065OsXqgoyfCCzjx1wpXBkCuUP42yv/PTFW9B+EVrX0QjvGduEWiSt
M7V19Q8UhuejVG0Co4tdwQ0WQuHmhYS7+7iJOojgA+bLYCxSaW1vKKC/sJ+fg+3ty7nZeNgBOF4H
+vQBXJfnq3VFFbR+OtGN08U6RBhVDlPxmzQ2KRAaSFpH1T1VaC1Q1ODC304hBnNXdsW6bsEPVZ2u
2bf06/Bxzi9PGPvTzZPIWBNupiUTpHxYXEr7xeDAyaQhoyadsfUDvSVRIXL6mhsReoM5UoRva+6u
F06aoVmzpt19fkib369sYJaODNMfaxdL2JrPV5tgC+M4C+nRM+hkM7Nn0OAicRRcwf/nGPSBqDfH
h6sVbt2r0FdiOwKti0EDZh2zDTPbl66OpwBcHqtorSVc2pPEkoA1MyxtZq7nlBCAghK3UbcbMzjR
/gBTUJeKbjj7UlVVCQtUNImqjijmrDCL4+pzDs0SFGExay5b/ub84KNBJs6/dG4LOvBryd9Xl4cj
rq81CBU0KyDrsaxLXLbzRavl7FXjxvFMXNCzk2U2e6mzc2eAphWnmKCm7zJgVTJ7mOAAapNKZnXR
73c0vNM9adJaZx6IvV1T1bgnKSV+fNPsBACsDdxyRM9Kg7XZQ838xlHVX3CtAU+LEP5spUBYRwsN
1/dGl6DQX7wcuuLqwKRgk86t7wgsusCL/bbXB/HHniHqAQ6O16bR6+LAHFqm6CS8HDveV9KtYP1Y
DnE+Fsi7RQUtQ5bFhFBVDgEKz/gLoIsBkjBkJn9RSI/N+Au3mLWYe6IPC+WrrfSizF1oJIYRDXRD
Oh9cy9W+3qzRWbaA8koPXlOjTyKl1R+u4vgzASXwHppi2nc+EFiQVV9jyMl6eZx3CBZJRSuZ9p/4
1s6Wtcd/1QxsSFf7Y+CO1P5RmhusGOJ6WpDOI55S/k2X1JfQ0HfRnHShZz7C97bF3NIjdlvaWZ/8
s3slExy8OjdwKo1g4BGCzsuZoBrQvRqWe3Gz4mDeF/JaRdK15wJRrAHlqq9V2kz6LyFHmVWj38ee
dBthNqTcAawXoCi/SofAmqQpayNRTd84/Wf1eRoJs1CczrIP448lbFp4OVcVGKIQxq/VSBqWOTFK
vdupeUDqaOy47fYPzSVPIlSE6RTciPxFpd+3WdtkGW/wskz6wobrovWTzHZNc+BVriOcyENoy+dT
EaKk1lVj4OTqzMMbt/ogweGDp6RTO5HnywSITS2ZqRQTsGJAP5UK5RX4Z9PDyK32V7UmPUWyJeCY
yDw+oDwyOeY3Poq/mwLZ8GVWKHGwIu14GF2niArow3CYOEElb9xIGUUSBIle50dwUe+kHY0eprMC
6y12BDA9TfQA3ozbEJOElIL6pL294XMKYBhKj15uWA2uLu5qtqiX/Aa29YgQn2taH8v0bNRxWHMe
rGvl7R0IR0/LOttVQuiIbK4R7xj1IBFC3fMtia5NF0wKPfVxKQ7cLEyyjHe9mE02RND3QAum+B1V
PKpyO4AsWyzTabO8vcL+D9klUtp9yOSXUBdzn/eF+L+xFS4pzoMmn5x2UInfVdF5lSumQ27WQ0ls
NQrvU5xDNU8CS35pmGYNztRYz5FABqdevAzwkdqSLy+F1lCbd/OGzpJUT6Dr8xq6HPUxBj3B8/zp
K2GUzUztUAvXOLa6Em57nlAEMOEt8SWm2/Q5HSp/kaNbrkn95+Ht+YNukfc0kAEmWnX9J1GRxHTW
65lCB13gVrVKkuAuJNwB6XUscsQn6tPlS9NiYiT2l6zOd9NGAJA6CZEweWjtpzSLhdyPOYHtbtTM
DC8jXm5dt5qeTDCeOT7ypvvoWnEraXvyz3WapVEUKLUbEjCFguURXxW9tIKyZhImEFOloyOhMmLy
82bSav0TsrToJ8/o4qfJo2k9pN822ph/JeyxL5DeDbtZrKQRoNZ9/oW/lKUSTCKPdQpA37ALneH0
kRjDfG2/gsW1rvrF6E23A517/If8sEsJIhThRCLILec5qjWFGeUH8OWTnnsJFVCu+GJRWvgzQFmb
XuBGbm1MS4/6ZD9m6Prq99xW7rnsWSRyX9cUL/0HuE70zKymhxNBW7CO1+yf8aMFchVTy3Mp8ppa
1N+eIprVEFKiZQ6lSgCKLeUK/vzNZGx4ynNMcP4et8xolfI3geaJdyYKHNkPkHkFBjSzVX1g1PlB
+mjGb1rHQsTrtNAFkfhBHnBpziCNnpxnILY23ufdFu4JoV8Vcxap2G4v0c3zRZGkfIq+MNt8MhQ7
Taj4TUwED5pH3YHLfHWZorkjJSsIE2eShNBmhkwaT4o8oJ9otmTOl86B51A65YrV5eUkHQJ9TAm7
GsP8Ag+JL94bLv+kZA7gLb+YNfcBZGFwJXYfG0o9medcjsoxt6V1Vh1gtGOJUn2d35JwjrGynkc4
7iTOaKBEtkrJ/sbxmbYgE6pxu1jt5/JMTkTDXDdUpS8Ri/1xfjkaoz1/51hAsuDBNCCIMGLJjlLS
cBbLj3ynGfRv3iH4b3s6zr/mTbdFv7W6+EaIr5rSommswsMVG1HfEZdoMLzcEbeEA7Ohyn+flU0O
ynibLsIXfU96fzMhSypVmQYE8tHFj9lcqzl3hz2Hb8bMQIOLZmBPoAQOJ7xmk97LwdXh/WVIstA6
RGnPq+gRnUi2IlMu9MDv+qh1CLcY6voDUFMCr1jAVoHHIY/RQ3cNL4zLK4iiRsSY1g/MTYrkHpH8
US7gGZh2J2KNU2wVXdLMnJsAHMh4vX6S75rRhTQq+UqFEIvTWmgqxuMYJHfiDKQeNRnWLgC+p9Dd
p2Yn0HF6090N3k2gKimUlXkjO+pptdiVu3unMh4HRYKFvFYYsLvQSg7VH42kiVDkiFugZiwFHf9A
kpkASZdStAP5LLRjGQ4NzZD37MmI9vAm4/VH+vFtONLxk6aEWvyVycSixIW2VLrETArYFVUB/Pk/
o18w5nd9qN30FODEghGoX0T/ERvWbRb8Sbri2y8pf8VDAiNCYcc1oACQ1qrKMtpQmeJnPYJR4ToS
P/iK153mOF/WIqZ4LGgmj4XiYatP7jTLnQhFslmtwttyiNar8TpS/fUnI+cCfqXSqD4437Z0EXFt
fbbqROOV6dVYivCTP8OzKDvaYoyjKsqHmKMycBjTl7iST9a2BLxyGFK5L3WDy9rG2pMtaeylQeaY
5N/vgPqw2hkCJLWM4V5yYiQ3DGanloh+/rVKsIIiNZMV5fxc4VdpOe4pprlS5uzC4RjZNRLpbDTD
M2OF8A9KGC3TDEB34fdPH/IlkLreFHfyq4Z5tc35wZCStNp8A+1cCGIn86svQtJQdlS34xODdEzr
mUrI/1gwNuO/eWyvpK3SZFRoTT3i9hZgDFel7QpCQsLm9mFj+xefIsyO1Pllvao6I31e3UJ8Ozj/
RNLy/LiZYqE9m3eTQ4tX5Kfej4nkFk1Os7ZmSbWYgEQGkJbJO7CwAVI0PLKIbzXMJNmqio5oQIdP
xF59W/nopGSk22/XTz49LXsTPJKrSIFIZIxwPXcsI3O+j4OcnP58sOqIbkc0vTsnS3AQjPa9iEpO
mUnPP8DXkq60DBaNOKgDmjhXxt2/gsHA7f6JgoMda8CS0S3tL92idzexG63lsdsMwxaWJnpcxtVD
rzUnU8PeMCdAyXJulHDVDOhvdQ63cZDe/a2gtwHP4OZaw0WKkwFRnVGsRkO1wchVN+IHVRFpYHKd
toAvCEE3iVjeCjnByCIUz3dYebvgPXFUsO+jA+V6l5p0bMRPAW2A/371EaCd2h3D7e6k0xW1CLTL
kSr/FHmCY0HV2bzTcq9IkugqPql5ZG7Swi6zO9ZyMysI5l9sk8HaBFAV+J9JVHH7Ul+PA1LfgW/O
G7xRWfJaNNPnjj7/xNxj9QuRF0QNX1XCQIgPEUZuU9VQnvvbl2jXZe5vtUafTiy4JAwW6A/1UYnF
2mjhS3Y5/sihQWS6CG0TAKKcft2OMwFkFQK6GWekyKUMF/kkLT3FkCfO/QcVLQdu3J3mFwQ59Jrf
rzouAeoM7U6UJrTgDYgNWxGMoGW8xTtCxiKbohxG4S1W9PAPkUfhoany6ItKzWWDBF2AW1bmA1dK
5vlM6b+T1j9J98WhKwdK3t5CIuWVrC6FVy2+m9mYaajGE6y2iMWuLzwA8soF4LCKM8D5zO7iK8rz
O+zc5XRBsJ55pMbmEtx2+wq8jD2Zdfx+2haE9LzJ5YpyMZWr2hTMGCU97N/B623jfFKEQqc7kDKA
NYi+8Oqe7yPibW1mm20vLCWfRz6drlmj0FR/1093EIDFMAaTk+ZNWBAmdZvT9jDhJIVAigFtKwoj
7vLI+nmVvrlPjJI3ICuLruGbvWHmXZ2SDEmoTZhHx11gmmweiiaGkzQVube+0ftcuD3KRVdxjgG8
rO9pCS6kf5UzfakwLJ/Uuv9/YPb1Ha5yk10zQA32zJnDBDhfhOHwOKj+fY/HEKCtHaDdmJqoZxQA
Q+pCGXKOf4sZALG8ybKrUrUPa8gz59dYVrK170hwUdLZiERZZRpvUKNgTGZAVMZ77NrwagV0W1DM
flKkpzRhmDmqHqvCHGYLdi0o0SYbgkKGQGp3ksqkBTE9/uMX3lEkGYbfcn8Vh+2JvVR6snBnvXLT
qCtUZ0lahS7p3L/hTXSzMGJRKBKY5NzlFgwqLcOl/rVhM+nSxroJxAEsmH4OyI5lCOEo/zhRUxCP
ErLg0t2S5gft0kU1Vn5SKGsyqcxj5l5qdSdYFcHFj109J8jtlfoLHLqgRcVcYGInzXps5Y4tCK0R
/eIZcmPut2esQjuNx7wgoZMsKrYYudS9UKQKog0VfxP2ECDNGgc97p3jMuhY/1+pQAQuQR06sQL9
PKTeSzIw7RnOrkMSlhHSav9r0mwClrkYXwUIz7o56NsDJx4G5Ww/Ityp+cSWvRGWMPVSD9o+u11M
ACBqGniM+AX5F4AxIrpt8lrAM+ddxQ81iOkzc/xSDM0jfSt3/b4z4qsErx7uulpd/s8jbi6XNSk5
rjEBXNHtLYi5Rf+L1hh3irgq/s9EVrI72qQANBaVpcfXuS7aIO4BxWTcDaRQlNKXbKFPT836tQKW
ltPm2dgyMP2fP++WWcqcqGBgXdew95MbcGYk1AoM/uGTEI35nX3fAHz9Z0ZsFdveX+L4GHTkLoqa
uex4BPr0+b+1oOvWKORIcUen5Mpih2xKuaGqCsbhsOfkvNOLvGieO83+pX4ECTEWY+DIHE55qu7w
zERlmhOWogFdUUfrE6yHPS+J0DU2cgxwmX7qjPiXgOtvzSh/rHC2tX2ucL6pVOnDWrr8kvhPFilR
OAxQAUcyIYRYherwIWrvZB6fLRynS/nEFfg3zqpXqE2vg+Q2hPaA3bqfxC6LhekEt77ENpE1MV/d
vV/uATzCcWu5nHOfmGMOVU2bbqbmcH4XSN9vodY/RKa5t2Ncmnuq1PaXmm26HYs0v0yGZQb8mTdF
oZmgSCPB9mqAXWdGc43VlI8YB1r1ISlwqZ1vCvwy4awvS9xy9qXmzHrZWxbAjuscGrNcvYP7tb2i
TZEPPKjYFbNO3q9W5EcFbiUPe8FVHqGqvxLooqmR6RyEJnIEu3+rDTJGfsRhCT865NnQMDCh9IXV
7J1FmviC+Z+AaU6YG9xrupAABgfaOmm8OCKSFHcQ2D3ppji+sfhTwwUBiQkezaQe3mvt4290j3a8
Q4S2tXSy4zTHSSxWUF1jGIuGAjYp39eYppy+1Kp9feqcqmeEQ8sxqUzK3dLEnKMhVwSMMgg5aMyJ
FUW5euw/yRqUvFVncWscWdNHBGXMZDmcg73Dh90m033GNMgYbcdv2pXkYJfeWx0OVl/UPAny+uhB
fRagJaEI9230j2hqmWxdiCQDs2v5NJ7V8hGXrTMz7nYCmcg4SMsadsbvzjF+2M9M6bxVFAt8gqlQ
4e10j62BrMYCYXKRUD4cjSYkW5yii/rHMfovNqqFcAWn+Lw7GIg/JgAD+tEtIN2SCDRuhxgeeUWX
EcuNhn3jWsIS2dlss6oLzW8Ep60U+1VpZG6wGIVLPd/rv6OVptuREpi0bcP2OhLlDTj9n9asNevA
SggeZVBFne4Y2SFM2/naoI/90mc/7xF7FdikJNqVX3QpjqdHcZb7p5Ck5A6jTZivJsYIsirc6iJG
zBygIxl0Mvh0Ic9Diis5sfFHkyMvdXigqzXPWDBvsq/LQV9raNCx1X772O9pODadYag1GlZh9uAW
wIks6ls+GSpiHasRrRaoPQpjuMw40/xpMfbWEli2LZuzSQ87chgJzWrhlnFnHsXpyFuromlkc7CM
RmxmXDJR90uegPJ7yFXD0rP4zZXa8Kx8M07GJSVMwniLhogFPfhi5CcXe4WpkkC7MEP0SIXfe7DU
ruptcYc1G9JIz2CymIHDnGJ2JzD8DdG5gODNCwEIL/A5XUmkYdLQM77D7Td+2AzVmdJueRGaHWEn
bqlmPaWkLDEz5pnRIv3ozB/Uk0CoTxMiMj37qeKau4V9THMV7KmXHq7VLCZ8ryCzDdVZM1AzNbbM
dKNsQWxeMrXxqcndH8ZDSR/YOy8iK8TcmpAhRKGY6HqETdb5i5M0f8+2NM/OESQkCYpRW3/atZDo
jDd9z/Hj9mIdswb0FAFsHLF27/JEbX+lEv+rQ58Ca6+H9VqNiK0TrLW/sEg+HZA6QiieBEEu03Bv
AHFm4pIQ//WP+UGNW6SGe3MQbm0AXlQE9yRdfBmMaWzkvOaM5n3FhdjPCM8GmictJe7PSPDueULa
pBWK4u16zhel6Tqa4Rgw6N/zD2ZgoiA14gICwiaE5cXBnkPevnmYU+fBa0ncD4PFfdDAPrYoqhJg
iTum0LKmg8Qf4GbWFYLkW+1JutRs2NtnAWGLbB7ykfqYBxgv08LP1aQxUcnJhCfI3SxZWE48048A
IV2D3wT5YCscC2LKk/s5+NGpvjPPqGagXIoqiClHsvxb/bRMgcVppzN3RrXk3wLpN3XeeSnQyCe1
G61wSalL7fYNsrMMq3WcwXH0Q7BlC5PYHvRgRzfXxUPOYhUFH3lajycvzeD1hRRs0U+xJ346TkOp
l9L/mns/kOevHXuLjrZoIWobqY/Tq9ZDN8EnASOGl7TMGh+jTSbhLvXjMF6rWLydWOWNHNwPMPfp
Aw7svLnp3L/07QTc7BOSwGi+pAN5L8LcAsg+t6qsc1vjPGcl3G6yt4nxP2Xpb8qnLTytj+yDbmXV
wEqYgW0CPLil9e9SF73T7Ik2QukJnfaEe+JJyGcqymIK9sikPNThrOUEEHZLc/STNvnx6Jr6u9Q3
t1pQ4rJCBGjfVwzDD0lkVWgjfHxv8nbILxM70fKPHeoGiYoS63F8A7OxrkOcvNFv2MLRaTlrUnew
HnfxMo3l+4tg1r4pZ+QZsWCJbeUeUOI0RUBmHHYNGp5B63fhHrORdtyql91/xQhg/OclpCignyyA
eYM1zFw8rNNrgdTRlQjaho9DmzkHuMRCTrlekzwaKCXMIUtR8URTsowSy/hbn3tuyfEjiq8dRrm/
5BAQQakmr5IPVIKv9LhtW2D16PxfvUlYuCIozSxVUGBG2XhFg0mM9hMXxaam2xU2ZdvEp50nqBhx
41g44ZNibaYm1V44bEUdyDtyEpdiSgH4qPyNe9ejayz72Bv4zRCJvedEn38IPK7gHvBrKUo02zkw
lDOYBr2ESKpxO+IFWmR6G+OXxMI6+yUS9d7TfLObT5VWy9sygdEfxoJtsKECHwgeGyFIckzy7SDb
IurkcnnAjYXRtLHFpQzf6pK8XidKfL8Ld7MdDv+N11/5DZtGtlHoBLjjjm+n6sO/S4XH/KBQEvcl
qc1DMSG84epUbmlVcFO9/xaX9UsowHv/kIs159XC0S5Wc+5fX3d4SIHDybkEz9jy0J5LD2/E/H/P
XZ71qZ6/nrKBKpBROVQJVvrAQmQsS2bHT9rrp3+mD9zMXKnae9FNDylfcqR5hrYcD7/NrK9Muomy
yvqGBWS0+FHZ/zp8iUfVQKzxieFEsZdi5RyaLo5aaPeKFsgnSJyvFWYDCBVdse/NrnRJV/EsEQ+C
FF8hXXmDK9VMZpJiy9+spf6C5Sxf5e51a7lCte3WmbQpLHH/A6QNxMNUGKoDfg5m6VoErnl8Wamd
ylr98JZpzHkfA9HEWRBcoT1LuNV+Vt8sbC8uYB5ZnH5PYKFl9Vr1zYIK3XPCrulIQ+s2tLH2dond
XCfxCnqrJ6khjM0bz+nDeNxyzALUASNbPQEe/50amdWYX4UjqpmWzglK/FqwijFDVwP0bMSY6q+8
sWLp1NDTT4N5cYNK7qEGGJ2qMk5ihyDpzNIq14TzBmm2rX4mI77sIodipAJNb4y7Q4oyfNenPbFI
E6Y/ADeCmRd5S4kvOCA55k/kCezOun0gTIok6mDPtvFYZhldcpDgbcMaO97NHf8jBUuZb1Wxbshs
AkPQ1m4gh8UuXUdM9dVfni4UJkDUpR8joducSYGrxIecuw5c5JxZWF7rK6cJmF7B30aI87yXFQ1O
Q220njVOEN6vSAUkkWAr5d8xRF5xTHIGOzU765yzfTcCMvArCwn1iHf8ZTLzoR2eJyCaeA3U0fHS
9AtIp2rHvctBgl20T+KrPac1yYG/yiplGhbTdaA7hkQTDtTU6+ilosCW44FHncCZP2DoBlTkAjHf
AgWmepZfywwsYPvtbyl9Y+kLdAu7LkvR+t8vU1B/rZUc0ClchE4TUDQ8FuURoQBq9RFGV9Q7CpA+
bw+4UD6wx2jB+b0QZGq3UdJaCOZogZ22GziQubuqoCL/KR/EineqxNqxi4V4CzTv0wdcDVfTdJRV
O/ZeynLKjlS2qbQ7OSDSbClUbUtKRWDE+1GvVWOlQGehVV9e4fDjcxlUt/Pfs/Rgn7u0jryIIiXp
zfymtg/Inm2ut2HJgP9wdgWQ310rGuLPN/cS62VZ3BymCswBg7Z5iWtbHrGOqfH+13mGXlVxykW1
RX4eUE8XQDYzuDMNJbbhchKSV7MQSoiQQ4XBZM7DSQ+kSu/DCyeXiGT2oUIoullh9WAdrWHEPsP4
yS/slQIRLd2uqqD1jeIjZF40PkLYXq9P1gJ0fM7l2+DnO8dhiauhBoDcPACdufsTSccR4S9CT/bn
bih9zj8uSZIvsEmHvngajHGn43w0IasoByuM8I0lpk2UITCZtxdnwSNTsfC6wfGTEwf6HZnuvg/U
8JK1oDWTdSejVzSJvFdAnwQBWm36FcJoWh2M50GCAcyjCH2vtTIzYjHkzbWXmdsd5TvF07C3oF/5
nMLzJ1XQwMXjU6y0SAkimF2XImQ0TJR1BjJpinoD0E8h35KkYdQ741gZSkBPVVME3kdwwLrGX1Lf
Y4gnmLZN2IEkkpgHbqiUu7GC03xKNCxlSL+U82/h0eu+vYVti3TQA5SMFsKp14zClFgSp6NOXilP
o0N2KcESNZRpkec5p0s31CnE6XfoBym/DGY2/nI3sRfdmNH3u077dl+howWooieH4qgZzsnHQE5v
aUugBBlbAoIYOXZKUguxKto2meWZDJhEZ4LTi8t2keKSHep7bIXZBpqfRyxqDSVXQoilM5ZDCHRt
cOq3e93hK2oXT37PqDPBugrSeXqCwQKF7TEflPyujCSOdaKIA4R5IlDXW58K6u5ZnAR4VMexAQVV
4QpunS3PfsGbTDOLN1AxSFcvH/TEoQnqfKRW/9KwymNkJoo2A4MgYemsVhUA7KZ+r3+MmyPCr9iP
+7Y9941hm5WuB7gK5I+4WC2oRcAWHYeLBRmKa6YBdx6IVI0ydmxDv0R6K0orAUZzu/1aY3MkhWdd
2tq9FJdzvQBxwdRJhVXseQTssxCk4+1K6prwZyhHLAKdwomL5h5NHFrWrRkh+zy2Q/uHb3G82W47
GU6oZjTPmUE8OF1v0eWWNK5JBZ+bRdNpp0ElHRM+TtnZhN5d6lINlF9M/IubXrT8D9Q1wKQQ1TXm
H+d1/D8ydG5hxYUAnHz1Q0frY3Nhwavy08A/vuFPwSyHSHAlUjr3EY3q112nSCLmGi3gxxSED4Mf
yKadoAn+WnX6/UZlmjs1cblp9JwOfpCWnNbmVv2Ic6GtEzRGBA68rzYYWDmLjQTdTX4va4h+W+lH
nUbXb61hR8/HVjKmgynZShILxqM1PsKjzqGW7FliXGuYL39BGS3jFnAsyMwYSvYM7d/TMhAlV9uQ
0e+6dTPVt3T1382b3V0oNqewN8rPsjUVzAW6cFhj67ZANGToMqNIqGEwrVG8GcvhlMgGAyKgLYT5
vVVkuk5EwsxUnBNzXCBEMiC+V3Dx9oN7P55t5sni1elru4Yoi4T8Jrr8P9QQpLjXUi+0L+x7sQEW
TeBCODN1SN/kzPA1hp226wyhor/GKcUWxfpInJAr1HJviJhHEpYsbS3b/UQbRf7WMaklGLsLcria
b8UAvf2MRQkRTPkeS0Or+PkqYOXJ2kFc2A+TKL8zgVwNRijdcKMNNSNGzpDtA85x2dQS1XoiiJ7b
wbrMy9UpvOSc75KULU2pcT9JnHOMFF6rCR8UXVhRya8Wd/XE+bUMwprxWgP6CaDsf9JImKR+SBqe
JeCLgcS0qjP9+llPXt3+mj8qZds8gHd2kuxdh1CsKJedPdcCZofweMwMssN0U0SeCCF3ANRtLYjj
Ov15wK2OJD2NiePpmXHANRwCocl47G4DjJcmi9jLgL20eyB2r3OZ+A75+Npv8jl0KLhdxYTc71hq
MuXLpSuFC0cjVtT0RTYAmbcGEWV0YU/SNOyKFqY4RN6xqZyDG2UAbKvWw9WzszY21M4W/6HBWFho
iqLKaeah+LaiXbUm2+PGAzb5vLxwGOY69yWeXOf1Vlk/Lntxwn6HPWmb8EDvP1Fr0VIh1L6jDaCM
+B5nucRYB9mrBdFVBccc3g+pPKpmkI2lHWGxQLGsUIheV/14UnM0c7KrXZn7GhqblOfTViA4nRfJ
UTDNGcDVNtVrscZULtvDvsYWuoZ4Ih5q4tA2Zfi4qJgpeoh9CJtjHv/hTvsiBmeWZiuwYbYjgkaV
ipIE7K3BS68MxBHMmvatQU4jvEf3i+QsgxuaZAtiK3D5nWRsVCjZv2w4SfWAG8xbdtaj8PdbkvNG
l92iKOjRCWa84J8eNZSrhYsVkOR257De0WzuXCPr6WKX+T5Mh8e0qr5e9QHiQW0tlSEQkAbI0yz2
zsVOTX1x6ii3R6Q2Nkj+7iSd/dk55w65lw0bDLExxI0mHZxK5nInrJCQeW5f4nZA4aralhTKgBlK
rPFTxwRaYJ45UpA7zxtWALeRlEHujVQk7cA8ESmCeoUcIMoAHgybx3E5jadeQ0J160CnWc8uFOcY
gQnjNXF5wm/V4q7Z9xAofDxm3lz2/g2ZygSnWwA8asxdpy9+udcnO81Kl3gX79Jd9ogZjVVKp59l
6fgnjWlknuzqjrXAlIrnoMziFiPqtaA1ucVEoM+aX7n5qbUTEY9X1m3Fg0CSVYsnuQ36Cpx/6Y+Y
Eh4EoZMRvEovHBbl9YrhsE7UpNJvFzxXfnrr3V00vHGem9Zpyv87A7wuUJ2CCMLkmRqQwqb6c2xb
rIuY08KwtqtGKSS0Aoc7K5hJAPJyH8xTdIXVfkKAsfR54qHlwiKUGUKCOPHVedtVpfuIUgEvwj3B
IFlig42ys6FrLPqpS0Yoq72tM/Ti+ailHXfFC1GL72B90364SS10rdW3GPJMOVN7RnkR9MQQ0KNd
SS+btBDxzz4aZ7CmYGdWizGUfUUfIo1wSz8hY/EBfWh100UfQ2yxxDu4bK7llcbhyxUehc9dyLT3
INvb6/ifBEQuk7L4U2ZzO54JaHpNrCZg9tmU/aQ8FSss7q+GNaWDX53s0qpTtQoX4aqy8qBxeqac
o+53jfYM5pFRT7sVQr34VdI5/9tul4irjWofhvxBSbrnJcASmEty09aEcNwYhqQ1NFFC5Kqmo2lX
4dcho2v3u/EbxBIYnsyKWVePD/YExuORzeCXMHzdaDQegOCURDYut/7uWhdEyG7uoMtNJ1Qy/D+1
ulDBqFkHuht0Uw+8GTB7jPzVdUqtyXlbBKsXRszIcv5ttZMJuYBIwc7TgpQP0B9zEAiLJvWfZwdW
dqr73Hh1GzQv6VrwG7PaaSlDM0vsshlbH/m4LGi77V2t/V3UlgNACKsMH4nOEdGBSc33WvZeVlVx
2VIJi45BQ5TVgHn0ZmMrrLxpnJGDyWG8Um2EU9PEnhp4vKgq3oig3Q7Y1qW+8Clv9eSHGzgyFhcw
46pjz3t4mTJTVEO2wnaxUY+0M6JWDXW0M8jgzvOiV85ILd8kRJMlTNoqBw9DAjhB7Ou4mzFXRNnI
/mL0RMMj4R7RqPGd+c+rggobvkLKVzZHp/TmXNesxy3RopuDIcYxJNZvgh3K2oiTf956Yvn5hCW4
JIR11KIGaPExpH/PNPnMWsd2mOaa9Xy6BKp7xIcixgyJEDpBFj9e8N5ZU0sD3WrM4QePkGHoo5pW
BtlMGv/Lo6ZTYdTuHuWRXd+Os4gZRYKghj+G7l9ys0AIPfMfy1LhAe7gSfVnYfqKKY4RYt7VkeDN
/SnZZm5n8c5YVt2bWmLhvQ5Fo5O8lqZka/fFLeSlaMt+RC12crwkjgdtrzrHrB7Ck1mwONNFXP1R
GmRM6NO6S9DwQZvlGb6KHfKSTehgWnc0WFTO4RIZEV9vl/3p1AgevMcwD0GsQoYz5GMFMbvO3O78
clK1FbZw+9hddBJ3ZkDr3DBK8BO3hFzEgnPwg47lHLtOnpXVHpj3z6heOtRj2AXjISQNGrKeFVmp
1LTgmmsa0kF9cITQl1OEuAwJ5y83dpIdO0u051hLJlDh4FCOTZhc9krwl92YrOLri3I1x+8pf4aW
OfaLiS/7QF97sHqYyMyBL9ZGfeHAprSFGOazGWaOt4VT6C2+sacHGVl2KzCNP6PX+Jy0JbpxsSvO
OqZF7IMRMOp+o0xC38N/oULKVTU5afIxTkSIQ2XRyh3rgroCDie76oI1GVJaicQX15eSxY5WMcq8
HMRtZ3VltGgiMNmNxRBZM3zsRDMWFns7zl23PJlCnHz4YCUgxRZFZw1eKiUndHfLoci5GwDTBSyF
IbdeBoeffXq9arroQ6KXWZxZtDinO4GdnIDpJ6Uj7nfI/uDGS2RQguXekBCqu+nuF1sPnxIZEfLj
DfUyfy5uAl8ukhX5arzbSq3Mggg1kFSb0GDDAfvCGwiZFMiM0p163151AudThKcbzdtrr7+Fo5wm
tw2yroh5TcH+23QavtaU7j8O0PtvvwRGgnSwcppcu9RQLuIVBoD/+9BsSOuVr1gaDvrlaWyVHvFi
rSJpumYPQqQNl01HIEa4ojXJt1J7hWJ9lVSR9UJqUH9aTLlsy3vH0b21Xe8pvQJWUC9YKsItH+mj
7Sn0RDK29q4f4uykHC8U6SDprWHckyzF3UVlA5mmmz7Ol08gy7nMIP67x56XZMIWbA+RodCF2j/W
w3TX3BzZRZFgVzttv6WfgOqEHMu184XCKcoCHAMCGYSAvqRoVnATbeSd3PPruDPKQImrsBOG8M3A
Ls1OznvrUKuEHcd9l7z5yMhW0SPY03bfD0YdBo2OhzJPdoxK1o5eoLbZBJIWc7vrvsdNA2H/PLot
J37mxVsdX8VjhOenZPM9esZrfUPLpV0+xGt/Ta4dufd9JTultVwBdEcN9J7bdjHHt9KZium+HGiR
GZ6xvt/BYe/nLdLF/G6dv+h5TK1TxURBIgrT9ljF3Ojn+nZUt709A6kYPL5sPJh29+pMWgWj8zvv
3+xUOO40YVCbF5R8yg4TH6YQTPBMW+3KdCDKbfzn9A/y6g13kUMyI+Tq0GUDWziY8F73L+3P2Lqq
KXDQ9Y3o1p1vYiZP9QSGgt78KgYWBL0dWVWlZxEaUGxveG2/+KxQMYiMioMN8ikRE/N8sgAu8qaX
Zrbrw+01Bn83henTz8YV6Iy+/qeNlct+tSH0ILfrpCtH+vxCJQJVITdrok133VX/KYFLg34XflKt
CcI3dGW1YWUF6kvzD7GsY0T1EwJeBheb0IAvBBuvjEqr0j31dNgVJ2kvR9fEIxMfntQtTpAfsVRa
OAjQloIcsSkzz5OO5IJTtg0Lgovu58/LeCswc6aWseKCGTArL9QsuJ5Xm9zumhvbZXXQH11gzebA
be7JsuHvwcLkmJGL8Mv1Ddrfmi2j93+TPB9V3AWW7B8VZUabAuLGNSsXOKj2E4rl94/tGxxGnFZ2
hldVAhwKU+PxFcjyworVBFDpyxDxpbCxvWm9FT5Ubv6uZ738BG5mbaI7JVB8S1ATqaEAxMiExnMz
PKiJc4wLWPCZm0ExKePTf9FIXqjM3tS2Hmrm+7lQgh4gJcB67wIJHXltKgXpsHPacAbPTRyWz+7J
4A0wPytOqK1iFnGBRN1YnQpXW0h6ZdCzEpMFHEKKlpvTq2rZpenDnwLw8+SInD8iiNGhSKEJ1czg
csUAKXF0gUIHYj8UTXRF4ZF2rs1grnC3PHNS1CR2JbyhOaAt67BSNHH7ZBPL0VSV5pUaYarujmJJ
xzxr3fZe/ULmXpy9Peu4N77mxiFZE0E1Fpf9/Z8ljBcJ0hczWuPgFNdnfMjCr8xcE9UKXk9fZ53k
3GFVHim8daVcXnE5Ap1kS3Tzvn7+rVrJzWtEwHZbBb6L6150dUAX9Zsm1+K+d3g4rwgGCHeznTXV
VLfZ2ZaD6cnumAeQQxogFyHyYqB8bQ7BHA0kUd3Mo6WBDy1j/wpgmk0JbYOQZ5cyP5p4OAxudKNv
jj1cOzCgL8ZsFZjBQD8G+hsljAS/i36E08znU18ABSw6pHzpwyCPFItWHUxiG274xz8XkIfsDE1S
qDL6RlHoNAbKe0HOQRrYLOyQvw6JYZrOuiXTZtSa6YX6qDDJJ7kAQEwU4IxnpXsfphChO2RJLQkL
uiEF0PofiG5xSSM8eEmeUT9RlByjX6XiKDzPWe4nDbP3Tozjr0dJkBglzb3h0HRQOz1KBiXRFZDX
podzxgnqhu9PWobXeygQ3XF0FgP9p16z9uceYVmghGb1tLUeeIAM4p+qE2aG70MisGAU+nyqwxaX
z/+FverPQMrFWAwdEIVOPsaojUYXMDrkYo/jWt3eTaVQO0BhOyMfu2GrKvcXVHxM1VOJ6OvJx54p
mqtlx2bVdbI63+dcdyBHgE8qvvCgS8Zrjnm5FfD+BkLNuEnkO1Max+T43ZGTGRAs8MIRhLbn9A4y
5iZqAD7jL5a4PKEn0JHPyaZDRY6VaAjgqZyp2dpI1Kv6cSSIvfMpOBSv4G8/kgrM7jGMGOKZQMDU
ngQQv0y18AXTA1Wxv9aUxkNsstY3yQ21eFlU/3IbKwnWns+AKJsKxSUpSDDynIlodPB3dGkO7SbD
hA6xIJVBGC++1AQcNrEH4v6KsHQslmNr35kma7s3h/7rf1rGods0mfCBg+vTnWTGSOkJS9OHMvWL
K0AaLohuCbGOiSyH2+IQBAobu96+6Bq1DC7Q+hMoMw37nnWiz/TKptUpxKcPbtK/G8V7QnR0JI7u
2IFgkiV7ARcK43gIGKBkUTjlMlttGJC/UujuxlZx9f+tDOoxSoaaDzYaM6QqTssNY1BjAHBxyCwi
u426s3S22L2sU2GnzVT+mu+covNpxtqQG9UR6kcVxtscPjFHpUnQ01+Yz8k4nWo7WQ4pidNpx97l
WbUpmyE+zvIR1v1uzzownanz+DdXIsIw1ayq1D8aXM9VxXOK3QAmOi1uKajjIoelo23UAtkYBWfV
YC1VwkymwGMRR2ctGFFgoLu+7LjncE/7fyFzFhsdvFU8fdTrdMS2RO/pyILLg6bUxYKw6djhts+9
TphzMwzdv9AyQWrPo3DV8kBlWu+twIM1Fu6XBXYkGps3HQzrKZRJadn3ni5XDU3eeYBUC5kwvCiz
zUzHbY4IK5HUJzfM9C7CQrnxdkw1SfaSnLNzatVi63bZXlhEszqzVJ8Bxver7Bjgn0el1HGZ0TME
EpmVHoVeMeb9h9yBfgMEYHzX0+WbhnIZk45AvW3DQqVqhH8OFc0L97mkrb4k45BUIgmiCQcSSRqV
4LRBqrqzm84cFfk6TA7xCfNr59uKz7hAQNEUYhLI3aEXvkY2CsJEwV7Nv1fuPMV7nug5wvLZNyGc
s6iDqsMfuohKTF5vUqEsS1eD8MEOkA56D9Q0JevUQi9/t3+hj5yCv0CzBS1SI5rDUjsTq9HGpS+E
YH006QwpOqcv8p8pAFzvfiGiDpPWYGBFNbzF0V+EgW2XgJYbyuke1RFw571zr7tc/BmtiG2xkAsg
rsA1r+V6a0ked1NEyc4BLDnPT9BgJqLT0NfUAs+bl1T2KfR+D1cq5hf4Jt+HH6Ce19N38j5dMLKZ
S0Caw8y8+Fgm4wngXAIzO8ETYjWyD0Oc1lS9SnLol4I6OmaaN+af4ndgNuUMaRqH/FekhlvG3I0q
NR3L7n32hVeVdN7Y/xSho0MQ0bxwIYpYwtts0L3CnztDpfP2LjLtgoGaBo+pEOOC00MUHMlT7t8m
JgN8fSfk2RKv0+8mCj/Bfdmk0BhIiPMS0+EVvJel5mJaPIh2OnY+nBITJW0B78NgTLcBOj94+CVK
adK0lI/SESVjIkHs3diT3648n7A0gtsFHHyMdFajDovj11kvY87HDVAUy15qkjQYkcJLM2sNy33m
pbe32YiMJnEpNzYilncucpb550tkAYOMalOTrJGYGFhfNBtXoEZQ89C1u/GKzvWXI6l4OYS7Dfg8
s+paTNvaiTYmahgMIt9HriJN2qexXBmPQEMOBGLV8f+VF//SY57hEq2hSpfWpABxAQQfFNKrXIEV
Uvu6RucoUaVMu9vb1TbtxQE4b6Pftuprao4HfSNO3/rv4LQBfH6f/4e4orTzWeG895mrp16plSqu
RSO0QB6H3deS/r5fgYqT7e/q38a29dMTe+5QyrMp7QWic4cHZrMvQiTEFTfs2sBiq4E2r7OufO3N
ifHVA3pybDcU83cPT6cp6TWlMKVP4GNZYTIN0LOS2kLODvOli1Hc/uNsMkCY8DSqwCowopKDhpUg
mkKgdZw1wHmPDC8rU4NHhue7y89ls+yMPkACNAOcZ7nsqR/phhpzhnjeOdlYhzyjKuyYkWbtGU37
IylRrYls7of4cGL3J2kK4c30lPix9kELO2IkM2hROb74i7K/yykofsYI3Zh1oC+2eMzrMgcFpUMf
+5mf46kf11VlyZI1K/tCq2VXedUo29sF1FDtiGIBMf41NK+NMScDwvSUKWMAK0jcIk7BS469VFeI
2SSjJaN/giQOP0XB9yVJwZ06r5ZakX2U4r2Tu6Yo/DCDAMXunugkE9tyraY6cmP71UJpgkS5zwpP
/+YPHUY1Q5PR+45S5OPHMktnFHJduTk13u99Z28Tc73KQFZ/NE4bI6c0Xtg8J+T3o15a3M1HN8AV
KIRytjdFYeoB96/NVxen+TeMldWA/kLzcAd7ItKTyhEWsuCV3fYObZTjUy6gkJdQLunEbjrpRLUn
FSszkPY8bVqrxp1syIkPI9O8Bc0TN1rSZ/YTl2fiRNNQHAO5JRzIFMAe0dVHohfR2kf0f1e2ovIl
w7Qh2FUxgOi2V924sHYOYa8CYeIt7/PY6m5pO4nbfkaM7uhvFanp1OFq4Zj3YKKmEdYEvpYVHzL4
+84NiWqW9a5otBbFoPJWHSswNq1Ovcfq3Dj65QsV5YqX2YxtFLJN9kSqeRRIZ+3PCorcQE9e8gQL
hhBrYV5puNsxLKYy4253V+U9b7uqr/AIQnaxE9GKIOu5wOPz5xjwgk89//vMlCVjflRwAOj6ABT7
XM+XPS6hOsey0RWRoeAl4W9JtX2iMVopKJs9WYs44VYPgocJqrYGZDMfhP8vn4re/+4mxdl0dFpw
wO9sHDBtbDhdXLFQY8GB+9JgbgtVsPTeR9uiCK56aUiif+8Prs3K9uVkvdnS1Ngm5Yd9ZTX9iE5A
HRWDv7rWjkBlD8Fk77ygQFVb/SddgPzhVLqkKo9YzmKljc+iwb9HR+z8hBR9d/hVlchnPutlNi2q
+Jl7kmBKCU3CZkoT2BO7QORsf/623oCgKNm4uOfUo76MjiX1mWTWH8qPHAC2VVErpUYEwJsoPoN+
6K+U7Sl01wXkXm77CebCxnr6kAuVONyO7/UT0UBtTaGgvu6XBR13ES3o69DHBVFupBqcACJ9nQfC
83f6XdFTefKNpImfKYgZAQ7gPWd5rWvhvM982Gyftm6agq9oPBDrClavwkBJIBUR1H39gOgIoDjF
FrMh/j+5d+AhrrDypR4ALTjWSCUU3Xm1sDIAEY1edIh4cmPvvX/IcZA6toA19lpGiX9JqBOEBzsC
7tvN1F0ciPNf/0bLjaMAjKV/TJ+oVrcfs8+uNEFN3oqc82s5YwSOCR3oqo8/okOiFL3MJRkpcPI2
7M8vgNYXlYdIzZdtoxMYO+6O0qkmueI1IxlSHQqjVjvjC7MfFQ6EfDxoYk8V2ylCm0t7jpHcnZSH
7zjvJEV+TkYhMjf78WQ5VE1YhIDlmniNXWNI/cpWMJThcfCXXytDzuQhwoPlxEuigdqpkeCPndy5
K/W+TFFUbC5x9cH8oyjsXMf78w3WfPYPXRNwBEwCCxShXoJ20lKe/sfjXRhV+xU7vZDkexWFn4ia
1NMm1sW02pXr+H7zILyVa1bCP/0Rdg4eC6jdU4qU7K+keoV/pPMWYx4VUtgUFXpJSVeQIkwD0Lv6
fQq7IzlMIANKuy3TA2XNqRWB5Xi+21KGAVSn39gfM7SwBZL9UyN+4vNlWlBMAdkb3ogDE8kv0wz/
GKT/zerXSLAS+vRUhV8qAsBwYlmUImw5vaQIiWbbDLRcL6gxCLvt2EaDELKsXoVFU4y15xHK6SIw
MYXpR/ZHvEGWnZei8XCRLZhvlS43ZfrZmiFcTGyeDPfZccsh/8pZYH4V7YA+UdHfTPZknnR4JeZ+
okfsDCEJE82OeL46uGu670GO49gnD9PwmzV0kz3jClpr78FFCI+B+ElL0EjeiTMa2CuzMXbEyGGS
JRyuvJu6fCcsgVViurRCObE3C4LTgtz7rYwYTZDmJr6gxnncx4d1RoPY3VGH3YZnU7pnOAXILsCz
m/EwBNaeGhpc44euOWGXgHrF7qVBNArkqDrK66Nghvr+wRx/Q/mqEGZWre/zQSVl3fLrRBiPcqfg
tC9taFox5ycqVn60oOWQ52g873IF1B0Alrx34F1XW6exNJMBTxB8F9yrU3+DbQ15vDSgwQfyq1pN
RiLYp7KzcI4KrGsk72MDaxFRQRVU5ZGK4lu9ENKq643FM+NG7U0CYoaZnhVpCOQZs4rR7ZtG+S/u
t8Yso+FQtSJ4vsZfWbPOGuTN/mb9fNb2rh5CxhamyhjC0wwVbocWv7Y79B6WOEC6o9D6T+gOGP4u
HTm2050MNoMQQtd0v9pRERZ4NSYj59Kbn7wjPacGh7WlkE76HR3lX6WU5pSzNKa3O2hJ34fmWw+J
Xzh7+Tqs2R+0bM+xfsOfzcoh1+dBHbEQ8VBct1F0gqXmsXJ1I8sAZ+Is88bZVNL/WCU4PBpaF8Z9
zHi9P6mBvPJOrs3QDmu+2eRvVTZh6iioGSwMlhhJiTnh2Tv8aA4frotUE3seMZYkWuVMzqADmHVJ
kCnD5I7NHfpKrCUh6TLBXqBW+MMI0MJbTOQg1eRqs8fLCcBoPVIo6tuiNlCAQ5tVn+AXrXFz1wM2
1QrLJ0R2Ooq7s1COgF/YZBTfuho+zkrKMYEg1+/TrKrXlZ2s5hVzFDVb2RmJybKwrYCVqw31yZR+
XeGrrAVWScVfnVQ6EBS6wGkJ3/WepEbzT0HTdek9Ht8gOjfVC0Lra6AyvHlHwbQTXBLL4T9oo+Sg
Blwd+TJPfbXbRaKvVFFhmmkEIG0vCh2A4ELHhJy2xQNQiuo7wFx7oynrBdkWvKhH+IuEKpwGIPRr
KNDzNOhjK6Qbf+gSPX9bzi1F3DczWBvYbhZ1N3EOmy69dt4XLa+R+0ejZKzVPyoae+z5DJefICE6
pOeW+TjBYo/hgp3eSnXVKfjW+HqjkMVG79GsbPQxXAbpHZlvNXmfHp2xIwqf+/RTgllDebVswWhT
OgdC1oO6t1PQ5ttoJ2ijVyxHGo04/MZZF/7MnxFXUbxqyofma4kNKZWVRpZY+HohYa/mKldM3xKy
3McPdPdd9vN5y5GWyZXkWRTssDIeD9Hi5N6QPDmM/I0EngdbyirQwsU1LBZCwiEgb+vuDf1MKK+l
YRwyvR8XjwmvrD4jHpQPQg6T3KwQfpIlFOWmkxDlNK0LvZ5Yi5sd2SHDKGoBgvB71mGiUXxxyFpz
92A0smNtAqm3LyNiDhXLqbjaWE68iF0KrEGyytSyFkoQ4fDxZripN5jlMhKx9Frv4RgKmkCZ4WMk
eEUK6gwTmdarxTiWSDHva9SRlYB/b1NSdrf5qeJAbBGYaGciyewGfZdVPa5pKHfcrbDh/S+HNmtG
BdQ+CQm/hU09psQ+cTvEnmDBUPmZLvELNjdsFM2CXeSA9XnVgTIK/63PKdW0S81NCPaPq36GcRaS
5ePwDUJeCfTxMK4WeiK1CkgeuW5pkw/jT8e4sSEUDfV+5xFbFNLFH7ev5ZouW+r9XdbuzCogovIv
g4+djr0KJBjn4r4AKi4Ahv35z8pinl8dmEBc5A2AiwjEmkpfARBuQ+MOpBwMVM4JK/1WJMdkpZ5J
+TWbkspyKj9M8OKSE/bUBNrh4UyMLJ2/djOjXFMY4Ti49dhbyc0uw0EdAeeQU+w/XCsXpm4t5T4j
rWOTKody4YbcsGqiKZBf1hJgsso/JJqf5VTTrr6S8Tk4CDhR0l44ooHFw2lqmqLVDDZ5D8QQm7hM
zq+4NQT7qEtjyaT3YhgngXK/oDp5DtezGevHFVo7C1QjcSMPbkOZwvWm4567R7Ic0qWNDplWklaZ
zAswme9Tc7Xq6Z2IJ7t7FDgg+a0OZR+DzXFGMkfXpj1xR8BIox0gl+mZ4v16r27XZrg56B+T59v8
WWNCzRRyt8s8pdMRM2uOg1vgMjKaZgFd/QADg3jClSzg+OKSwh/PNwW9bq0DypgMFsxYkQQACePo
FZhjaJ+bEgoQ6KBLBG9EBWkOC2/zSKXrNOiRLkryLeag5XavXLZWbiVpvfbaXPnvoBze8bTI/NH9
Z+Jqx49OTC+YwVpshV7L//qEAlkQT8rGIoVbwO4ZKKIHmaVqFIAs2M2AQu2N14LuxZn8TsXx/YG8
0kPYmTV+mq7pR2R6Mxt2ZeXmCAxDyoH6q/xuyEeYFBGC6lLsoIT9EJy0cWUKIafWzARGQT9fKIl8
i1pPGz87CK+uZAwMDcJxThukJhvaGepfMNsGXbaAVck+CNDpnAb6ZCpZ6EUJfSk/1miofvXJMFo1
r6gxdd/2/yVhUMaKvACppknDuZRGMWtmczh9mgDYhQVy9NJUYiqLL2cl+dU94iIXCmaIXNg4Fy1s
kj+rxzsVfLqIuy6xDH2GQ7WqBAggq5iSYMC95EIOMF1zbhJNxgq5Lx7iqLsGyNgT49sSLnjXEVD1
uVawavGK44+b3/CSDsBT50snaYp4GFOC34xBnkVXoznkydPov4MO3Hirvd/kN8rIYgza6170Rxyw
1Kru4nZkavDzJH4bGm7NygBsoNrFpnZQQNQP4XcPvzRAn5Hd/GfYx430AgAMjMgxWX6L3RAqEHYR
74JHMuMcrrjSOwMWhdM9MWirX8utdiHFeXa9iQsJYEIW79wO/crcuIbhl3G/Je+mGyN5IdvPRYwF
tcj/vXZLHvNcjYnxXPw6cTd/mplxD+3mJouIoACrci/ThvbUsRShZm1d9acHfigosjg6ExCqLxMU
8/QwlYF/MzwnVE1S05oNi4VhQquDKT69w9xsMSD/0RuhLEHxLyztijmEvM51NG4adR0R2U3zV5zl
Xdu6S72AzdVimZWbD3R6D9v9uEUUGLjDaI9qkpv9FxoSBWpclCILRFG993zedE4vSK+fUpViCiw7
kWvLag+NUr9BMXX8vq9krqxWXbOYMgWpjA+my+CYjz97ZIfKT//yKy6DIQi1B2agtvg86vs1tA/l
k8eSiLe2mKCl3J/AL4+bhWmdx4P8JEQ91ZCmt6U/S/14/lV+3M1bJP3dlJXJgM/DX3QuyuMO8jBA
sKqOevcJvP+O4rQsUu1fSmgFUIS7GERiahjL4ycqBTo3AAR2kCpp3dxYzp/m9eftDxr+wLdT3071
lqQYnWw1LKF39kEh6mLYjONLkWSmTHzPD2qTvKWJRDv/O0rwh5jnuTGcJJX9i8GANEwfcYro+C0I
dvhbCceQwXnL1/BLUxurL7BZDjDh7+QUaaMPUhk96QMmlSgYllrS9zinQeKiAb3tlWV8Ys7+8a0D
HWHN5+1Fiakm7zvPCP5fdVL7NatUJK2ocynJnl7gqvsTifG13ynwZb2IY0PtN/mZG6Qd42umqmI8
mMMergF9f+WlUn5mjP0GEKsg+axX718kKVm9bO0BAoJasqmFbS+9Hd7Tnk7z2lnqml4Id3wXH/vm
VdrKEPlWukMw/VfR6BA6qyQuW15a1xLW+9FSZLz1KNIxb7l8jNvpFVlq0xL22Y8OrsI/sOb0hmJC
unotnyOaGy4eBVVRkXAmvji3J9n6QqpjRnRHDStR8hfBrjFjcnug0QkuRxICS9hhBypG+JDZn/Yz
cgT7fas6re+S3+90YGD8IsbY+b5SDs0E4D0df7Jso0QUGDCkB+t8xOUalJyEyQyvclII2n9g7B5R
glwZ5pVLHPIURCMWFAhGQZtkOVn8BEHHrH0/9Nd3nn5L7gSfX99IZOWfWE1ARuXF4Swr++oocpnF
maap/2i2JDN08/pcOd4YxsMRfE7ZtQBAijOrEKESVtASFbWblx4J7RJ0Ni1bhAeuuEddBPn7TM4V
6B8gEgZQ1hHLFv7BMtt5o/J6/NyHhhE9oWATtNMD10BTDEXZ7sMTrVoa6tLx25Tkqgtt2nthHDzd
ScsL2yV6f5MyP4w7DPVW/pDJsuSCgvQvT7w1L3VjYSCVLMq4XLlngmhbSJEe405QxuXc5FGC1bJD
fmjR4SVZJOYwnFT2A7q9wggoYo6cBylcTGUyBuYt5AXU/MV6rmlVTbRGWddrQecCViF7V4l7iUDd
3JTpdwMd6hJwqvhbiS3M8sw5YYrpDegw9C9wqOl+2BbhysPyk2OSlf7vz9kGczuXOFujDabH9Xmj
qMPHJ7P4vnmWye19yfrgowLfOVZ9CHaJ0jLYySFoUXeCKnpq5N5o9V5XHCLfJHQjIxR3ZCYqMYi8
+uxtprA/K9xW2YRG5wGUT5Rjt0eQs2hih5vWqlyYwGeTAccdco2GFFa+5aLNDKsJJ5VSQjoGTkvM
fNkf/vHyBA0br+xTUbW6K0GJZnj4aMaNCgDwmgOj6faWU9OgwcOwdzcmsMHKiiZ6DY44masJEsO8
H5K2yZhb4NyEIRVElDe0pkZyj2bHH8FbhDErbLjqGbfePa+mT36NdromETFEb2HF/kJH6sHv6p6f
1gXLz+K+4AuAv38x3xkQfrg7NPnbKmfstxIcV+KVK3ZBXcM3uiM+slUxdzjKvi82kKBTwzZ488z+
blwzSG8PMxsvJboO0JdmYGWdB6uNzCM+eXRq82tnZTSFUGze3nqfzXtvsY9gRONlVAEZ9EpGHDCD
9Z+4gmS1zXvMGdZvFO3BI3yXqf29E3slRKxNg2Sz9RYCc+X9yRbcVS2yD2o4RpRQ7JkwzRvutYh1
mFqZPIzYNwKmY+gqEI+4vMbqZXQ0+nbIADg5ejb9CSuQWnOpH8XHmIf1xoP7BNrwV1U+4DagiQ51
Yk6c3F59JdPzh04nqWSK5pmbBJpzxLeUyFmzvRJvZnXXwCWH37bdho7Qhj2REXUtVZgbg/xNKXlm
/mZixCMfOaDjqmfleiK+qbxgtldwAFJPPN50UtthoUmjthNmXXEeXboCFAUO9IU2WrMaodYzPsmp
T+ELJTpfvjsPFjXRx6167uVInvXpcJAK8ltZGsNjQ9E4oER+CUI1iMsZrOfe3QE3jhusk19Oa1pc
EcIjBSbiaRUq2yQ4ytqv3ocQYu8nxs00VYM0j5aoXmcS8Sc4ttSETqVEdmumfWMaoVCoLvDPT1ca
t8rYxUYUmRGQyMRg/54aNk8Pu1CMXMngBlExkGQfg5h+TguOqDGDwM61wvbdU9uCxmFnySHgFAjl
dNooPjg63vGGqZcunvQBR9erYhxtXecpg/MLhZTZbtrnDt3oYRhVLKEU4MZQlvXoXv7vcl848OCZ
tDWS3DDrMjH1JPXtUZyCYHoG28pCc300Sg+hLstqsSIVMZwQ8c83cQV7On7TfPjVs1dSrmHoKtt0
zB8xDjKWR6jbYALuzAUJPps/qC7O8a0z2gaUqYKNcK14X04xiwrUdqIFgSiZbJQLef2ZTQIqeAmH
MtfaS43f287XEkW73ExBmJoRo1+Lob5tO6wieH/qYIN8iMpTIKcKbGUcSTFOpKW08hKCkvktMGQ/
0mk/olmr3vS2v+9c11Qk4biQBE3JTxmb6b/2Ra71PCAkv+lDYgd0fdAB0MyofcOLvBjSEp6WQc4p
0ghYatgMGHdXbChX9Z03MP3HuDJ3reBZEXY12K41OrXSXP/NIEC/+vsnK/UAwuLyut3w+Opki7jT
BawObbNq9ZnSYZrkRJwneM96iZaTOScmTBiQr3tAmI2KsCD75PLWO2tD25/mxThnZwSo149O/yxi
/lN6ER3SnBGCG20YYNbnfM2kLbP6WwZ1LxeD8iFL42QgjP5lu1g6pG5LEYhrzOOSB826A4Se+8nJ
B6nK1qs2032fv3lOWuGFBH2jzHdTu46gLdaLvr1rNYVbsYrgarpdtheftQBtbqstHYPSuPKJyHiS
9caJeqkUhtaNr5A75crRlTuTqQGoTwqQzR0Bs6536gUPkmDRbKVAoFbmVRMPx9yik1kQhB9Xk5p/
1LSAJ46pK3hYrZEbViE34XOSDATRqsDOGQXB3Tfe8zAmE2SLK+C9KTturO4yBFBMzbsi0bl8+z0s
TzOBE0XERk39MyAgDokiO2YXwcpHkAuMPstOY0BnkCiBXO5055cnbA8pFKzPKiD0InS8dZiE7wAq
GCp/CzfUvxJaxtGTZmJ+WZcVaq8u97MMb2MU6W7cxLmbRe1YCUTDOvvjzKUdMFlvJ4DWtbohjvlN
FbQmMZ9sFYJEs0b9ZF18dQpUpoUapY++Qev9+W112b/6XDo4XTZKpIoG7eGVVyRkTvtY93DS5CP5
oEbMDQV7MMQiNMT/Q6D6iKpLYL/FyBeAGhS/KHfceKmwVREnSWjx95BFTs5jMxHmuRW9CnAQ/x+w
YVW/tC4vDPkhiDiA5uPrsTuy1xlMdEbk0SIs6i7sHEKgiCZyfLTNWE3ObAT+SE2+P9nOnkxzLhI4
x7UHE1TjR/sJIzWrzCWpUDnkskOTaFqOl6H7dOO41Hgumr+ae92yMMm4bMwvRGMjgf6Ro7n9d25x
sbhtildymFk+Men03951znD2Tb2U1Q7ObCJSZB+8OCLgCyMzXfInp6SiZ/BD8kefZWL1K6mGWVpb
3G7TvRg8rWRkbRJdIyOzpl8SW9Y2uW1hFVHOAgt2SZSnB4iTdTUNHS7kV0dACqCo+CXVhdrDpcPX
pwFlBBY/tDDK+PpVfh6bbQiIaCrzh+1ABjemymt1w2KVQ7Wt6xUEaEVEje9DdIKk2jgTGOcS4mOc
z+7t+nT6pVK++ICkdbAw8+GjCTvMeIuT1HBdBMnq74Yvar/EN8NQiLTg45JK0cpNabUa9dhFodPA
54LwjhgKR3Y0yQD2Ajy3IOedshL3UZrOtzJJeSfJg1ksEaAEAmJt9ORzLxp1L/K1mUYlmIIGN+ym
fV0F9BnDpf6bxIBKdTlx4Lj7X6FG5ESVHZZdFaRddYM/vP0ZF8YU2RdgRZUPPlgU+q/ulU90Ko+p
VPLas4iiHoytwYD1MD1Oho7lxtqza9t2KXK7VhfRMj6lcRb+kx5Xkh7CYoc9pwmhuV2IFSyYs63q
cLNvsvc5ZXWkvKTT/G1KkFMXXpb4ZepuOhZqEjZ2uhD5RomZh+akx7To1ggQzaTI6AgqC70kYwMz
RFTW8ATmacGQAgR31VZh7P0QiHTsnIsy2kHKQEd0DpN8w1QG5MxJe8d8KSa5VSOHxyZVP40C2Ll5
U9tokRHqi7mV7YmKQ39kpFbraLEG6+omipNAMY2O95Ae5LViBJLKo9OC614J/42o/zhO5G7ly/FE
w5S5CAclhfo8Uq/HvT4yf23adjmwAPn+mvN55pFSOvNl/dhZhSUFPOgHOcW/DyNGSFHqHozyMdHB
9EGLa22fLzGjHkT9E/tsi+MxU7G1KMtoFexobwYCVQgoIJ9x+nCW3I9sC3lRYanlxJ8H6fiy1jTw
ofnrFn/jodTPF42KLZri1qA8iLeyoMYIt/DX6h0Mpv9PdwssKUgRKM4XFo/y5/wRYFsIXMLzJokv
VU7NDfXMp5NqVHpBBg9tiBQ2iu3ZNui8aN21GlQvUT8ghVajLLA6r87hDyaAo7jKm82vOC84LmRF
YUxESX7Au1H8bk/IP+Sm+olauEOXZCpUQLP1JYPal1Iw6zkFYAj8FW+zHOaMAa+r/1hiFYrmQVcv
Huq0yXeaOHCWI4eWl3MwVceTzVjd7IjoNB2gJNwAGhVofCnDyOj/YA24Bskb8QIs7+M6Ye7RBG1t
2FfaSlVhfpeHQHinRSpdYPF8N2oe33IyQf8=
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw1n;
use gw1n.components.all;

entity PSRAM_Memory_Interface_HS_Top is
port(
  clk :  in std_logic;
  memory_clk :  in std_logic;
  pll_lock :  in std_logic;
  rst_n :  in std_logic;
  O_psram_ck :  out std_logic_vector(1 downto 0);
  O_psram_ck_n :  out std_logic_vector(1 downto 0);
  IO_psram_dq :  inout std_logic_vector(15 downto 0);
  IO_psram_rwds :  inout std_logic_vector(1 downto 0);
  O_psram_cs_n :  out std_logic_vector(1 downto 0);
  O_psram_reset_n :  out std_logic_vector(1 downto 0);
  wr_data :  in std_logic_vector(63 downto 0);
  rd_data :  out std_logic_vector(63 downto 0);
  rd_data_valid :  out std_logic;
  addr :  in std_logic_vector(20 downto 0);
  cmd :  in std_logic;
  cmd_en :  in std_logic;
  init_calib :  out std_logic;
  clk_out :  out std_logic;
  data_mask :  in std_logic_vector(7 downto 0));
end PSRAM_Memory_Interface_HS_Top;
architecture beh of PSRAM_Memory_Interface_HS_Top is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
  signal NN_0 : std_logic;
  signal NN_1 : std_logic;
component \~psram_top.PSRAM_Memory_Interface_HS_Top\
port(
  memory_clk: in std_logic;
  GND_0: in std_logic;
  rst_n: in std_logic;
  pll_lock: in std_logic;
  VCC_0: in std_logic;
  cmd: in std_logic;
  cmd_en: in std_logic;
  clk: in std_logic;
  wr_data : in std_logic_vector(63 downto 0);
  addr : in std_logic_vector(20 downto 0);
  data_mask : in std_logic_vector(7 downto 0);
  clk_out: out std_logic;
  rd_data_valid: out std_logic;
  init_calib: out std_logic;
  rd_data : out std_logic_vector(63 downto 0);
  O_psram_ck : out std_logic_vector(1 downto 0);
  O_psram_ck_n : out std_logic_vector(1 downto 0);
  O_psram_cs_n : out std_logic_vector(1 downto 0);
  O_psram_reset_n : out std_logic_vector(1 downto 1);
  IO_psram_dq : inout std_logic_vector(15 downto 0);
  IO_psram_rwds : inout std_logic_vector(1 downto 0));
end component;
begin
GND_s5: GND
port map (
  G => GND_0);
VCC_s4: VCC
port map (
  V => VCC_0);
GSR_30: GSR
port map (
  GSRI => VCC_0);
u_psram_top: \~psram_top.PSRAM_Memory_Interface_HS_Top\
port map(
  memory_clk => memory_clk,
  GND_0 => GND_0,
  rst_n => rst_n,
  pll_lock => pll_lock,
  VCC_0 => VCC_0,
  cmd => cmd,
  cmd_en => cmd_en,
  clk => clk,
  wr_data(63 downto 0) => wr_data(63 downto 0),
  addr(20 downto 0) => addr(20 downto 0),
  data_mask(7 downto 0) => data_mask(7 downto 0),
  clk_out => NN_0,
  rd_data_valid => rd_data_valid,
  init_calib => NN_1,
  rd_data(63 downto 0) => rd_data(63 downto 0),
  O_psram_ck(1 downto 0) => O_psram_ck(1 downto 0),
  O_psram_ck_n(1 downto 0) => O_psram_ck_n(1 downto 0),
  O_psram_cs_n(1 downto 0) => O_psram_cs_n(1 downto 0),
  O_psram_reset_n(1) => NN,
  IO_psram_dq(15 downto 0) => IO_psram_dq(15 downto 0),
  IO_psram_rwds(1 downto 0) => IO_psram_rwds(1 downto 0));
  O_psram_reset_n(0) <= NN;
  O_psram_reset_n(1) <= NN;
  clk_out <= NN_0;
  init_calib <= NN_1;
end beh;
