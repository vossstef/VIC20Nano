--
--Written by GowinSynthesis
--Tool Version "V1.9.10 (64-bit)"
--Tue Aug 13 12:31:06 2024

--Source file index table:
--file0 "\C:/Users/stefa/Documents/VIC20Nano/src/fifo_sc_hs/temp/FIFO_SC/fifo_sc_hs_define.v"
--file1 "\C:/Users/stefa/Documents/VIC20Nano/src/fifo_sc_hs/temp/FIFO_SC/fifo_sc_hs_parameter.v"
--file2 "\C:/Gowin/Gowin_V1.9.10_x64/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs.v"
--file3 "\C:/Gowin/Gowin_V1.9.10_x64/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs_top.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
c8pz6+gH9HLYNZcBwk2+tJbYjm5y+qGe7o5nU4kib2qu7Y8sIi3XI6RTFRdCbn80IkWWfjSw+XvG
8L7fnWwDPvhvgu64SJY8pyYleLwzLBGevFGwGkEf1HRYjnkqaxHbSb+zzteZRBeOTh5bWRI9bi7S
Z3o/J/6c33/nR1yEJa105wxfwu14h4hWUFbBHcEbplLLe9Ae0vFdyuFWFpGhSAXzuONPY57roh3r
km5OJ515H9BkGCUq3ZLAljQoM9H7SRTMqyvA/VMfz/dN0w52e5BUgt/C1g7bVlpACu1+c9HckNya
kpXGbWxpUYnOA3BelzlfC5j5swPBaso9vuMgSg==

`protect encoding=(enctype="base64", line_length=76, bytes=15360)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
AAN22e6jl7D5EeJYqz7MfHFoKkz1MBcuT47XDJwWIkzVlClOQ79w+upKpBHav4wtDkzlSV/Ip9eX
yKMKx4wXL0RrB5pSdS/f7ACxVZfVRlrzD0pHAX6qoDW9bpQCSFvSlAoG4vyNyimDDIPTSsQAGQK2
o2GK84XE1CxL95bkyiQE1hpktbgIMWi9CCAGSR7M42Y0pF2vvxjSxE/33lYAZ8UjgVkPwaKVW7Y+
Wdiz55RTbC9O3GHub4SPrOz7MLS4Sz3qqnPiv5vuJ8u3yN09WQSwNoDaWRUzQbiBlALvhTtAJ2ZV
krwikYD+GdLKWc2bRCIGn/S7i9pYqVgWJkwW0dW/8YdZ7nHXImGI8VNFmbSbPxmxQwGHi7q8qgym
IikeQqobmwrwAa7gIeOrAxu8Ckl4r7JIbyJsDOlbJ+8rHJ0SvjWAxfsgU4pn7ndx456tkD2YrGTh
B8w4j9SG4HXUeWBu7AVgZmM10IaANRNvcsd1kftrjnL+90BlPprzkYQyByCwqP/XuBJ2LWf6Gzrf
tyek3RisgmdIiabgoUM61vracgMQEPsDIdmQaoBOsnkGBvoTH7+J8NAZuvKXNkmcvqHVXjxl9rXp
/phFyXjVwFmFNvQ0ABEW9E5ZieQKovIrLWJ19Ql180avasSaM91fRZ4j9oWi4uo0+kl4/nvwqP/8
2n5ACI0DhMDsVgxgSrEpBv0KMZ1+F3jDS1SFDwwQ/9Ogr44T/W8Hmd6ZDwDepr/f9GVaQ3aqHXld
etKvYp3kBWh3ScOHVUoO8W0n+uP7cEfT3rIsXHiBbiDn8ur0Mx2dUkeXkpFgGOtUOmm2aje381Lh
qWSuTlZNUHg++x5wWywvEqB3fWbOx9CeRxzCQjKsnuNxWUnA6Rts1UWAl/YEgcN5GRUaGCK6bWDR
4wO1at8/CVAKyPKAfI3SyPJCF1R5mmC7CiacYm+v5kgy5J0VY9RA9plNlhWQ72DVpRtZmTorkR5s
Iat7HaOfrGraUcxdKQ1tgfHmH+S3MuokAmI53/WCjtnKE6iKqh1rfmBsKZr/kCb05wyud3wM6zmL
lHEXXC9SknkqaDqYUdEXvO/kG7982CBelaG6yPBJmx9CFiiomUi/fz3MSXE6Zm6zFdk4BulBkjOc
TgpN+7KisuwHiiQLe1EC90u5jeXPfRkfpiDECbA8SXVDMgEE8/nFmz/6yD25y3Rzya7YmjCOTe+J
xvpPZt6RsGOw+HuohYo2q0xyUlJV/Xdpko91CHUjuQ4ern8U7rEkQlohQYxPrs+8uGt9dJlfZz2v
JHNo44caYI15VMgZXyP/IVjGmbSp7oOwPc1OMPMaGHGd8HRtNnbhMTB12RROusfZQ2krw7TjzaCF
ZKS6n8lbdSpYVVzW7+O1jCpJca4Gv6o60pJENJLAu6lRQJ2ac/yUzS43CQ7PKmiDPGTCU9NmnIpF
9aZsQ9MI6mzpu0syw9Hnr0MZj2QwMaqbsVVPvrUkTCx55okg8RMGaM8JvSrYBQGfM1tZR43e1fL8
T3AmLpz2rn1C9ZK9piydgcqBUgw3m5r8wWTWgY/UybJHHbSe3/gsQKTMC8jw512gAXkuZ4HUi6Fn
JUlTWahkhxNYO2+qtuOIy4AltoAG7jr3x8S0ixRqDWAZ1swTPXxQwaPfI5ey1i97tSIzRgKuUDnq
0uzU7Oi7uB2nJSPO/4mSj0Y60xiQTse32m8aRY1Jn1MP0exjZpfT+4c5ju4AJNqIJk7i2XF+ine0
5m2Bn3eaGGHCbjdknBYIGLsfDNL+d+amE0UQtZqe2ea9G265tK8MNRT4vEfmviE8YH7UxSJnkIzm
li7KizsWBVQHo2WPMm/dbJYWySrE+1bcREvylHkBA+O2gOh5+SIye3bEbIK5XBDBQJ0ludW6oTiG
Lf30UUeW39zRzSh0inGG7YrwwBT0sGaUeQuhzMhqfPReAUWPp0nXIxMZbEQE5v2kkfIRNe9gXSZT
pR8Wm3VySjU3ZfioJGpuLYDlQsbIH36pE8sibqOcHIFUwR3QpXL9S0Lk9vOJm37+b/+nSKu6MgmI
k8lAbWZQTemjp3J9/aoPbodLIUHbJc0rxuqYuqKeCqgYUVUlqBlzBAUhHE5VrFJoBO5iHvX+NPCy
Fs8RPVL2XzE3d5MjDQGw+4daHeWaWd4bU7Wigbtfa0ezcZmRnoiKwvroCX7SjkZo9PiMEjS0vS+s
j2cNbTRBEVv/02z+5rLaArqD4HdbTixvgY7xA2E2jtODeiYQd90gJCaS/s5tg8f88/XWwlHjSeCL
D6FmuZ6Js/oAObzcSByNl52kRdPoQmfM77/cBCIcDTe2ydvNwWgHHh7+e/A7Uq1k+E2kJiVe+XV/
xLrG6fqNk6k/PzMX9mESEpXZKx2hJ74SUmiX8ADM1s6UdepL6SaYHaYqAngKk9Ur4teq0OjJTa94
eL3+Rq+SSaJz4RrQPUlM5k/zUfHdCLZt5DSbfhCFHRQRLQKB2h/BzUcYtoEAHGDxIgWDz5GeGi/E
XlCQqVjAD1E9XhyLkTeM0abYzWgEwkJNcCvmOnUYSqXE/VRtp5VEOf/QNKFRj8aNCinCIMw6Ig7e
mat1HrZ+CrzajFUyjTNN31jJCLh+1SjAs38vqvqdiXBFoiVU46Tyulr9rqvHbVcaJKeA87e/3Am5
0LzUmfgg25peeFyByYzIqJ017ypNUoQjJCeCXB+A7Ruhn4MQEcBrCJVnaRVUECspeRSPXPD8ivrl
5WB88yDUOfunOP3YrHmZDXikSwXVyXI1NqYOGM2EeIMWpCmbQ/cQ6MNxRTHetlIXS8ihsGOIYnaj
gIMPy7b1fNTOUu4lq+B1QP2ApF4v/bOngnoqFTpiYvScp1k6UZ2wJp9n/XTEbJo6536Ttf0BY49k
io96QoFw2zy9ooKG/TKwlZLjTJKKRHUvI35lmww/JSDv9GdPPA0OHgZAHkF3I+ih8BiOQK6GPGk0
Gp0BGThlB7H36AJsqH2UA35ERakll70LEMQhgtfmb+kynKXBoG9R9eRefgtBtaYH1hP22gWbDHZ9
X75UF5vUEONG1xNLUJf/FaHuwy95mjHPCh7HnKrzCAdCb/Ws5D4ieWpOiXDEFEDLdSN3Itg6uwJM
54T/1eBiXMhIN4ckAYvh0L6+oYcvNTaS3evz/R5YPzXisb5l58oaqxMzPhUSpdh+B0HRHL8WNcoA
OJA7HYFIbguFARSyrksJs+yY4vZ5QXQBcPn4EjMuc/flbctDQ5UmPDFOJTqNHj6M9tRvlZ4xBf7t
TJ5+my0kPPlj+30Y7GSTM61twb57xZ3Vf8MJqZHY01Ef3s+ANtAOHIkP2s5TDqswZgYrvUnqNl/9
EClqTHHgk0cZDp8EPfFUasveeYFuUv+oEh1Vot/m4mrSYnbBNyrsXX9IW6eYRJmB4L7KCBtCVMbT
xKwYBgqx4HP14eyJhit16iRHyjCfbOQQ+Le1hW/SL00II9JHSN5KR2fAubqy0s5P92BS6FIYVVL8
w0B90cd5jrKcZcDJfTgJrM7h7jB+OAoQR3e5VtXUMSAqjby1SqnzHJzI3Qa6uMlz1gTl7iUBGTYy
OrHdOyIRWs8uqQopd0jLwpYKW0H0QM08urVrYuKsNsBk69OkNGyiJHZfqOdGQnpqIo8cEzYgeRyt
cx54fudEGrDbmpsuP9AdjsU8WLhPqoazCSnIg3faqY4L3NHj9cPf+Vu1+rF+nuoMQGiQQPu9+m0O
ZPu1nTZZkVC+bP94HKNACLozvO5HnJDprXfMV+o8bk+5vd9o1xzAi8uJ5VqeKqRxXfA+UTFwIRaJ
2z2XyPQmT16/zaq2YYBOtcO71ib6XerBnMxGDHe/tqHhwbIC7i9yUmkTORr03B/FSmRMKcQSEiIp
PJ8/uP7zJBpmwDTr8uDt85bMZTQFP3mgc0KXK14c+gZOpl91va0N87L3Uc/tLdbi+iNZNHNxUzd9
K1qDQivrPJ9IDIA+pvHg/PvMTdSES+MlQA5ck7naBhN108ogIwXARSwk1PmhC7feGN9p7SP0DjxX
4oS1CXIPrfe8a7eaPnzv7oboXKwSlpIaCE7r7O/EDw4JABoh8rxdYPWL91v4FgATCQGPODS73UL9
v+RWpk9xBrtT1wRRyDVNCYdEXSvImgxYyEjSTVygDlqDZEtuFOewXxocfE9/l+WqGPqBnCIzkcgp
vQXHw9yjIvJ4B2KPq9dOKPULuiYy8zwmqRev478+JCecH1XCTW/5U8HqZAjvqEUMlfGGH0eycK9j
2n74EP8q9QJ+BGzMhAJv52X+JP5SFGHjJK7pqk4JGMlJk9Rk+zt78TEf/lZZcaddpl/sMK16Usv+
JpnSGFsweHRbk1o/iuNpxFfmtH0Idp9pTBGd+HEKlLgkulq63JL2ckJ6CLb9IZVgJaBz19X01Hh0
/t5wYD0WT2lap0ST2F5QeCWSUG8/oIxVNrdTD7QNJjE3GgWkY1CvZzWlTjYNnLkRkwV5cKCvTubO
Xbf5Hpu/ULBv9R1Pp+7rm6FWkkdobMg0Q+Q/meGVY5So5myAQIyS+gUFtCFCqC15RGLpO9arLLYn
bJRuaZmaup5vfIgcBchiOxu6PX07KMNik6ESeq70CArJji8k2wv6lQ+OMugkE7oWSSwj/4DvI2q3
vpRfhb8/RJR2uSTrz87YYh16htOV0JN9JL5zcLQ27WVG5J5cNezzWQglckycAV7oSgtmB/GDpF/Z
le0uRwnJJB7vuEKh+oJxtmDJsDjMLb1hLUPnvKA131OYj3ifRQEB6CukCe7VvvlUTtCQKK1DgBC5
OOjCVhJ8uHggW4QzJ1aZa2HnwaUAd1hlgD1qFcKvUhjFSwjkms52AupN0HZju3E8FzldA71LJDrM
L/xgNboY6fepPAJYtn5sJ4CBWxLQwr4rK9Toa4SA2qJmJ2qFlMsrN9cdqCAH9/jNoqWdi0mwCIVz
/D3y7aaTsBTiPBg8ECOKeOKu3uTS6IwEbOWWFKCYEc8MKovTnKqSvDVJ7JtqaM4n51QFio2hkxJL
27ewmiFlHfFT5ItUpJjwdpSpp0licZVn9tJxn7pt3C/l5gEzxSSpnVdiMOkoENQZK6fXGzUsIr7k
u1Scw0hyTl37Ho3cFEI9OQdpTxTtszPrD3dSd62Axcc7oNC3cwCAlvKgYssdrGd6dzuonO1KhdBV
aBrM7IPNg0Mpi6QBSWlzMjmFjO/iPdA2/UaWgUDnUBEG8BOXObN7ffUSJvh2DZ76FgHAu5slzApv
OVLQD9YcJD1qJEoviCuypUQxI+p0Ch6W5E43PQ5fQNllk9TcmMis/PzHAv55gtl6l4VwRy94eYxA
YzWm7s92wRyQrv4cEdUF2NYpG3r3PzZRQrO3Yu5Xs49tFb115BScBhw6ZPq/onbLct3wWc6vxBhh
XpVPA/BuzMQA+vzeW+Ca0MaNtJfMpvSFm+x8sJAu7/sH6iWcDPg3nUTNA73WDfMuX+tFlBUDgm0o
AKcyNC0kq4vDGOzxft47/K/X2DMygsajd41DxcBhnNGI8sCW7JGTBBcUhyJde8i8Yyt6va5wcJZc
d1mIS0ulJOngx8FnzHu6c92BgYoEYlXU6Cxpwz0XEIdefNS0v4h/klCjGKh5YLdQXnw+oVW4hw+l
fgEKI6ssmWp6nwcStq66yA5FfvcR0+e8rCjO2jTzRoeTSZBs816vBqrkqnMtnMeZYMH27CfCrGWy
cmKU+7nYyR8z73LSuuuj8PCLGCHMLhW9O71B+ZRINKRfg/8BXvgnjF+nPvhMZAMl71Vg0egjiOME
vfwcmkKWE7lnlm9HPBNtNkGk+e2cgikWgDlWY9MnhCTtq35eIsiWPFnmBCpHPVLG9BeDx0hcg88Q
0UrRZbFlAT78WARrol+O3pHM51h16lEYELoMBVi+b14stuJYvqep7jAD+cHVhVyHZVm/Smdz6ZMp
wkfLVeGE4cSIOBm0FaYxpMjG3pK/bQflmC0TPkqV+WNO6y49ywpVP9R/R83d/njUGfxxkT1W7eiF
QuAHyzKtQXCJa8MX9CTAAlBYUPqSN8YB0IwsGQhcwENmnSw0wP0wxgfI0wSwC5d01ZxgaYaw7C+H
R2L7X940AQsH2AsjXPY5hvd/BbCnnHurRuKcCMsQ9Men8dXRrugH8E0Q74G0SkSMCzULa2yKuhY1
VbLj0+eQWwPl+GftvLCPNi5ZPpH+IQFxgNV7OX7SUFB25gfNbqbtBhJovSmf6G72yLiHtpmarhHT
I/m9Lv7t1NibVj475mivIgm1lzG0SlG+J8Q5LA9t9mdAPhiHk1tJzkAuHDxLviagvnQCYqCbW+ay
/Lv4+q6LN1eFKMDEaI0mKkM5UvDasEn2trvBj1wX54GUFC6rxYyLBI+gZmcLhvGh7+2Gv1kzSleB
paiwXwKqM33O/73SnTZlgJz6wJIfbRaMFqB5wvKxzgimdxI2sbAdioE6Px9ywCqwnpLG2FV0qih2
9RXKkd9r9oQl7WwtGgrr4k8HWs1kDROopKtvRLlkkcn2h40tfJ/ZRFc+GGdhEz8iX94w7Aetk+rb
RUFqDMMWlxr69NoO9IyTMwtFDltz430r1p3N32p5DjcVpFcLN4gP9XCXB9sHAmueK90ZcjxriKU/
uFbL9JlZs2OVFZ3RKzQbHOeVmkqbQ5Z2OI6j0DXFxqJwI20Dd9FzhIWlaWjDlIMew6l8Ky1egQWT
gmHgyK+GekIGQDR9eywLPuZpFvwDTxR2PDbvSUxzSXN7Ecr/M0FyVHps4WdYsk13/uy//8GlHAPG
jm3/eovWjMIWc2+ATLdQQjGaq9xjQs9mFyadY/qby/UlVwqz5wMo9SiyIwN6MwqhxbF12UshISt4
Tcg9QQewlWchI0WesgnGh5Pl3iDZuR4bO/X1dmiJqmZg4XVGKowq9JJY8VhNEO/Debwet702Pbjz
OJK9t9SICi5mrNcvmzCLRwYFRWgDUjCr5VxDyll8tmFjX4DMMsvpqp+wHVmqWHmpFXxZ/jWPepM3
n6Gzt7RsJ7SiLKya2/H/p/xRnOmEDf3V1tzm1Pwj5EwigmF1QKS70htEKGyCdn+X2CL6XCgESadi
EcAuEewHGHsPoMsSNQykxmlMki4yjsl4Yts+gWS5uaoV/Dc0DXMG11UwtENLI0qSYZVe/77c/wM5
vTVbLB15KiDlmw7WJ+gaNSEZQjTYKRm9dcAmAbV/xSV2hIk5zS8EciKUFo8z64FatHuAYTaOVNv3
7RgY317M4tei7ax+1uqiNzytY4IqXAG19c16yZONPtt/4qlntPwPl0fO7D3pyU4Mm1Ygpvp+4y9q
waq2B/g4Y4RVMQ+J+ECkiP+minFG+cSJZhK/kQLEuKrrsvL4BSwP0kMty38uEP5y0/6P+S6ImDQx
6m8PH31CyXYBhvAonZw/9r88g3QDJM/gn9BylOj0X2LeIMjNe7yIEmR6rUJjbVmcj4hqKJnhrPuo
fSznNKcCV1fQZEHZEu1BSWeH2S8Ybd2RmEeBOs6Ogb/amu1XKTQ93PuauXfZfkxxhaSe5xCf5BVf
+482hYOnaEx+YT1MFN4YMaUTmL28FsLmLzvVTmIRBrUGtr1vfLYDG3Lra1A+ScvnujcryT7YSFvu
5n9CTmUQmO4dsRzB1DLiSjy6UvwOUgT/17nJtgIEJLrGaGimtSOOGhusUU0IPiUOVYujem2PGGcC
+w1Ck6TR6Q/SN/3A3i5F0vLFQ2POzVUL/pKDG+9FRVlvRNm+cy0zEea+JScLwgoMn2Rk43mFexA+
lxg7Cj2aNEdi4RmpzbAKjs19fSTe1FEwQUuysBrl2gwY8fhmR8rcE6ksdIkgM3K3NEz1loL29ijQ
bRtxI/oOcx7SITmj6DIMLhfTNXjuki32ooanSvlqZ6r8HT0VxpPLMb1GayoIJBJntRd7M6+f4jll
377jyzay0yZehJf7VnPiQJK9KFJ1OgdXVSI9hwjfvNcIULYNNwoLbs+VADIenjKcY9KJq7OIs46E
Jy22d4MQzMIns4vXAZS9IpX4ZGuMsHV0k5NNUKnE6oyulCDPwrb0A+A4G5yHswAUE23ui2fv9m6s
x5lFDiV8eEn/A6/dzQ+RFPanEti2KUBRB1+9/xmdmzPvlwLU69I11NbyBZ4DiZ+yJW0dbnbGZIuS
qIGUtfQkIxR9KttumYQI680jsZsdXbEP9OKWcPs24itjM6kMeQO4D2ZoXPm9A4yX4iOb1VW4yPoK
qiBI8kVLS6HLeWl8B+LheHpI/jiKa1U7URIS3hVUYKVk6TdwtFmr4bZO+6U1LYEPENZP9PCb4BJg
sFFYAb7ALgM8YJaSloijfi0uYRCvFspmBTBdyP5tgVyQX2pnptfunitURZQp3mSm9uZLtQd1fUie
N6xDyTtzXF2v0OzoJE2E0SLexm8RZcIZIG/3eovgL4JoFykoMvbSk6g5aqU/RCPw+aesWBklDcFG
a7u+mCopmbBHwEGXw8ALOwRfS5Ipv9Sz2afx52VcBlGFyonauhT8Pa4Ssv7qyDdQQ1IH964KDwQ0
CY3nieDr4Nu5BG9a2r0R+mE9WjoQzaaMs0BAUsXA2sHPdToZTcXsJj+01BT6iDz3irI76sPC5NU5
G8x2QZUZajkjnJOlkouCtdoR/fm+YWbCWeGdzT1u6g3w1+++EEPYvVkpjAL86z10f+FY5g3Vfkm7
Nqif2XG3DcNmVpBUuzouPXpdkw58KDc2QTPYmppYTvcc+x+6PkQlIzBULwiVEgZqyDG2pWMpweI9
N6Y77ZCJNLVNvkMhPt+8q25MKkLnI7asmhnSZc5fM/+H9Xf6Idl9Xirwz9vOYChBtAU3o/8YG8eC
jPuZ3Q5+fkkvV96V0eAm7OjVOzFchJQqN4XnzAfrlpqsvBA7aSw5hRLHJqxxaoGQ+ihBzTHTVDPL
KMCj1xy11Q7nOCoqizQ8qM+73kNyZwr98ytkioh+F/XzBsMmXT9s89gWX610MGkQBLLx+mBejIq5
zm8owyTjqobXK/Pau0+qBg0krkjPkh5gSEhLhAjh+94CRChR1IhgzZSynh0upfSz8F4fPOw/82lU
VWW9vI2LNWQDm9MwsmghOdthMbZc/Dbh60k+TTaJaNXuXEE1xtxbQik/HvYIEblN8Ix4LJmQcnev
K0GFw+gVWbQqr4hUMoc4j25RvFbuD/UniCgAWLxNZpfuvs9shuOi3yB/RmcmD3PmV4HNOkwlJhzC
KPP51TKW5Fm3Ba/oasXa9B+ZpFGhT6nwJq7tV33WCrt3U+mFs85MLJPWK56TqzD/crXoJDuD+Q2F
JAcf8/ATagF4x5r2SBv0PidjDDE13LHC2XX5MegmzRm5XnlpN1r0uURbHtjIb4K06DaFgPQySUse
lODvjuT1+3RAd78pp2SFeltsQnIFS1E3oPd48mDYcXtEEjx8ANSAV+onk9pybJHu9gSkaV7dx6VB
B7w+Pn0SC3pEtvmbd+QgGSY4s4aQ1myWz/9TeWbqLQ5mq0d/j8YPA5Q1pBV3SZYqLQfYKaJJZwDp
tKFhKocEhdmtuWpSQybcAj24hITLS60PtCyT9Snzwh6yuVG2nekJU3keiNpVgjcDyNE8clMO+LHt
ytiz6E9+uWDTOYUVT9I67wIqqCSPAZ+Tokc5O+ZnraRubLKUaj47PLMuX4j97QsubEAKQ2QRVWn5
rBa7zpIF64dvs85cbpar+WavNKsNRwcZEK+qf/wtvCiSoh/hbcox4rNM8MPVS+wdvF7LU68sFyRC
zdbD2CP1o9v5XZSykZceTUCf1z1rXL46nmDiR2jOUtjCB4gqMSJ+BfoSi3VsLMMv1zfqvUHsPLjH
lH9tgMr8acYGvP3xqSMrniyL+2Czu2Iq78IatPRwhGAyZN9UYEI12fwGQZTyoRdf5gGzjKuO7muc
87KVg2ps9eD4yIfXmnz0FsNa2I+7djSN1L/4v4iuxI6rDYanUJT5O/1GPqGfKDn0Aiy91eGMEp5D
aYyhR0rkfnSJL9yRCU9i7Xcdc6I1vRH7sFczbDgl8Jx+chTpwh3tXLjPilFEh1gAYqyaZR6KimBp
PaamYCWQSotZcRy5s25o36Xb8jVIgwMLnztTC7BLJOkG0UzzkWGhjyFWZwcrSopoyK59VvJx4fmU
2rsfeBxXao4XUuFdwgfuxZ5oTAeSAEwLs99w7BqgieHZCA3ZP/oIP2o1kmd+rJKLa8byPpMJbTjF
6QM9a6NC2EI09zXc0jTfLEB1nbag6WQx/1gzlK2HzFCrkdbk9Ys7FiwCpYnht2IdQPN2NlvdyoHH
rgIQ/3wnuihsp/KCJ2ioOQ9fVmgAEoACdA8EPqAo0yPKYaXycblR2DWLQCwTHXP3GUHFVthgoqHG
xfoYqFfOCaBOuKoBcohnhocZMQddv59Jq5GsikDVwgNks9f9OtdpC8VYDuZxjMF4Yj2LsN5rAZHy
POnnk1kluImFIwon9NdoOlW1gwt1ZT6ZJv5OMd+cZQfNIJUbXi5L5PaJceD6D0IAsdJ7BKCC6E6A
8YYXNnwVBXU30GSLqmyOIji/AUh18Xh4rHZQdIIyV8v/L0xys5P/O9Y7Fu1JvR2f/ZPi8t+3MMS9
9fVVGwcW+QtYb/m4LniUCP+BqgyImnA/47J0kOlY05l38rniBSvDaD70jZ6+8YC5X3TAFABQpD+k
7CMCDjW1fHWN+MOuWNs5I0Oud2cfAp1z5crFyKNDCmOgmn9MtWtQ3c78D3KB7Xw6XfDRiD4PeXSr
pXz55ZP7gkHuBIwLNpBOdWA56vWLiMOEqhOoNUIdZmHo7ya1J4LcSD62NNIUijKdKVXWXVFzes9F
eaDfMo4dObyqTJ5HgEJIR/BD9Fg+J37nkPkGj7tBjorTo7opTZTeEuA1cNjy1A3tjiGn85ewNhaE
jinbXv+SEJrI61KskMCGrtip3ubJ3icSWrItDf/+M/GEXU2zziSoHJKWADtzubgoin/QX4K+jJh4
uFDvFaE9AvVEjfuHKJXOwbGNy3SPs/4LTDw8r+qceEzx91XHDJQyJNe7V9XJherRtOg9caTXBa+M
lDrRWUgXa1RREmrjvBeQzk6gkcv+X7RqykmUFqNWgRgdieo1B7LBwYHZv6wzE7NZp7gdTOs0rU4R
vQpCQV3uZfPDagnQC7rzk0WnSiS2+XfZfHv0fCvrdlVFOt3gp7YmycsbzSYorNzuddRl5fLVzaHG
46jXQiAjUKw006AWN8urZgmAld9exoXdkvgy5uVJ5aD/kZieNWZTQbQ8LkbiJ++lv/Rlhk4AkBjf
qgA5BUG/0JREDaCHJ31QScYelCLhXCCQUd5atdaoB5mi1eMPnrr9KGX0gYbxPwD9uauRCof4tB3S
yDxYe7sFbZuciqYceFIGKH6+MSI73v4EhaSpiSBfypmX8CwpJs7wUi10MULQ9hCM3L7CtsKpysn0
DRV2ISDHp0rQJUcr5L20/yCJ6W1+PNGf+4fPx00cmnmVDvGueLjf/M0kBH9mGa/eXx715d0IR8Gd
meASKb0IWMzzjw1fwDz6/zvv0Akg0NxvvmMWbqb6BD5KS9Y122Sun6gyBbu5IAvpkE3et32XAwlk
2PHuIqdFx3iwfFr/mT84MGu7jCF/v1SYcPlpTOHXcIiY5o55aao9csHK1V/1CsYj+xTl1DKHk5CI
vbvDA9IGOKVzSn5EsS6AVSSd0s1CRJYE6FaD/1NlUVluoIngHflcb6gtftxrWsKObL9Le0ZwoK+p
LK5UWyjNmyA7BGNwU/c3nyYqqnaLeWHQKKB2fBya2u60oiuC5u7qg88y673WIT+M57ntPWtuCmEk
wZp8WC0fjQNGm8Wa+WTWjKkHcRk85Lj0S1Gmi2DDOvapeqggeNrkbrirW1GK/82vGp/Qa8gFFRHS
aDHCMGvI/4bVuvDMCECm3KrH5b1lceQgSsj5X3jKw4gBjvE+Tysbmqf1Q/7mtuTlfmOv4r3+lhhX
yR+3meIYt6riUbZyByDfBswyAsruIKRI1JDZe1KevfaosNVgNa/zFh+zRPapuobZabhTy1YAjE0T
LPn+NsyiZNyZF9sX8f+Fdx/XhrZYtuCwrPVjppFFHL55HGOcC1KYQ/NGN8REX5KYOIG6/hLLj2bw
6J/y0AzDKGjWvKgHWIvRTUC1IFkGSCMAu3BvFy9LkzWLIj9meg6s/IYmXXgEAunyhkBap9WaulXD
NW0jxOeRgrlZNgt8ijd0CrWfD0Bw+qKK1ko63sgQkJgZgX4iA/Qh6WUUKSntJfkIYUekgT9ERe4H
/+EQpDZBB8TFHcZd+dO0gkX+RYw6fusKktGk96A9Z1JZlQTSYcLZib3QoGBQJYm5wJSKA8xPTJxU
aOATJtABO/L1qi/ID33hC5Dnf7jTi1S8ac/UNWnNL8kDLXYgHsAuTvGrYzetOP0Iw9KTzOTulgrz
Gwkr0NrjyAt0AFcAlx3Fdlv/XAZfJ3HHRbQoI9K7fhcrYi2NwFP1/S4/InfJ7ULZ1SYplD1z2CBt
qh+1vOMshzDg9PjhzOnJ3B+rergzb1+PUFy28JbsbA7Eorb0jm+3KTKojfe1UKArUgEFZEWgBdSd
wrm7fM7PHD8Q/eER0uwrjmdx6Eu7TiKI1kQ92syaQ01IX64ilgpzVD2HY7WbazbESPlb3o2Kaatu
RqyDSsYxcI760ZpBFQU2fgbJ1w1kyiDfll7ma4aw/EMS1xpe8YIGTqsRXpglmJwXK+PWkLc7xUPL
r2vfpH9RtSfAPlBzQIEQuLggeSdUUQZQoIWefhd7Dpj7mDaQMoylo7f5gn4klSyxwwccOT7rjfvS
qHmkQbZkvjUADNWizBZZpaLtM7YrdPV06hOlEIRCps9t4MEeXKqsdwtWbtsTzx80U9f1lZpxHHXg
BXJI5Q7izdJm1dibOa7K665AgoI3vULk02ACj/pVCJmnlauqmBzCEs+zoYaTG3CznXtUq2Lus1a8
Ptequ2cKrBgUEyNi482A6oPKnoJUQQTe9gUAwClnfbSwae2okKj5bzC7Gg17MqMhnjU4cWsFGUhH
z3HWcZpDw/x/YHJ0EsdLXqSIxlVmaXyX6gfKR+Zv3cYDj/wmWt9jTLdpQQKNIkFSLUflg/Re8IFd
2sEt7HIgh8LzPOIBZTLVeTM0CMgevngt7xXArcUjPEEjfqgM/0+AGxMCeeLiQXDAWb1B+BhR8onq
oN6Qyi71i08oOfrllP9lUyohCD6wlaaTnKpcrhsNtxnn6MPDi9M0/eL4UGLkQB6aquNdvug5/bWj
mc1PUfbRJjmakumD+GFn6swlKWICvnD0G1Kep7Pwo7tNy9708EjdbHu1muDyKbwPLjqnso9lGs8u
2Osyr96+UOKYUPiT157Ssed9OzuxahRMSNxo0WtF2M6IVPcJ1RZT10KNSm+/hDEhkSDAnhGrFerF
e8HELXfems/Ff2wo2VoHkM00o2Z5x+/4wTE5IgyEDliGKNVGw8xoZ+QzosNgM6wj5/5xOworid4b
Tly0pRELssSEwoXA/wlXuxnwUUGN29P1NV62Qh6UdUu+SrpJTG3fCffJ3d7CV+ZeGbZZo4Rvpjbr
PZeufGRrSjqUi7puulHeIBnk8IB9ZHbmKdgNnOXQaFbCkVVb+6Q8zC3X7NT81GgF8rOoxfrlVWcl
L1WQrU3t6KAR3S6g/kuj427eiCvCXbrxd698RaBPmoX1xWTRIQyEiXuyn/YDnRWvRBxSRA4pk49Q
+6sK43grmygJf5+/WvK1QehtTzLQbUxrcuQ6O7kjPjoNZDioZtARr+jHmbqKMrOuTVhOGeyMw0gs
E8AKlb1cM7LYujuCfRzE5cAf/z25V9qk2ZS2dpEdY8S+Kg0Jr0Mzkz8El/7NhSjQx6YZUL0yRTHX
4Km6Zud6iDS4NymP4qW898NVW1/PpvMS++/Qz5lKlqN27knLZhevj1JYDo7tJeA+N8DWcUf69yLx
cCX7p+UTkPNHWIkC2pHBxSW1d2PbOwX2Y/+bej0LCRGhxkUmn7cMSbz9hcXHaqIB/IAdb6NtQ+mb
axLJDumd7qya3llaTbkY1ap46dS0Y8UuMrXFavrwicy3/Go7qpQblMW69AB3v8qCSySm5E5t7bzP
Au0R4NOcy3YvQA79c3lNCCzkJHYAdAuEwz1QD4TLakGx2nBmUfd2XIgQYGcq/aVX0nmy9Jm2Tp/Z
/+YH80Nf80WWNU19LiZRodyKeqpKbPErmVbGBb0Aly8xCIiK8n8Qy1nHRGSFIppgpzIKEon1NDRr
1z6SIAYgTSs+wsgxEw9FioqL/Iv9byvOZKlt0lw75Fv2L1h7ul1MJ3otf3uxC3N2brmQAmivXlgj
oEH67JxJkjOp5XyZ/9C1rbCt2tQ52CiEcULEhPaMH3xSWlPrkMqGbos/omZvMb74trlfVJVqnQDr
opiA53Sw9ncRA7X0sQBJp2zjIgIuMdKkG5sct76TCxEou69jhDxZ2C4gsEyM9TCAgnaD8Z5KwQmC
uI8k1VbmtqZDRrWyb4kA7LiaVo9J9UlQS2R3pi5ItEvLgtIkRSJ3TiCtj/gUbGvQ5qWY0qv+mTif
R/q44QHLVmbTAZKlDmDEHtkhGib/GuvQbfy4zlnoVruOKNTVyWqKjbDUWSHtHzs9DVvLlkWyvc2m
WztYzx4JO5X5jvMTG5W0lI+hV+rQW9CVt7TDe/LyLsbCto5iMDhrZQIpXQ5fwdO5WNv5eb6fKTGR
WvRFDAm9L74MErdlgZ3p1Liu9/mRaXscxJOYUT66MBBiwEzcGC33Talhg9wlFcomasQRmX1vdEpf
tLZCsxLEUmxcEp4OTFUZQ4GjSuBRamdZmvVCC2uMW5BSPA11/M7n4BIy4fYSTwKbG2jiDZeNyKBo
9QkXJ3ivxysUlGNnIm94BWv86tAE3NL+7tOINWnpyyVwPDNUcbi64BFbcA56k0bCmRQEhmfZG/fg
MbPrEk0cNsMZPl4QUIiJB/S9tbMa0uYRtUqL16HjoU1A6yUlwRyZ1Z/ZFVdpqViLzU8af2sGSmGc
hZxl8ZAFlQ9Wlnn11LWJBx0ySqD8qzc9L3pHskyL5yIBG0BQa9IbSPsYpCekjvsvcpznfa4X9Jts
G5u3NkOE6HomIxbEzHxIn5pdcWxPiIyyFsGMfiEZ/jaLqj7+SI0c+ZlUArVjNcMCWBGBJw3ClqC/
mh2r1Zs+kEimXjtcQz1AGsXBT+okiiWPQfEh2/L91tbeHeH6NDQwn17VwVGD9yJAbu6oks4yiUdd
q7+5FCKHG15yQm7z2hNX4K5CprK/+YFYrQKrxSEvpT3emOgCj3AuSl6MH/a5QcOHpttD/cpYWtb1
JI3PHgOlllMPgITtLnobKJlQYwMyRPv2vD/1IJbapQnWqlA0yER/+p8Micz3WsgLZDT1YtNyPjrL
cV9wjEvCwE0au3ctS7hth9i7dUDwJcUS/a3t96+MJoy61OuMuYREs0Mg4OCMwGjRe1WjchHZcP0+
EJhOova7PRPbWZVUYO6Va4KkKtSMOWiL7vD/eJ+Fn98zXIfd2s+vOWgC4QpL2qO1OLPp1O/MbaIb
C52al8LrWcMy39GJzn0HsOlni7BHC2cuBhRU7sHqblUOkJwuG+U7+crPJ9KQRQ5K9XhJESfEWVXd
+m2yvGsurUP1K3egQgQyQr/mxoIUwZaMb9ZINKOMdUrniMEvQhSROtOen7f3XuHhzgcCSLzruRqV
qKbjDrBJV3V+8VIYXpkGqi8za2HVPRVD4Kgfyy+74yizZRz6+zcP2ufrL9pI1QHHe9+XWpnH/YMt
eTEiuNRNc7OB0LMlEfjPFbcadxtp85z/68f2W4lWyg7BWWrJwOw8e9zpDA8aGlLfynm+In+6LZ8Z
P3FlShEPSWZJFMlIIRwHW8XIJcq3bqViwm8OcvLkbg9+68kiFQor6UtM/8id3ZBJQe+jOrp9t63u
nFe1JKqQ75bVMmHLybglvk/sloVaS1UKLNYlAMUQxTGMuF0A3lZE13nK7TDycg893Z+vLHl4Uvag
vG+/i9VcI3/swdK5L3gtCfnrOaPaQ72KFpPxY/X9biQk3uaw17DFPUTO0mrkD3ULPTA6AbecU+V1
sBHkpV+MIGnim1IUKTmkyazJVXneyqS8FsyWjHpz3eme5Uf4gHuDGO3zNVqW7/gvmtXGnc5idA1i
eMI4CfS8dp2AabYAuqTHO6B9/nZQsvU2bjOJOw2kodPjpPVwyLipYnxTW0X5yRbEHKhvH1Qsb65s
K3b53WCTH/JlOS10e9mWUr1MLXICnMJ2Ps3ju3B8A2Kp3QU7piVmiDyj+WEkwP2ygHJkLyeXPFnV
H+Msw27CaHp+cJpkbyzVXbGfEp5/R/IBkvRoryDclGhbs0tyR/U6idqz30o+XTCrmQAL8rnfkMLi
KHEahvr+nOvq60KnpmTW1C1z83NKe3DNIHl8ghDo6FUrHGXgZwo5C1SaGQbWjUGa7FjE/E6y+ng3
1QFjaeHEsNCe5fO+ZrIBORVfQT9uFDT2E468v/5tkBLWhT+CGbcWKn6QKWbymonh4vFMvSB7ZYQU
FfLeEdb+zvSoFVyRCs1atPsAckRA4V0li8KWFq61ur2Hxwt3v4gyd31gzhKckSAZxAriiY20ubQm
s+QnoVAo6vj8gbsbz+OlJo8DwEbv4LQsUJSWduNR6jY6zfwnmUpbi24iR45uaII+6YQDMSoVDpq2
il2O93kdAiaV0U0tRIJ+oTr8LYhS6703aU2TlVsbnFBYAnFrC1S7sh0gynDXg7LKxFqc08aOmOGl
5umqnLNX9ZoANyiJlvSNO5mZfzcvksNZTvPFfpKVvQ6ndlLWi1LsTzqCbWIILtDZAeLEUhYoM9n5
4iUM9upReTDFjEcVVaZm1CFTGyjd/GUZF18vsHcQMVVgpGzHHEVfOLeivVXAsndgE6Bqy5CDnjTa
TIOzsiQrjUf2BnrpSELQfhKIqBIn40VEZ1MT50Rteh7Rvg7UDp4JgwCdgEMnxX40wS+FkO9iXMcs
Is/0qlf6HyhBDfMlhI4VtgjDd+34+/QYyTGUXif1KnLr5no4nDFrmd2Oi3pN07XxsQIQBf4KzVPu
HFifpEpeamwSiuEk0M2s2v3RMjPREKwIJLSH+Yg7yUjd2Pr5PpRh1L1HNpvqq8nKQnvzx0jvo0Op
bbx/CI4AiA839CHTJAYkh4TkMNpgHlROI8gDAyvyj3MgwyTdgcWeti+f3NS9Bs2t+oIwZGI5u+GS
2fx+lq9+LOI5mZoCoICbfh8OEfvNKI32Rk7KFSvCEZD6u3LF05rAomkl8ozD7qpWPy1OwR+rYhMG
6LM3k0K5Mvxg7urC06dFHTrVUTeDH7+xQyaBeR30GtP6ZQOKIql5YsftplRR0SWdGlC0B3Fu1Www
TSGwl9APYRwXdq/S0QM+3H/L2GPtVap2QoX659rnydIl2ha/uEvsEKvNKK6W12vTDnMolHp5e7Wx
D/OnZlk8caeP9ZrYexErs4y2BJr3UT5MxDe0G5tqQ57t0yqRcF3njjC1NEMs6T39J9vPVSEZBRUv
L3oswtPAUSeqtDPgC+DJbIFf67pVT1QGuHRmYPgJnPWdUWzz8q1+W7L0tYCXMh3HAeqs3/RkMb3X
rJUQjDfcnIfChFyiFniQOrxD3v9Th+lC3KLugrnSJ3JGva748+TYKaePnOh46BUtK+VE7AfL47tb
WkShR1WIuvy00yfZRB5Ad7GI3SHf/74y88PZhnQXbJOIPS7PiDAAX9BxruWH2/nd1ofdtAxNCU5u
vY4XconGktMz7mrJ+SYdS1BmStFOmWM8jTPd88oPJbCcqXTk7qLeDB0o65Hxq2S7Vm3KSkXCiwHs
i9KVaaVx+Q2W+vg8sxEEselFVsofvGkLlc25nMtScuNBhUzZD2mZ2lSlrH8gF9M7+8Yv5U0EizLv
xD3uZR+cRlt7iTf6OxdO31kg7LNMFwA9fcpR4ozckinA+xsK7UeTTzT6CNLIVMtowBpr1XGPxZnb
WC5uEJiTfw4Z/4Y/WccRdJ2pZ/NqbpXgZzMgjOi540vBQahLbcj4WVExrymqRVOWswB1pLg/Tqeg
ISzYYUr04prmxc7BI1t/kIsrmrc8dvTujcHMZYHOR1WRMkbmXTlPC5n6ImE/ca/1R0L2+3u1G1zi
2uWL+3Gn62SaiknWsDiX8vz1HdXzON6KRLIsu9krjS3T6scXYQrABqHCp8mAwWN7tpytiYS7PmVU
qoEyW+AgcZ2vm7W7XPnAy0aknwhqhCgwQduzQYMi9Kt28DaEzbLs4RLr6jDBbeiK81p0MBOHBiZr
woucrxH8TwbSq4CwpO9s31eYaH8WCAFv7pFspqagtFz9KgITWb4ZUnI7vyaUaHF+i4wBIvlObIad
JYKqePIS/OamKc8mpz7Br/q252ON1iVjVow4kmenWMrMLB45stCJA0bLh0RCGUYYF4nZ1R4VRtNg
HDuoXnaFaNwfro9EkwqZDvVVPLaPx7WlaXHU6n6sLegthBm5sBSq3nImsnt3p+JkJqzZ0G+STHqP
LEo4BEfOCai+X6VwFIB/CSciU9XdtUsQGf7JWqRodd9KI7LcjC5lk8K1tZMcEUgSwuBIOVhccIfT
TjNDDr5v9BhQJ3jxrl3Zu3BBC26Z8CXdNp6BfI8BJbXUqy4QPWEQyGL34JPzvKOTy/nK4Bl4g8sp
s9YgvgEuB3pzVSCcpASAUI2bF3ZEcTmRj3AGLTO308uRMfo9IyaUQUD0hv0OPb/QPLuyTuoqhu+z
j75qgMegb8SgXufD/zdVwiE8TbHCOOwlh4cpJyZDH7shdGXZh5qQIKhns7fND+cPoAn8TmSSutwp
a3CowukzattieWhEL7f4HmV0zYneLIpnDBO2yXhZXNuFYaPuJt/VC4OlywsCxZRkzByWqwTWRccn
lRWG1aHq7akTDIJlYz3Gr44poSQgFFErDdzRCfIV4bBsdbG+1Kpx/OEZbW3clVqj/KPxqgaddYfM
z4k9SxrUT661b5TaKT3SE3C01XIdVEfFqPoAnli0JpQy4zlj8/HH95H2UyRx8oUtimdbH4DOOhgu
XSE26ILaSNFxCD7twHB4bxGOKpLMvv2uKRNwvDi671Sk5wKNU6I6YCHbK7yvjKmC735A39bx//eQ
OXXJ9D+xzFq4nKFouKP3eFfOkh1tPRpJjzAOGjwA8I6bPT4ArjUNLBtGgPvuAc75OsVfjizIEW1C
2HiBTLq8rsBEwu3Pm2Jz2IoASklK7P3URJjP7V4PYVqEG8rIjGRiX1ZQQCKSZo7+rw6ZcJmU5m2Q
Ony3+y9Wy6KBxTx0yyYjEORmE68mztnS/Jo+LJ8z79pimCU/FOUpMsX42vwzl40Xnvgll5AS+8pB
2GU26X1diYj8GSvcsOOnNxHxBtRUVYQWFGIFq/TAmyinlW9YLmC0ISld0PPT6tFyZtxoj4xedtxB
CpsKpYOuVpnXswQ034hAHL+JmvBsflvCHgvWZZ2EJPEdr+mHXqhpW9huT0fzb3Wfnx5hBXDhCqy2
RZAxRRV3uEh4cE/+HHu2aNRMG+JhfLCfNG54wBNhrtkIJMq5QVqMtJ+mq79zfKuc+r8cO01z+cqP
M/I/4v4HTjorcn1KVLaxEHfTqbBdciulkmbzoWWTqCqMogqJ69TRYKAJqmiibbfCDvzos0IYWz7q
+pZ1z908a4hxjzGMVelC46q558S3AyjrFoNREOF054/FRVGstyHIzq2yuP/3DoahAa39uWBUf4P6
DpBfwYNiQ4Zi+A63corOJFUV+18+ZvaHs1chwHtnv4Yt03V3LkZsLDRa+IIzYIFcIjyWOxKHIib2
1Zl/kABexhFDYK3n+p1L1LpcWpPyJ6XMbd0lS90VGQgk+hoxwVdaQqw2HszyJ96IKJw/PiiMhMxS
8XO9A4QY4+veE3nD7fpLgEjqm/m5fJETLa/oo2O0Z33ADy5gy1PYT4geZSKV1wNL0SdHzZrMlvUj
K+czwG27tRS/tpP8vf4WXr1qftmQFJg5t3kD2zrDcaxJqIgRHFHisZbJcyE/4I3XkiNIbcrwioEo
1YTkO89iZ8kJJv8Mk+7oHrOToOWqxpv9ktgVd5VvlMIp7a1RziJnc8ajcjfCHkNyqMYwuRkghnKM
CkA/B7uloN6RTUIg6NmTcP5sxJFofBM0S6YOcGNYNQA5oew9qxw39d0vTupIqc5cmWJ53xCgdEig
ZfVWGrON0huZVoCak7HJ71HZO30E2Yu7uqJtLM9YGdOqfebJqX/HSEwj2Q+1hhX+nQ6xJtoCUFjF
Az8UwGSFiqvrp91tg4zVBX+ECykPXThErNsMdleUxjWtp9dKQfTFZZ6WeMszRxdvBhHLs0l0oMkT
s8zZIvDJoLc1OuUSUjvbl+ALRcNK2p83Mt8geVvW6G5U/CWHBtdVTCJQAu3IrqfsG3Q/90bwXvki
o96OkstLyqENLG8lhcwHLS9nWaylqrVzU/ypZWSJ1IVHKq/UcZlpQT4s9E1ynpTfqFmyklw0EB4K
vpk4+GSHwbEpWHiz4TqIyBejpzgEw0h9j9H5
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw1n;
use gw1n.components.all;

entity FIFO_SC_HS_Top is
port(
  Data :  in std_logic_vector(7 downto 0);
  Clk :  in std_logic;
  WrEn :  in std_logic;
  RdEn :  in std_logic;
  Reset :  in std_logic;
  Q :  out std_logic_vector(7 downto 0);
  Empty :  out std_logic;
  Full :  out std_logic);
end FIFO_SC_HS_Top;
architecture beh of FIFO_SC_HS_Top is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
  signal NN_0 : std_logic;
component \~fifo_sc_hs.FIFO_SC_HS_Top\
port(
  Clk: in std_logic;
  Reset: in std_logic;
  GND_0: in std_logic;
  VCC_0: in std_logic;
  WrEn: in std_logic;
  RdEn: in std_logic;
  Data : in std_logic_vector(7 downto 0);
  Full: out std_logic;
  Empty: out std_logic;
  Q : out std_logic_vector(7 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
fifo_sc_hs_inst: \~fifo_sc_hs.FIFO_SC_HS_Top\
port map(
  Clk => Clk,
  Reset => Reset,
  GND_0 => GND_0,
  VCC_0 => VCC_0,
  WrEn => WrEn,
  RdEn => RdEn,
  Data(7 downto 0) => Data(7 downto 0),
  Full => NN_0,
  Empty => NN,
  Q(7 downto 0) => Q(7 downto 0));
  Empty <= NN;
  Full <= NN_0;
end beh;
