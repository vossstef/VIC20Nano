--
--Written by GowinSynthesis
--Tool Version "V1.9.10 (64-bit)"
--Wed Aug 14 23:35:56 2024

--Source file index table:
--file0 "\C:/Gowin/Gowin_V1.9.10_x64/IDE/ipcore/PSRAM_HS/data/PSRAM_TOP.v"
--file1 "\C:/Gowin/Gowin_V1.9.10_x64/IDE/ipcore/PSRAM_HS/data/psram_code.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
FRM6sprtAK8hxgIDP2bqcIqgWPzLdgykXAIciRyDWgWLRTXYyMzJifs5djxRqnqA1KG8JEw70f9F
xx8XeZpR4BbA3VqdWJZtx/uAL7VDRIGtxyH6x48j9egX8Uia+WvVlSqFxqUbAq3qtt/1SIHCy4an
3GgAMMwsjTNws79PnLiFE/kc3YO0t6lyed3PmKOibprE/XbF07oZEFEsF5sLR3l3DMBTNvYPVWY+
2t5th0BH3Mnvo0C5mPvApUq4pVVDuOsTM4iNMgj/xWCiU3KHgyTrGsdWr/VHUAuoiR9cY6BUY/G9
nhyjAKiMjef+nZ8acH6xey4NZwO6Mwa+jjVm6g==

`protect encoding=(enctype="base64", line_length=76, bytes=310448)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
+jYcTQE/5IfaX8Nzvv1O4JqL4AOHlFXWTGFphebFVHZKjF51s27yHoDevk65iGcGmPvPVP09q3Eo
+BNirDQhal6EDBeaOEWRAE+lFRvhOe1I4AA3yfN2Z10jRMXHrDuSJnyV/6cQgt7uvZyhUsi3WA9l
kU7+DJoHL2d39yrNh1C06iAVvS6WBsOgfI/zklkjb61X5eD09i52kMM+/IS+rovMsDHGgdW7LeJM
vkQN7z5PqSSfG9hq9yjls3BSw7f65iMLhbs+eSvX0e6mxC+Oq3RsNkfGEPcKEWgO6VIDP2ghZi9f
fpMiTAFiBWYI32x00iFukr2lllMo6TFCZme6mn9ye5PLnOKgwWCklTJ/MrKQGo5TouNU2H8YUCJW
faxzNzpVE/IlD9ogZoaEfWifw7RGbpb8+PAFWWUbqvxb4ngzcCRbjEKM81m9rVFZssjikHN1uLZO
y6IxwhfJ0e9w6V37fS7ExzWnKiePFI7CTkSXsZM/nbQjxaBlFv/Fm4qSAGjR8cbAcatai0s74UFr
LDGLjUjZocf7xNolNHpzx7ECO99YCcpVPv1itSy28ld+R5L2U7gJOED6FC8gHCP1CMFCSoCvwJPo
BjLI5GG7VFRPgL/XgWX6z5qsCvcsworD/F+1nreG5rTdKYo0IEtgCLDU4ng/ZfCPmE0sEcy6l72/
NSLfG8Ev5c+BCyxRVZoRXDfomGe1HDb4YS6fE2REgM2FUkFHlcHX9RhBlH3WBcnWnoaKPo1I8GhO
JlVQkOinXReYSqTYyu9/yJaSjWqFQNzFi2PHGmlhSbmWgX1x1t1GJ3kX9km7uYuDbzCuNUZg9Ggf
vpywPGygkJvLFMyj9pST31ktN+fX9viC4SlgEGVtAJ0fdziaGrlyWtx9KeVLvmuU9naUzoERTVMh
v1rDEZwakV44noDbNsfG1qcb0g6iMmYW3FzZe5LJk8fWTiw0lPynPVzovXxGTuIxdGze4O2+ZTwg
gH8r+204kLCZbTSRjrLaPqFyf98jtl64OMCVT/oRW6YKSDPlNLg92mnu0buEHLE0cOB51Qc9IY8c
Mbz4hELAZ1HK6UOhiNMd3iJSUITcXQ7l0eW37ckfe84B/GiHxdDoYg5QxgN2JTmMpUgJi9GCkXJg
VtLzAWI6/QDMLEJbm1/NeoydJu/XfOv97KjRMuMrP4F+BJwfGSAWIinFp7hW0EThGT/J0Tt5oYE7
erGwQ5syBSpn7YyUUZh2qBjEclpUh92RqJfe66Ct+RWLfrwtWzq2ypW+JpkBKCWuaHSKv19QKMWE
nLfFlPOj6zDReu+4XzGnXHqlOTTl4/VF1xSqvF1hsKJpuv7cglGA4UQpus5Pif5gXXiJfCp9kw3j
wQ44FSQBzmsmebyN2uH6h9EKi44V5jbf29XCksACRwuLQUR0wi1img8ZNEVBZhzzEkAndsOhcUza
+rYjxxpq0Rswm3FDclDGzwB0OoPErdrgjmgvtiyi/2OEfLlYQKAtHtuMfOKgaiFDlvme9gO66y56
6ZVtBYuxq0VgHKamIiOFbNOSvGhWZaIKclI4q7zswDwVlA1tFXwJ+kg3xzIbzxFyh/4NfOEHQUwj
aONCZ50ZP+PKt8oe3Iok+oAp8YZhBF5Gg/FHT3PSRpCNC/5angcBxuVo0eM8JCQ9mdxW9cvXzGbU
NGdJOzGjwqv9/R6Q+auCBfWBhruahKTLs+D3T3aIY6vjtIb/yZWorM8p5R1kkCs+4lx3yBQnXcUM
0FJjOA2lusHEhvYp69IP0UEEcqGA3bJeIZsZudSB5nt1GbKPhkBXZQAe6E2Zc+DDmTI6bx91h012
3fZpKewQtUVzjEE+K07vnf/cegexz4xKb1M0YkFSYHQjTABgCNgfBHndBGM8Yg8cVWfZWfP6hwpG
i+vbM2N9gMn2hRExC2hxRPmQnfNhyD6dZKQFF0XMRQQiDAuOqWUqjn5LPvG6/y29W5MP01yP5kGe
3UXYlh28OXX80pBgwDwo3SbjP8NG5j7E7yTqWzan3bcbIT75vy+TNKdo50X82pCDzccUNRyhmKyw
tH3qQgn32K3JUHGM8AsoEGZmwB61dpCvhmtIe0t6xqP6hmdnA44MQM0+NUD07iPVizD2IWbVLXdu
k6HHH9Nx7m9dcUjZTT5YqDzRRxNcg7gXZWOSAOHpPsi/npZbhUkgKhrVwNsx+XmrZUP8FR2l6uss
EwmrLSrvTXYDCZmNuSSUgc3kQNdpZ49gP2ZfDvdbWr0PMZ30ttX511EN8GDHj5/0xVlmF/iLVd88
ljbsczo0vHHxDASAkzUWvCkbRueV+0d3n6D2lfwdLwjwpmPTcJvMfv3Nn2v8dL46Or5I0+/hYom9
eLs5GNoglwFNHg4lty4l7QG1NA5boaVvMLV6uL7tJT0bg+CAcDdgZj7zIq+EuqaFsMZnaX5ksMgQ
TTJZFNjptBz5sehxPWkz7UuBv9lp6UpOOUhHGdgpXS83CTHDiNqPMhk9cPSdshez1YHgYblCSL46
/Wfap4PzpTim40tC69mHn5NHIgwR+CS32bHBqbLs5iDUcRRWpexovTcMtSrviSnI80KGob5U+Hk9
BN3G13K0LAwimhKbQ7VVTF2vgsURrP2QISoPAy37/UI+pX3jcC7t3n48d7IgwUY/LVh5dkqkwv71
Uz0rrg51UuBoHbpPAt6dViy1kjp2/kkSGzVe9R7Vza1rvOyoKICFpABjUOq0HJP2ELFW5znzUXFt
z/fWhWH7x3XoCbDm+UWaUEQfgOt2If9AEcZLLmPepuDW/b85bIVAQ0vEl/l5+2zP1zQAUBFGs6Tq
WE8Q9+O2LgqFTBnQt+s2Bb8vXjvDddJa3etyqYUSlMwXkgCdyy/ln055hTGf/tFyobEh2/Qpdjv3
aU6VMdLUHFBwW6+nC9TORDGFD039SHhrCpmC4gmJUM2M7w6tmr66E97UCLTonNulpM6JqhtDpQiZ
2X2xVsBnlS+DV808Pw1xmM1lRuSRm1MnVzxrzr8QeiQZpEUIxzEx5MeT7dnX4v1/oFjzNOuF0Wjd
Szzkp6ghpjfAhGZ+l91jPXZYv+q+NBz+DePkHej9T1EY06wF4A6GrsdmJBbtrC31nmvE8lrGY1+r
FGvMxAUrzcQvpUn+4TdJYp7y5Q2skupSgn5C4ICPucf2L72pOj7snLu3hwU0WYMCr5ria7m7jo1l
4LgndvCAl6/UnhaWzwQtBH2dIi1h7nFgV2rAJvZXs1simQu+nsGynPODoKobDMHX2FWndYpkK5H6
wPZlZT1x0HCBlL0nQnHaptw9d/VAMYRJsPXkrnoaA0+aT2NeybgUApEGg7m62m8M0MQWd25S/Okq
e9xi5f4zWdtSBYOLLbkWU8xIN5jDC3QUvPr876fqSXAHe1P8QWW8HmMDhNj2EVcO0PXv60RIL8ko
ReN0CNLFEr7fJBiZ6fFLJbNyoJXOWqcg8bnn1GHrCtf+ZCEN6HVyKxdklnHIF4n0xfZr9JWPrtX/
sDOIEM128iKLooSHUNvO5Uyiefw7V60YkyWW7bsyFt3ZVpvP0g9Fl4KqfpVxyWZm0D5FbT3pzH/x
4OTfyrthBH2qvwozQTIP56UixO7muU6oKq12HQpbJvlipnrqB6VXzKDdCBe0mR8HgvxtwvnvjlQi
GE45WnkEyPONL9gG7eXx719NA7lCZue9jo4wCB+75zEaZuw1kndl+pLMHfpxSivVN9mElJPr3ONO
vj+SoBxfSoZ4nlPFWZNnP5RzTG3zjBJfrMvJM3E2b5IFkDtDtu6dG7OM/K9xKnRMpGtK8mfZsPpH
v77sBRyfrd8HMRNhBZOogkdcNBoFsO+DD+/mj6zrODTceeR0cUJWtqJNCslTZvgfXeLQeWNhxCuT
RbvBx44BSiUhNt62ueNCDtzIPic9+5EIUrRVHTJo9ZU7j+No/WxzoxrynBeUWr/dU+skgsdUpBV5
WydnXN48w7Vl3t362zR/fdKZTgHLoKXQP+TqECy8bx+yQd33KSyJk/JzsVnuCqi9LfHRCNfKB0W3
n32hQNjMgn3XhEK20DO/i3ZnE9+5A8mezLjtr2OT2Wn/iW9Daud/fsoH8iTI2FJLmq4aLlFMBglL
rnG5Cdo29WJztAjp9ukmVtr6N0KcvMci8Hj3lTszwtSBlbAnuL/cv34sMm29VSJkPsPT1Rr7wdhl
foED+J+70PGjTFPNLkHfufU1IjR1wohwTri/2KHa4yZki148Z7N+qgaaSRq3YaBwHazJum/eTmhB
rD4OE3DD/zsNKmlXDg3GfAb/7QE/RdvPECw2MG7be0WAyrN0j2fV0anM0I7waOSYWIkm5hTMyr3M
MeY3aR24Lu+2+S6o2nPH4UgVmth4R9ENGp5e9/1mrVzr4fmZ/p+Xsoz/bPXUDa0cEv481Dym6TdU
ugaakzAjTcivxP9ObKSCjqcj+F3/EVm+DRv2FFHzpOHoa5sMu3F+acPaQbs2jIJC+UQI2aoCrxEx
j1gZCoB7auCVObkCmDnKXbc2nrB/1ArO8R7RgOUGWpfqRQvIK5y+701KpPY/9Cuzo/qQ2qV3Xkp1
7Wse+LJbpveZJGzCgRRpRv6NCk3v5BJlFaCb+TiVUOTxYoFzw71DLXQ4CK/zPEpTJp6RNJFqJJSS
gJR7l4149/vs3tFHwL/PmMyrjUkisHMHRcQYlfyZh2XKc8em6Ol9z4qEkJQRjp/K1pCQaMbwnNeb
Q8E81R+IQh8lNq/XmyYvkhNxpJ075fSWbrPhjEltJAZBkOFPYC0OnUMpGhg/fuWP1i0LyISi2EXN
koKPqws+pMmKE6Bj+oxM7H3wURGhoiaeH/PPJoZsEHKCitemrfiZm1Sop3GEmbLaA+xEAdOyTyS2
sXPAa1Pyk5+ibUr4GK56DNM4nROMf4yEkR/aEuoDWKD1d5QA/XyYQSKQr6FmtYYtaeyon0CD6Yp9
76I08iqRbLsjzlMJQRpHKc87X9qyaKs38xXiD4fUpF0LF9/EGCp/8YhqEr7UWjMG5gDI8GNoo5at
D3sj3aHZ745kIw90/gVxry+LiLyrymluQRgh5sX7zYbm9ML3qU1/5mYGLN/sw02uLbTjQk0iuhkz
x6ovNDsqy38eLqJRxlRt9gRtBU6iXw+zjh2U5l72ekcvjn5EFa/f92P6Bk48t23VIyopenSs3fyP
g7ixCrd8HeAUT4NtF9U/G6zKgaa6fIyPwApP+0k6b2YxNqfzyaJnU/ERSFG1GIgGTuTNUZXBSX5w
boIAuKsg2oJ+HtLPu4yQ1gf81L417sbSrSTLFK+LEZG2Vgc+QZrlA3CsyhP3lYSiT0gCyHVnivG+
kAxcwmkbznrnHCiO+Tco5i6CzrHyUWF1PWcZS720bFle2Pq61V88JraYVs5vN4WlTggQXZlfznlb
IIl9Hzv054Df+K5wcVfwfkV9AcpDwKB+nnDj3C7JeWR0eVVxStuVsyqnuhwYR4gv3ops+cY9lyR0
z66G/XhpHPakBK/RTb8M6G6uunM82ZYbUTlc9vbzYGT1Z1WKin1Rw/bk+qAQBhBaG4SUpW2YbuD+
9FtlCqMcZ2HdAZFrvCZGjenw5ouHiCc2lGky6OG+/K9NVmSN3xx3dlF5xWMHkBfRfhxQlpySVd33
1sDCR+spVl5MuDhwm/1F7WkwYl8d5ilYE9A/BReritz2wPjwawJEBqps4NT3xfjBMcIRQitXWsdA
h/TnKhM1vYNeR6sXpk4DesPCH/iDJ7/pe130wjyMGJZ98FHMUYPy6MGzaD443OekpjT4gai4lCKy
tmKWGOM5LAewuvigyK7OuH5Msf2OQAuWcJXSA3dExAbmajXPojXWzl2Rb6ArUO+zNMDNBsEIKbZr
7GKmsoCKb+A60TMw23psrqkTlLHilHJovRg4JJS0xH0Io1qdmhikP89vvTKQDBzoFW9TsDoOnZna
V5UsxYu2rR40KzRn36wL5DSzzn411FXnq4Aib/F6RlXxtK5+KRwpMPlzbUQH26OuN9IjqLa14+o9
XEDQroSUpT/oco7XYS6GmIqznRF653xQxR1R8J+GiMLsu4yv7IWInZKtZYNv3uuCCMztKEY3LHgE
rmqMrPAui9W0VB2kb4aST7LRinpFu6PPs0kzj9/LxlWmop60QDzM//oBqdhtM04R1WbcbMM/qvrd
uReCdHQ3ey73hA97PgWf5hVXCRMr0fBb4ise4fIfGBHQTA8vp/1+fCssyLk+TqH9FNhEfJr9v73i
mez5HiUdmndzNBOh1HO+VD45zH01isel5tiVKL1hrQjo2OcvFsoawSiKXtbE+Zd7bE86EJ6PcEXI
mBiIVjjCcavO9Sw3wmryocrmumBPbnp6iy2+hZ9elz1v8/3LAOIBmiJHLnx58QyJRiAxgKh3tC4c
d+y/Mq+A0td1I7yk7N25eTzd9MefwhRoCIvU43Wbmz43yeBQUy7RJ7x8+SE2zGy6AmkBF2qNX3K5
fX8CsMZ/JbezXUV04Up/gbcoOvZG1ju7AbQKWrAow38QKdNF1WFajU/zDs12etd3ARKL0VQr8+MF
Jq32xPLwDDfOYi7wB5J1dMLz9kPdbkCtqoriaGJLV2MX5Npwg8AgwBdg3WPVGCHhe7mLjGV5pp2J
MtCGhNbcX1CLTKC7uGc6sExSBFA64LCgjJrie2B9y0AlPTfIkUTITUmTg4dG+mxuiPV0e2eWiLfS
V0MneqrdB0lduRaZRU8eDxuKhjvN1ZMH78nqUBb5rfjQrlctHIh1MoFiQxcTbYGdN3og5z5UaIjg
yVCfz8DLMcthdhmTovK3H5rwHJMqJXKfHLMsz+bz7bipd6+H6nsBkOA9jQlTPCQL4X1VK2nFgTFb
UY4xeJM11zXtbwk0evkBujNTvzeFtwkJ+u1FypRo3YWz0dr7Dq5pUc1+AdtBqBko5b5lFb70fCor
0DDLR09WoQ0e1mr6WtWjq4vMPamfc9QqUhM/v9I4VD+ZAVv7jw6pV2Uc5ZXKTcMd2KEYYy92C+/J
rmzjeQuTa972tWe6hcriWvYzAMoVNfmZZpA70ERlClje3N4Iih/JAdif53wjppG1GOWACs161Fwf
rK9p9QnUCYHpiL1K/LN/Y8PBKssPO2t5UxNzgf2+J03oJdmY5q44Gwx1Vb9zbKmnO587d1xqfXwX
ewQu6vldZXRdABvHmC+q9k72v8mZRF7mO9OTApo7ZO2Vz+20kZ9+eq5uMGozHhUdK0/WwCUBkj54
cQYC5fttbYMs2mTyJfihbyW/JdPKPdBk2cBpY2hggW7JJhEDZdWLl8yj1UffXCJvBIbVMVaxUSUs
No9b83OTRj7x8febKAsnNpRnPYBcmcQSdvLisI3E5s4gCTocYJwCAaLgnAnkgOcOAonmbo6vzAy2
GEckwgTVy0WgV2hdKqYiNscbLYWJgF92X6vqF/HvvjxX8NkXseTd85hCclr9p9XBG0NW0i/dePWn
iJWNDKIKa1N2nPjrlFmjUepc1LJfFSdNmD3D4Ac6HxbxjDNotxRAZokXOtU6VEEG7L/RLNPmDa7o
ZpfCW+uwrtAfPE5sSpivyu8PSPoNreWFaSvLmYXLXmafStypwIGWoo41njFs4iGYXOGz/IC/TuLz
wkrBopzMI3dAY9am7XmyUiWXnn6Z9DPFYhxd1jytGfDwC7CpubvkBTDL0xZTBJx7pZD6d8B12s7G
psu+IMeImPi6S51wdYxlrv+rHBIOtb4Gbuhfhm4AAE/6ANlAd67ebiZzlJsfJRNalxaZoTY3KMoG
5InwQGRCkR/qbGFwh+N477pD9DCcWtkv0cS7FvWUyW0F7bKV5iGjcqPgN2ctFbB9dRiKWM8pIjvH
VwkBJrNNjvJpzAfT1VXx8TwcoHkvYQjeihjvONAEF4HrMoYnKoeUsauETJNsYfigsjpwYx0x/5t7
90yyklEVVmSEvpznnigjTLqGMDn7gjgc+rA0/+ahiqbFwzJVAnHmdmWqhIwPFh7WqUsWVdj96+Ld
fBUiqI7YpoAlveMvTtCBV5EcNzRCPxLLT5DCNHSnVRHRLKSyWFaa+U7x3rWF6Lk8yK0YDizoWDPU
eEnLQwNgbL/OjECBgLSz29zIKwyZbdips2QEAJxJ9sZ32jAhMGdnkpsXaD163A8Q6wDOfqdcY9LL
SFMP6Gpm7cHUridCq47P3wzXYUdL15ppqkJ7B+4ZXVxMeys0Kb2oyQwJVQsunj/oYNqgaer4sfV3
B05eNi5YCPpufR/Ynmh/Fg9h+4czndJqjyBSnKO3hf2vcCEbO6iZ0T/88KaaFTQNK7Z9TwTUXNbz
N6zgAPOHqZImeobqvB1h5yKFm95/w1Rnoi8+I5QHQudWwNIUeE/wRg71U7/QAgNaFf6BbUiE7w55
Vt3vIsak/zYtbZW995cdrd1iyK3zbvUAgVeZEn8tlDuSUGKuBc+eEPWtMltn5sK0ABeUrxXpXWdz
OPxIvKow8vmeXV+aw1FFQIUSpBOOE7/HGxHzZy4vwpqvnKFWHADvNdrtkfgnXE7LHEts/bBKksPa
vNdGzuRt5wuRwwZxASIQdr0S1SIOKBz+OtywKozij82tWX3UPz0Z+vZTIFhD3ZjR0roLyPVBd9bc
qu62RKNqkIucktmAvj2wMEnxrzwPwoTj9bhC3kjJU6MWyhNdndpI9V6Vu7AVSL0+R1IzS9xlhqAN
oXH2Fg0pn+Qmq9d8/sHpyuX+X6dt+B6bNhr/TyCdJvl8Y+Cc16lWu6nE4DDOg1Oa/gmAviCDXRM/
Fkv2DIiCyCNfkA/zOjYAmligjTrdl2bRQUIvhX0GdPLf9a0QjK+2rT2KA0kMb5Ub3HDD2/2s9ljE
VItA0PCzUGzuk2wFsysFnSWkqlk6J1Wd4rRPKO8II84H1T77cA8NLshI3aO8va0Pz6srtj8g2Vrq
qCVarmFHmKzXWRoeM3uXtiTxZamsp8f6foV6JxrITHysTGmFoFs8lmSJft8y8bPaxzJGIzu5aAZN
MlTfMF7bjAgwNkz9xWQ+zUW3P/TntyypJLRuYK7x7XMS7N5Jb8fm2d9W4W5dCtuHD727Q2esw15L
FgIZceiDuFp386yI26+xgYA4ooFscWtJQdMq/yLcCcMgdOFSRDaxl1e6uN7oX6NcWLcONevymVHW
2jeU7vXIkeINJ7uS3xjqm0PeTR+60DflT9z2YsDxz1vUYWHjT/NOJWMgQNAOCsPxNfByh67VyocK
U6qfwTePokhVNq5qjn/1cITPkIDaN6f7BHZsHsmtLUHayYoLGF631aVxwql1CUqUfa94gD64qpu/
i57fWt/jltBvKz8z/Kro7tL3gWK8N4ZU09odRnPNTjoSVagoemVsC8GtnRGlaTExAyK6jnfR2oMV
QhtK7yWVAC9xsTMS8uUBTE4VHTKi922gdk9TwUe+4Zyc7yR7szMu7HgeeXDE7DENqGl5sL1+bubd
z6mA0+YlnzrwH08vJiT3cBzt/zDE4U3CzS4Ew69X6y46f6XcrtGJHf+kzppXGxJSeQv1UEkF8CX2
F0crO3sOKtBkU5ilRvaqYSlNJlKCW5K08zEOJZjsMTSf/gpP8MmroVGzq2M/8FJLzd2Qch+rUPER
ax/df/4YAVCIcclBPiFeySfIhr69QPZYFx3XzTUDGL/X011QTxO+C8KKNkG33YcuOUZ4UXcAmT2F
lCcxzmDR85jNoAVJXsv+0OWHeUX9mNo5tLdrzgos5ao9SY/OJ0ZzSRcaM7ZbPXaSiu7AUOBA43bN
CY+SUfYVnzEEFe0wQU0FGFotDP+86EFtFCr/ccFAb3b6M7HYyA2Ge+A70sLlTKUpPLZU+G69soVs
0cwfib7gtSX4Eg2qbxQMUCHmVHUwCkBmv8EFTGVfnxEl9s29J68T2PvSNchiAb3hjj64a5B651pr
WBrATVpnCeUbQ+V+yeOnSj8PgFngYUCQ6NKLG0o70IaOqCoXR7oZEX3jdJDRcUOB4cUgjsjzakIP
0+beXZJ31Za3Hv8uXdUWgKdyql+6GrPCFv1/hRoS1ntVXLedhXkHKWoKZweDLUi9OLf0k/cJ94Sf
ywOK6DNHdqkj3cDjssfPvgKo3ktuVPGqIZlvhmcS3xwZZZbNe7Q3FqLDq5rcYbFSo9hbHdriotZH
cbwzRP9bNTLSLfamVBF6IOz0JoOJh/oB9RAHPrFx0y4zM84w8IPGtgKZEpWsR8OESs10bX95/ckW
mdXahKgs5HasGQmLvw9Qt4fMc7vx4DEOGbHy1/lKoKgAIIQUMfA/xqBWiN2Mtnz0h+LCY+Il8hEU
I8HtyB1SpCUyP1JfhFAe91JIG7cLBV5EO0sMtcQAzPzObMc0leGKsBo92oRbhrcRICEbkP7h9Myc
sTh4m5V4ypnRFNU6hsznufcdB3WJn1FaqBMdf/6s6+uai5DSsSjtQnZjGl6D8VFflZQ2v8EVdDv4
A4nTIJalmLnPFsc+yg9n0PY1Y5vy+gkzLRmHBv5Aq5TtMTUpS/QNEh7nPNml3blo27Uy7UFmtOxW
V1rpAHMCU6XPvigR7r1BDtY96JvTp3yxSzUoROe9U2/0KyLhOHNZVS+XhSrQK3/Dmw8xYWHJ17tx
lQSo+puWWtYSMDg5hx/twZlPnPaUO9zMzC9qj3Mi4B+jnQTd7xNxGutMSCysI7An0GIr6GGgwyRx
jzARSWE3MxY3ssem/jl+HIXs56t0NcTQ0S9DX80sHgPh72TbHcKXZUUmfHvUfFPPzowYorKQcX0F
TeIp0LmYjRseFbsbH5JqWCS+9FmBr9SongXmMdLcX6MEPCUkVhflynUprfKJRkg5iyUtBy014yuZ
xaFCgAUaPWz5dRZR3gi8xJzAHDWzmn1EnQitwsQ6vDRfzPTFWp1EHQkMNWT44YA/KR4l4uldQn5j
3Ka0LxISNKVg46oBaftHo2FwQ6OgjuTKPm5+F/BWyyAAdST8g0DWpAUXOTapBDqoDEfx3qCql7Yf
0229E/Nhd9OEoziG05M3N6ynZ1KfsBfiLLOTFkGXqNR9ZPvH5m9nQKdgSt7Emhh2sazq2EuMFCE4
hrYDgSIMjDhtHmu7SPqg2EtCVwtpUV7wwjMWWZdEhoTlqynUrReqsX/3vw2bN8qUC5U8ehfngjEE
JEfOJKMkDiIYpWrsXGZgpHTlPzQB5yh4m1KYMlnESt94WsfEKp1bQcpVlieD0JpMepRiHmxutrIn
wwB1Kt0ttzi0sa3KT6HR0SfgaQXq5dS8/y2LhctAzV1gxY+lmdHj3b451MwGhPXRtK6DUHbD/mSj
1S4v1bQNpD//qCDYUoIPG1U2fWUC5Km2/JZ9mRoeRcFt7MPBOH3QqsnTvF+3WKI8W/IyMFUwb7Ea
XaYEmdPPraQwjQjNyqWDB5ar6iq+FyumBt8wL90y7fKq3f7vpgciDc2kIdAaMu1RWdcJO6L5/cg1
hQO4gRcCIvuozwydYsGbsml/t23f5Ab3L3t8e3kONvXRKnsD35vey8e20Gb0qodeOJXyaU3qbR8B
xQbLtdAWagVb8jsq6EB7SyYtdDFxKnnzRVqVOhCYcpvcr8Fx/SSQzVBtQCuFpsFTD7/0CDvk9m+g
mTosBf0DG8P1UL6R6UmRfE/aur47HHpM1B3gGC6G1XWsI6m6/+08R05hCORpiO+QN8BmVOBF/jBm
RC3hosY5Yr81wOicab4H+gw90ngD2X5K0OOWCc0QDxbdZy/azycZYjO1KIA/jwSW0EwJUtQRDcWL
g/Ph9mDon8sW7jmXMkG4nCOwVhlz9l9fvubj5j3oPivAPWGAFcT1lfWz8Z4kplh6dIaGYAbPnB8t
HXYvqNO8iZ+CYlNGM6qMW4HV34zNxvTRHCG182JxJNT2mbBtKUw2GyWTXvThELXpKTFccm0jrvYQ
QWvFjHKKI3RpqQb4RS16kl1h/kMaRiwAw3ToSznTA1YQETPTzcyf/l3a1/RXkvy+Hgr4hd1d0BWh
ybXcZg/buoxagkcIdNv1T1m7XhZXI8UIximnms9QssmYSNVFwHeuBI7XtqJ/d6d2UzRjF62hyiAL
gRuzW+wY9jnvirFQDjFouqZyX6tJp4obITSyMVWOKDhj4pcr0JcEbyfi0EEhaHOkLWTJtQH7uGRR
WYp3NYPk9SWN7hhsq8I8pcDUyFeCPkzHtcj7gPkch+jGZBE9e+xhXb7CAB/DXLVIQ0m+IBY2mBWI
XwCjdo7jcX/RRim+Pcvtb5GB6Gl/gprvEpRxv55AiAfhRpLL+fbo+J6crSnPz24VoyXU6Gzbh6Qy
dWRyOBZY4YMgAqwsApewV+ZkQDjsBxxAuRXqk8T5M4i+6Jov1y5Baum3BA0iNDAR+RV7vrMtglcJ
qLdgbDTYDY2kYV1AiWRLnWyfiAfkAVI0eNMdG+FWOM2X9RqnU9VqR5BnzA3vTr++ShImD7a3hNyO
luVB++mIy72AcaPXoKuonfb6qhHSpkR82WyBnEpSD57368LFIHzXpZuK/uY1aIXpGHMnYQ2P3bLY
wo6BM+9u6H7xwxQh+8oyhOjeV0l/VbTMhJJDDJ9yretYCHOZQG4XsnmzP0Ba7pkix+FEPLaKgOCb
mqOnmcba5GD8FviTzn20cbGShm5BgrH18ExeFn7jga5IVcYrZubyrnoIwRbUrzWmUA/smspnQ17E
+/uchWNkcv2qdotyX7onHMmvazFy3/puEKyOuhfNdACUeWh3Vyw9Q78yRSG74nV2BZK/iBQgoLmG
o17efeVB6OoJVtygXq3Ht/JLKWEr8B2wpeQRIJjCPaezmQsL2YmwJCH8eDqZO5anpcCRm2lPT7dw
KMiCp9r1kW+BqIt3qJTBSwZ8NJen8Q50pgruhJpdqP1p4h7N/zPPq71gIEESDRDfGE+Uc/GYxSum
Ej7GGWnsMZU7F2QX2hp87H8dbiZeQuh4gooDjQSdj3E/V1EhqnAT2RfJgIfRikjTsbFfDfUDXsr4
cmmV5bmiIoWypBsDSd8ADwLor5CnR3h/9bMjLjXC4s6uhCDmu0Ej02dgmUzYU6nxNyJgF4S0/H/6
x0pKe6uYTi4kVQoEJnQv1EDp8QdsaH5xA8/bm4drlGg3y3CarbR7fTDUnxpNtQE7zXSEanBijNga
A+6JYi2e0eKZqoc7uOpirMLc3wWIOOImni5cLcl9gdNf9k6HMMapZM5zhhSwQmqHHkGULK6lstX/
mGYPPuaaOZ4gRk+jqNCfwtzlS3kfU/aKjXK96QG7CnNDxYYpSNY0fE2414WqKvDpOePFX0ZFKZh6
0U1UzqSeODPX1km1D1sfmzzlCUEWpAuF3gHn+lm3JlxLde4LJ2WhG7DdoAak+LDeb9zoO70hi7Me
CiMBxwQgbjqrCJHyp0pcplr7mwB9O4ZvXqPduqWlCly8vU6ZLvJgTf5fDFg1t1mfBPvrLhv6V7LI
wT4xXA0QzrLw9w/5LUWZYD38cIL4GE/Z+dgCAQju4ovWjjDthj3hSLxs3ltb0FrhbmAYFMp05QoN
+Y8POUhdVuAauAcsGF90NR/7TvRocf2WCI7Lxn2QJuqMhQzNjsXcM0bmA30hyQpZ9Bd0r7N4RtqY
6LKFCcRMuoxEOu/2dp5VJPM0qfpAmUI8/695Qt7mOC6CUz1/g74H3arg8bgRyJsMljcTyChYy1M+
dldeF6rwlt5A2fhkzAG2llUdY6unXyzaSBti9aKxL2Yq87DEb4ks6pG+bbZ8/xKGFa9PqRzJdCPE
9S4y9shSId/btZbo6JgcLaeeehRa7KEKnZUQXmjHAm86NBvLereIfUCeskpbTexHwi3s+gBxaNK/
QDJE/dEcmqM7HYhPDFJR+efPZjK5GNgATjTdtRKx4ylq08ZHaBVVf4+6wKfJaipsskT+cUeDeOyl
Y1VqIo70E8tEbfCG4I3i9TvSpJoo50I0aEM5gbGhVbV8py/IK3zYO6meZC2eyuwBvt41esTRyOCv
iQga+9DcOuuxZQ2BfmGasOZ7fAL4mpCwR0jr0Vqo38psCdHnFY+2yYGPmg7nBweVYtfkfAyc7B3d
4ju7PekqcjM+rbmvlDXk+v+zS2qzvU2LEHUmR+WpdYkSQLEJgGt5fhifwRBNwvNFXYHwGLFjW/EU
+49sDCjTb7s42Bcx0gJVq1I6IwDxZICJqb05SJ66SCqNw06tmPNFxoDIPEVFrbk7d8KNUnWjetsd
2FbbF2UOEPf9evk4kLv8srLyt07iYxcLirxAWt/tPVQltS0qfR617HUfQ6F6eVJwsb3d/600HAL9
T9svC6d+izY8ab29PTmBtdAj1nsHvy8ZhhdofE+XBsYpf4pY7jbv+vyrDXcsp5TiaGJE7z/XOx7m
tmBnlnGsMbtlxGmPE9vWWXVCPN3ueBHPclXYEcF1yp22AKgGVAmQPSQ3ZlCy9aV6sHEGowdsxYMA
7zL6dHyNsbBvhMuFq0n3SEZmL7xt7u1oTO3Zn5J5DAvxqpPFt05vZ/7EtqPDNJUkbesa5ZN3sWfo
BtUI5J1mBX7OB0748BLMt0J9gOE4WSxHc0aXT/OxNie+r+55S9MBNhpwJCD1vYxZUPtDUB/Xwmi4
CEIPBkqD5DJyWyzo/gNuDSAcjAjHJBaCAFr73jnPqUd/y8cO4Od8b16gCBj/K34mUPl2si/GTKca
oBV1vFM3nMFJUJOwfvwI/02TLLwlrQ2NTsfkUCIGJ0OIZag1QIaAsab+qbUxH48iU3jKp5bZEg7C
ensf3O6vGMumTnxZvAwC0oyeryPZVdWuo4MaqenmLvlOnCs49/fclITTH5NdhGfqpBOP7Nhirro4
bXzZnJKVvKgds+kgsxds6xH+rAdlpefUOEUEGMb+zdO81Ga8FMBxf7ZeCYt7KepjwQelWyLBOn73
58cAEcqUqIws8HjgWEvfsGT3sEy5VjjfUqjOyh2BW7iPK4qUs4UkhK5B1tJ21huAMdROkoasE48Z
Rp76dF1tmla/rIcnjDipyKcr/Es4fOP7OsrE/zFHmtVmfGrE69aKBn461G7TPXR1Phy5QF+7cSID
UPhoFo2w1grKuBIR38PkYf6y9QXpv+KgKc6/3LPmzSwE3cqYv+oLhdpX8LDJlfT1GUc02v88CNR2
GvcGaMuUlRsgkPR/WYhBA7n+8nQRd3F3gf7dN+M/d5g7TFI0/c0qLttW0GdFb1OnhXz7lUxfO6Rz
NOF0jD62VI+HEbW96Qm0JldjRrl4Yih84Pyqs06oAIBDxFIgCbshqrsw1l3Bcs9NuJsqdsfYe5kk
httOhcRUrFrV8FY1PYAXDHg3RDPd5AzE9yGE9EP6sFPeCJG6prvftqSefZC0jVhqrOySHROJOKXA
zGzvOs/on8N7vlC07gwJAGBx26HDbSBSagsFHTe3QjM6NwWQGJtIYKj67YUyjgWQEAntEYd0nOeo
p2OdxuMvJBTY/2m8du0VBoVcfTTYaDNwDHK+/4AP5MfkXDEqnOtxOiSu0iH9cDkun8ciFQimXm2/
R1Vuh/vy5me+KQHtu6+6a50RnjBfQ5LjC0aVAraElJaUMLVr7KGZcuhJ7Gje+NQew/gH5MxzCraZ
2Ku3/8RhPiz8hrgt8110XXB29bVApxKStNCrXXTY328nFjtjpiND1E6YcEKcJNBVdZffniNWAVXv
Li2fbS9ZZJeaA0SivNse9wQaOeZs5XLdABctvsmEjwInS/3SmRCiv983cW+P9j+YXQb/Tm5PB6TW
ggbzK9spSmQBdLStKDMWQL/VQVmCJ2VacHVP44DyLRwKl4MavkL2uwXSjy3TstCTaUcDXSDlt/cz
pHgJBDB/NzL0hhUic1AaPBDRbTDzvigUjtGY83NSLSYxiw/wEfXV+RACVKaBef7ARQ4A1DcbRdms
A0XwsbFpDzQRgj+ejZapC03HyFEOm9p5FMMQRE3ySQTghitAv7J5DGvLyIzpZR5q0yubHP6A1dy9
wdstQ5l3JwgiUUeUXg6Y6fZND0fo5WD3kuyxXV1Dd2+/lL7gAtvX3E6mMsVQXen/LE4wVMyZRSRl
aTPiEugYc/u1m9cgQ3R1BUfWESjrZT2Xiyi7K4IzYHcQ+3FcDD+mwX+v+y+Lwqp7NHlVucmV5cpo
hTcNfHbexfwiTYGqD8WI0kcI81Gvqv37roesNHTZN/EETADUEat4Ft6DblXSpZNa628FlKUDrM5/
BzHJP6pp2/ZXEqyCELl99d6XI/wPna6b6uDdQm5/CTyMRD3lDUF9Npx4DXncaM1EO+Qa0K5rJPb2
q1rSexdIk7ybgSBcB786ms7LhtifZxZkSF393RzodwtCXmHNG9KQyoRaEEVj9ZV0kceXnLGzMFcy
bPFEmQHvHpBujsUzFXlXI5hOsj8NJU/xEAPD3TKFME6rzHYqtri6HFzkpcxb34U0SueFVHDXOghe
AU9y1bgrZoXMLZ54eewu1nLnD/f58iz7hFfyV1fYq5qviDj+fAG1BmtlV2PPEBjvFkBkblNxRfm3
LHx2hXEuMf6pUuq3ryKkgIFZSWqJsRXO2j5NjXts17p2UQllsSKS8xoxiJB/IhjZIaW4D9wtwtnY
Hda7F6B+l5woAnx5zOC1QfYi/BuU29bl6knWHrXVfjrJzEfrmdJHw7eGUdcWQbR60sPo2CpvWVZO
tJ3Tw42OOJMjQsvDgNKf5Z977r8IjCpTaWMII9Il0PaN4VYzmL35G1UriM7trpTcW2nJgJLdGF4g
GIu4H/RfT0zPKwp8TV9Zwkw3uy/2L0R1fqPA/jGB5LAzCDZWU7Rn8hotgUe9yAZ5V7rKJ/z4vfiS
Brtl1X2cEesfDCyyIAUiGqOn+supNtQBRzIbe8RyktTW9FPzfbxO1vjRFmHnEG7lC37JHrX01+3F
fBlYiJGM+xtL53PWtwadZ0Me0cji8eLn1Rg5iueJ1yaURI3qL2NOOSn+9f4WfEZzSTYYphHuMyDg
M0+3/mRAoTxqK4S7llsXzIbEV7SOs1ffwAU6Jsw0YPmOULV8UtddaSkh14ksCTOQ7MPius2/udrh
X++g2HYd5Ze1D4f9e4TK83oT1jzSuKGnSwXEcNjMIH7rkL+OgZTnst2BgiXivnkSRBlQ+ap2wvOZ
zcWfebLm28azPfaVmuVqVthpZCr8wpuib4OtQqNaofzAKoP56EgPcvx+Kc1OooVH6Q0U53NJtkTu
wWHkXf1kRaaBP/ABiy6CR3Mi4BI6tltKodA4vU7lJbwLkUGlvm8ZcVpVXqwVVPTiS82NSyUpc3Zh
oZup1AONiRfS2wqiKeenEWhrj2ytKLUmWxbutb/cXFUKFJlDKxH4Ue9/8BIpKBACcDmiWZKOLhPZ
/J1C9UacW2GqUYm9Fqbjo3JKVmFKDQJ3e1vmabKPE8MC7+taiwUDB3UXJR/bckOUoDbqgvprK8ZD
hOYH8MncO5jblG0GjJBXG8hTlobxmI20/YI3enOWvk8L5aColXa7GHsu4fvOFzS78SLmpqEuwn+O
giYtHKyNiG0okhPVHGaYy47T03db6i5wegVTqhtwflxaGWxnfF+/Qi84iE+994GrQenENLRU0Mx0
3bEpaisZ1B6EAnm+Yp58z3smNAgU/1NHBjejYIF+YbYsemj9BaKmQA7yBCTG3tlwv5rgrXZyJATk
7D89pSmpKZj8QMW/357JD22wlT7GfarszMCM2S+eL9ENDI8t4u7RSCrDaFkpMnsN9tslnSuCM30K
5eGB9gFdBGF/Vk+cWtVLYDxoVK+CTHHkLOBR7RKz25CKmzmFsSYvQP9GI4tTN4wZk2xFI3dP3yMk
Izmg+p5vYvMmMKMJaET4mlZGQ4VddnmdynqBZcFmjog4wxTgvcTEm//PSJRq2ZVX0eZegEdL18Vk
89YgVnlqDxXUi8ulIRbbo6e3M60ixIxATBl12B9Qiv7st5gMAa07OgSIKtypue39QqJTtYnz396z
4sCoowuMwuaBNn87xo5aD6fsoTocWeXdFnaFrxId9qFa/6Ij7iPLCya45dVlCG63+GIQjBUIFU6t
jwKQAiumERW0caYknWaNHYlnxAQRi3CYZLhW069p/G/wWHc6NmNcAvjFAJNoEamW5hiV3nw3hmCq
ShoBJ2oM2sQtz5GtR2pqbox2XUA9QByNvHx0uZ7GekvcofOhdxuxMiKLVKYj6IkfXRP31m/ZcE6G
KPMKrZN9XLwmiTF4UytvmMWZGw6qKXomiKMUd33+oSaJGqW8BYfHWPZLdCD7XTadzESbe/heIMvX
wkEgaJ4eUAXWdt+NUB6IDuxGEh8p1nXE9/U9NqbvvHQvi0a/9kJxQy0IIogC9onDw1E4Sv1y5InB
Ye1dpzkS0Eg/XFrxPTOSzFC7OJWNcuNHivFk5q/A0WXWWXLf2yflJ52zPYTUxvo5w7fw9UWxIYHl
WcyYnZ3uAN6sGywkqrwUENsRv5E6vOUYkV31OvusIKyzlj/Nxco+Zqo1TGB2GDdTFXK8NzOSitws
F87rN0X0XxtMPs71zvSIxd69g0ebkljYeMsO919vjuzHBXBOT2hCqEb2bYOjZRZSMFKfGu50jE9j
ghurn0jGJDOO5FjxrDkJwEc4BDB4/dKsh38bjpHDSIILu6yf5Gi8Jyk4ykRLvQn3lhmCGXZkqPMt
xpORG4WrXZLsc4/1TNA7ha7OqJ9WRcedA2+nncxdxN+3MWTCLbezavNytK3eTwEnzOMMv8jI8AHI
nfz2SaUkcjmrBIsfdNpIAwVAqRnkeHVxSGEpxhPpiiWaA8ondtqF7KX5LEDn3EcImcnleYOr60le
VSNlALs5PVThV09jBwcJDklQVeVsA+K0QaefZ5AeABygSTVx7YzeNCXazb5bzSVYY8r5jJB4u1mO
3ndugJv1VQXGfnyorMkilFng65FTIGVsxunZXaG0ZjGWEWWIV0H8vKVT+L96pO/vTmkoiB8gb9cx
FLktjFdqm5A7w/Vourmao5d/OLvftoofq8dIuaCPAdb+HzvgXWmtY2lxMEoip+aL9DZqFvoiaHff
qoF6k+VE9apzVq41jBpmauoIqfkT5nNxQYXPIcKwKwLCYV3uwcpwyykWE+3fRhbIlEM35lbAVzZh
c3TfP7QztWC1T23rUPCwryMXdORcMNC8TViPFlKUkgshkbk+s9omgOy/h1qynPT5kxpHpZkEvY1r
k/iyvebbzvMOQfCDBkPPGnC4RHme9IwDT+TYP8sc/forO5Z0MyvN2su9UHVlS4jKv4UVnFEIjEcK
5PkVAs+r+OoY41D92OcZFSzk2s6Dc1IOExi0WMmKxTaQXBWVsZLnFGAkufByJHZIOUUhEVCGXmyy
Hw6a7RlmHXS/N+WsmfAQIFfbi2LnDVoMFsZKoVmXVHIqbjGNIJUDNrfSeP8rrNXrAcRC0mH1r/aN
wFjJT/T3iKudHPUR4ss5V5IDcd/4CvI0QKtoOXZLjYmvnsrsLJXzVbW77Y2L6D5BlCBxEbhH5541
9DxoMAGzZb6fZhWVqmYMppJyqClxRyueSflE3gaRr5M4nverMTRp6Xl0DpV4EH0U4ONjWUguoejM
0AYzrEgDgMSv/ekvyVX6b5ilBQS+QyJj6LsLTk49DrOacNbcS5aCpJEx4p1uFPmrbr7bKyh7mK9z
yRG/NQMV22IU0nCwhbKaHIUgdmlNLxabtB8UHNJmdU/QJADspNLyEbaACLaZZ8mQR9KAQQQMyL8i
dDpv5FMK+3GCuULvJDjo7YDzJdbgRQGptS8fGtyxn+9mgFkJzfieEGHVCCTFL4GDzLqcP2+/sG8c
man/+9uhqg33rmxiVXHDsgrRIm86GHm9zOKq4+JXaIEZrIx3+hYboipUuT8S1+Cdt4msXEd71tDB
4YUyKSVSYWKiCavfKsYdTz9PVhLedCbXBS0qDJXgi0wIXeNkdYAQfeqYfAJt+u4oVt+Udgpyfp+i
tcCUvkMVy/GLYTVtL0gSmlvpPxOrT7v7dtqhuvmWatRf7tBDFClKBjC/sbDNB2pw8bvVz/uZ+0Dn
JYFNGMZVIj6D78Kt+LyfpiLpYGmcmGjk6j+sqaVbfFH7yCm04yMoQXKtvmrpTxQiAqEGjSZmR6uw
KapdZSznsTS3RoE+ohi2izEkm3m6QqOSpUn7EZZXn5vmamvK9c3G+XK1lf69vyS71kHq/BUNJQGc
xQ8ayUoeD5BGMuJh1bC2TBxnWKOsoz9WS58VEB72EInxBEL3iuD4YC/yzBbboRM36Iapl0Gl0p6w
MwuF6os/cRtO8Lhj+acjQxb27C00I5m/dSVUwwpOyTsy8k8YoQx1OUv7d//DGCaSleozHoRLigK+
5Nw4TX090Or5rZ6/fDxw7g12gF6kxG2gBNV41YsPjpe2GYPDBP56pio1o8pf5W7b+hXF0/etQS4w
zmP/vMO2lTEQDpTIEDYKskPAa/Q+9mVBJrDHSQu02DKQAxQE4X992UgT5/Ow6jAmYVwycGskH5/o
zTdN9+ocSJ+x9aSYxJB9bpopEm/onm7blJ3UHRsEGGrrsXxUnWeRF9Ci8/VtxbnEidFShJgnjVrj
vNCitCk1LbioktbBwNw0RbOfmxqjHJZhnZ+jsToYZ3hAGfCHnS5BatPq6xpZ3RGRaeP6/ryCbPwK
F+zGgDI6rkq/SoQaP9s5/2QrTchZk4dJn1XIL9oiGQsPqDnpvc2xbzaax2BUBliJk1VNlnmKetW8
86ZzWO0B3w7bIa1+h3kroJUrx/iBjo3dqSEaSFIr4juFIxUCZkdnzrc1SrinSf2yXEkId160CWpF
HXEPR9hbamUs5guqQAAd3omKRfA4IROCyf5sud3bxWYEnoSJ5jMd0wA43rdBuZdq6hEL5R79d73W
npVsmL9YqLdKxPfdWhrOqgXIc9kXGHTHJ0lq604s5N4SOOF6A4mSNh+VRbsq1HHGzHRf9Mq+953s
Bc8zENaG9ybr38RcYCK+Zy0zvGe+GH0lwUzk3kpvqkHvRNo8cgmoABKmuDi9gNHDvAOWIcq+3ZSn
3wno4uGclzGiokCCoLqX+06BfhaPiQQ5D59G9rklZqHe3XHBfvEhVg+nrTQGtzXzEUBYTROXmCbg
WYZUYDglfZ5FQkszXgmOHPrSGba8DcasPvaj8leJXYRDrDOdzeTn8rfLx+Sr3A5Wt9qYmGTCzNiC
mPAxC7HUfe/8HyIdWjgizOdE49TLb4I9xjs6cARCM8hvSn+uEoB6kMGs2qep5yK8diSidvJfUqmN
oxKLt6DBJ3BSL1PoQ0FuuJGoN/X684+y4dfdwpHJ5DVc7QjCflng8dq7CTmoV/H2hu7Vn/pT24a8
c7Hc/xO/dk62Ly7EraoG2VNLjeKL94MeVlSHFkKzNvVqIEMvuYkDmRVpTksWa9WYxmehmpPVAp7M
C1LYX/GKxH0JswcnlBSomQF73vMv85t9y+pvY0jWTmxDLthJ/aOErizO1VakCyB4N6T7UxJ4SE8I
K6eYwvhgIynS8npjr/A7LRCc4WbpBemhNPoKzNyCeJvPOFujwe9D4Pzi36smObctykpebEB/tm3h
wOn9TzT5sgtiPmiLgAJ8WNj2uhNduXWOfSwEpYWMwO1ZxHCbSsHk4E0Q3HYeMBEHwEdL03p57rrU
eAIaBge/msL/Ch3Gwa+ttszUGON1s/mYQOMyzzr7x9arpTeI5gWNc93GweEVJukUOutHZuYSNaNT
sp3qDqR2Fa8mcq1AVFBRPK+9pGGPK25HAGedkip21ea9/QMnxaQqHRRtOabOFZgfbdX2qPfuMvmg
APTEJRa8pqfUm0yniBoeXLyh/mBwULYSVRnNeux0Rd+sNPcuHxUJjWZa/rQgjgB1E0Ee12AqV/kZ
UM+NdxOp+ywFVDUKzVDDyiDJ+OVVxmJft9MQcVku/1OtP9Zzh4NPqS3qa3LsZacdyC3UKQ16q6x7
1vIdhxgkOEW8AOCQI8dsG9ZiE8cG0nNywOkHbMogUCm6oSuGmFaaIRyOB5I87rF8auEZPeHE0Ay+
64SMbJ/3dCn8uSiWls7PxXUBXPcBBC0q+aArUL5FnGNAXVW8UK5vMoNTuOfbba65Nhe7QlNgkMQD
IsU/bj6+JKBtOkcIUHfJ7byvmUYpcYrx2kQK1mdLrN4bBPSlW+fGxLILFDjHGWr9w92cjsjlWvvD
Y4QwvxewHkPm0CmEzVLxRT4LwHVsxkggjseXkeG9wmLyHzmHR75Z2Az/HOwazAtLbEvHBLAZ8ywQ
vOSz78GZe4EM6uRUyUYnIIBNoNTlx9ewrpHa5PYmVCGsLDRwzU4JV68kf124RtOOdh+LPn2ioq+F
MFei7HavMekB4FjsZ9UuVioh6l8plMSVNvypX2FjFBQPfimbXcnh4rEu91YDdsYwf1iW4qi+g/RP
+jKtfyg8wZpCu+qGe97USAt7A75upZ+8gvqXRS9RBC+5kRBzt3mGcG/4J4Rfifn9x6qCTv9ZU6Do
jOZjY8sy8qH0JmM4oKD3S+otZPQcLuDhLbeDUF+iwID60KYQoXR4FumObjaaYso1hmGoqZqfszqH
DHyfP+CiC0q0xBht7bzNsQ0Rhe+byp7w+6xsM3HCAAjaA1qySX4pk+JGcVFFLyxyQ0Gj407HxKak
S23GXoCEvwhjJTVoTv2kYWVPaAdxZsoe+egwJxjeAo0+PxWdotAWwf6XI+ZoY5VH3KU1D9+aZ0TR
BnHj6qk7AgKziHIkjh1qgOTCMUQE9oRnB3vsVQteE/jqIFjsstTrjgjc9/V0zkTwX3DJxSRVZjPd
rO7SlcUt9tzcX2nQZiYItOZh24E0YliMITyLOhOnRqw9hvRTKF+3d7NP4DnF5ncgiisj84lPzDRR
nUqZbtse6QfSVkhZOA1npBOxPBxrUIRjHeZdzNXgo63q632JO8StJsnkHVmKH/bpmMgTa090VG0I
94nEE4k/mrJtzjUCY45ZJ9eIOPFfMgva2kXtrHWVZVdD9ejqQkWpqR6qrQhjbuEVgF8mSc1SGaAs
JKb8PqwCU591qDw82HTLuA+PailkCmGSK9JXHS0oBicu6MBzLdzZyYa/XufgbwxDbbll07L50HID
yTfnvusVYS7cMqovyIIP2xnxW4lz1ju1VdrJ03Kv7dlxVs9Mlq1LbcEqR6/lqNQ6o+OE0p9YV8Sw
BZqY6i5FVwKNoCXST+KREoytOfmEi57wB8gmzGX3zXuNbaLSrCRNNTE6TBw7lQxe9FZV/gBwdo4r
owlWWjEjHjQuYsglRWtlyLycKMfI+IRd9TdYfcwabw6Oy+qCQyudQgHnmkGVbmhJMcp0N+oVNoR2
ubeTmOTFOlN4R8AeNz37tIzUfOvdtQmJhyrcr81MOJIB2a1HZxfgtC/85e8JQpO+tRZorhnbryLN
aLHx0S8fIQq1Z088XoyZc9ehaT7mOioBpm/9PlKZ0wcU/VsTibnQlShYgjCveDRwVpZVfNs31Tg+
kUIaJB6TI39Eb783gepwGjCIta/BF6Bx+Xk990IA+xwygLsWu++t2i8z03yioI0jlC1H4nolEVPf
d7NCXUJMF/IZVSIYFvI9dzGuzXeAxw7V63lfMmIYV2alpAlr/caNHyBVIQcyjZ1GjF1aIojp+Ikj
NvJmCPs/v2/gj/fyfGT9BKXauwP04QKPXcyDCJVPqyuhm+qNX+4wUe4rFMWbr8eus47R2Dq+SnqM
UxXYhgEVzYlEwzfHr0fbSSPjH4+JLwdbMslbnji4dlTlT9gsHBejVBuSFtveuAB1WKV7e5OXt9DD
npb4FNsr04CUVH738YxIf0JPE4cdaKuAKo/On2bfxVdlO/8PFWMbGtiY6fWFsQqC0sO4SRSfPqSx
eG454QcpsOrS/gP7+3CRgVqO25bElUg5JRvrEHwuEmIMLJQWiSrgx0p/xCtkvNkjLELP3WtUM9Yu
H7Bvyks2WKskUg7xjqGdkXexJ4bxem7lt8h0LuVSS5IoMLzh7edoA4uQGBkPP9f59+1uwih2sCZO
90WB870nC8DHbtStBea5XEuxi1AtD4p7XICgIsBgJCYUNcmD8fUvWrJkuyTWnmQX3VNXJEQ71oyK
WqfVfyENfJZQyDcCrJHQU7kdorJ1+39PjnuZ2orYlNynJFu5N9UJxa00RoM1NCZu+7skUDiubHu4
0AImmPDbd6a+Ex5mUfNyUwLxtiuJHhysow1bJA3XrEVaCkUyuuvstZIpMPBLI8TaSb8vts7kfrmj
0F0kCawJ7w+z/hHJpekuanBcM0CtSJqOxeECkN7kxeBx0vpcWWc5tEFiGhRMaXX8Fvf8tTaeBWdb
C081rjHc9WTHr7WN5MM0LEf93vYETpeQCkuomHPtdSLHceO18Wge9ixd4N1nQHnSwoQaxI3g2v92
cO/tDiHe9QzroPMR70Sqc8C6TikwJ4ynDtbPEa883j/gtAubCaZJHy3bKqJgBAHzvbYJ5Dz0w8Ou
Dq0dKA4W1thYdxhipKfiIu4Eo0Ywnalnd9svQzDc57XxYhA+iyRH7Mj1sClpsPKsBPpVipWRb82C
+1CPwL88V6Fb8+xKoO6w1XcLpbOkBBxf/IHAlmrAIgFB8CZakXi0iyJJg31yQ+tsf2/UFLc7mTUT
SKyL3OF6q5QBsdWeMRnoPXRywQe9+ej8fkkV+haPPbkb0LQjComtfq2tokb9e7y8fP6E/nW6jWIC
Y2TgVlxK1Gp5B2qokrGvzqwsqR2hnymFZsqsrXY6tjvJwJhx0QlPEbrHaRXWvk1yIGMBCVBilDBD
1RMO+Q+o5+lmrJ20yLY4EKvbuPYaYZ53/Mi2HeGYoZL3/VaJWx0wSyCYKxGq8g6vpFA2xl9RZLnV
4+Am9ASZXTshWYEsLQH9BpqNfDKDmW4iXGcRJJFPaYAO3VlgA/ykECH1JF8qeGZXV5WgcoN3yYyj
dorwwAy7u+7pE/zWxz4RWiPRxDnlG+BVHifRc/CiFYuJlwHp1GkT7rR7nN/KJ2ecn6PuhT2oFOZT
0lvPZgBf37N34TdxyOZ8uFWffrefSVAuFp3JZ+RYJM4gG6R/wqigOo1eSMyvgBYUzJ7BJpL3rzz4
9Dg98Cn6tzBKSsS8oq+yEUFrvYRrbqAhSRrC/CkA0jWwe8uG0vZ9ujNDzAW1rayGDB6LzZctydqI
bjZDIjG7reUI2uAFd/e1DU406nk4pvJbtOUdlX5r7ycONrgBdZlNjXFVlboeZTGiAu47a81iiFea
MRk970N5Mjqp/lDxAFw74x+XMk32+HefW7m1n36j1jy/mrRjdrPhqIH/P/biJmoGMgii3hnjnOqR
JzLwlN3wTaUSmQlEk2SnkcePaNRqrJ0vXD925F4cRQuBBnQ8aEEto9ou57pwiXpWwEOFsJyBO9xf
Xcc6vvb4VgS7b0LhsiYwHc9PPuyb9yDrD0CmaIywVRBbP6v3NDmecorTFQjtZ3nBkGR7ODX9TblX
IHue4t96seJNB9rhioTluh5F8SQcW92Gfu2fL7I7+v9YdjU3E3iga9OvERmN6dSRd2fGBP40SCm4
KsP8V1CIjTmTrs+/HH4qzL5sFFaPSlyoqLoiPeRKiYJ287AQxB0kJxTULgCdTT5F9osykHshfvmF
KuviwaqkPCSG7zqWxetBADvLYfy9N7wRxUMUSyiPBgEoAXIuPDCETgGIKl/tpSU6W0KR7sNXzgrM
Q1hqfAEYyIWdLh1auoBp5VakA/tTlgPe6JD+G/5OiFLWyLxIBUgDqnxyZtyIaiE0JbAtzbp2M2au
4oAEsD6RblJ9tth+KzjMvLcK1k7mg9TTJzx8JolGWh54ZCXd1EKT8AgViletlOPEATPtUwk504Xm
X96nCMY8BbqqH3OVCljCwhB+4FojvQZhW1Zrw+qVqmEmhXlkjl016LCFX0DQst+G+lI8Y2jKlEzM
0QThhQYITUvkJIQWoXtbVVvvzMUN+x/4222dxWtFjcPzhUzMQBa0XwOIIjzobj/7upHbNCwm4RJY
ArcsX+qob3RxACYy13+o53pseZ56JR9rv/B3sX4ml0k1q0H+dMHolzOpdFYUlOHo5VezY1VeSv3m
b6ZvLP2L0vIl6Dnbk6T2bbsiZYi+ttRVBdEEnY2tKmkH564IhSp7M+kHJexhQ3iN4QUyLc8xVYur
cgpWa4WKAFuZBnKfs6R9e72Bs6UUgiaSEmnRK0XI4FXLKjeoADoYJRoCfvGly8L3YlBYQCTF/8Bu
88xtXFrfOoKQE3MCKby5O4dsgpXJQbUvBE2SuhUqBw8/xnUz34+oJIDwFcjVhIshmpj28eFodcVn
j4RR1C/QXRPjThxZ0Bf411Qo5lc1vc1s/EnYjg68OoxJ6sTIDiiKATkcI1ZAWqdYneQcFnA9l22f
/CmLJl8EQVB3CGpN4IUVF906iKn8yaR80xqDqX8tshxQcAqrMFJJFWn0d+wOUKT22okd7gQgWn+u
96sOF/1hNeYLEoVUsGJuFaYa9xCnCWEG1v9NqA9LBU8Dv6ZIrsoIs+/o9EGR0V8lmn0vOs5wiFZe
g6NwRNMaxtKFEdGCfalGqdRrujTgp1y4gIKy6AaiCdFU4GiCWa13O0uNWzTUvI7ILv2MdT0BxBs9
dgXnvC0bz1G0M15AcY9/FWHLkV7Tk6A49L+wZG+8sCd6LCK8G3fnqM5of9Gb2VkCMQoa7CMANjYS
HbVpQKCsG5EWedPM/5tSMCjG9W+iYRM8wMNi556XMgJ5PnHAWSKaDieLvw1cRFHMgzZ6DhvIHD4p
1BYkqB92YmWOIGxabhbe8xkzdDaxMLgjDg0ZvnBwstaq6Kz9ITz4R7aVXBgKU17cfgGfoRyAUS+d
NeatvnVyaWvfV3FJu5ObBcKUlh44gG3SiPOvHBCed0GeTEu/zCyDhkYj3MTYPWciGTTueg3Od6yW
N/7pze9indMzctAJLSWlFoLXxcv9Bkdu4l5MlpeupOQwwBBqKehX/4WtDUxD2UJ8xo641rqmGCLM
Xo1A0dBl6HvD5TyRuiznkCQNk1UVwNTF9qFCXr1We/bNaCcR92McoWkxJMgKiU0jBlYCZ2ZaVMDT
4nN8LaIDA/VLhYi/6rNbbQhfv5HYxITE2GKDwzce5vJzmMnc/QZ5qJKkS/NO+39O6EV9J8Ag0Xoy
uf4SHb5KRvuY0I5D/QsKAqR6kqwaeItL11ddSSvDwFqB5gZhnDIkDPX61WME+A2PTgYYV5/7UzxK
ve+17K6BQT2xE3aN0fxIiGUEzfMxCC0AlKOBlQIl8PDDaUrZwFpN0/2okoQvUDI9MBON/axqVyPQ
0+j4YJJwchqHaTNBsTp3pAwnbiNQN0INMMWAlFdsSdywRiekrAh6KrCbx+K2C1PVbKigJWJLNH0k
Z5pGON7GjzE3NDLiEO9GQ9QRwkPejlr/xPmW1RaxoyfKHipfI482cJFHwV8Nta98qtxrgc/GtWIg
dU3yYXWH3hiyv7S9vewh36uzgpdJwXQllmC0LrJLSDh7Fx40KB0c3ELIVA1U8oIb9OXBzgH+yayl
P1/a4A5Ccc+DiP7COetT/fOGubtKp6H6k4lw7AFW7zdqihvtR0G5J/+fKzSMqt/1LXMF6MMWwzlI
H+Fp5g2pLEgjdhgkZO/raFZPl1K3+lgbeT6Nhq/OlKnWFmBpm9qUedn5L3+fnD7kAYGTYX6Z8U+D
8FUf9kVGXasrJq3tuV+mi6JBprIFWGZ54ckijzb4epesknoXM0onWm1ciWnVjM6dSAriA1K29bDe
goN4Vfo4nKHcgp9KVvErFiW0Vcde1b+aqvwX6GuXpCtT9/su+SRIHry6DhJHLhINrLrM4FPhtpdQ
OZXc7UYhwlnF88ZPCbLoFT+U68WZuRSUfTgK0ZRXD11uz/1qeBaugpA4PHWHBoLkKJd9CDFoobHX
3RnpGys8w8vRgLyofhFKM73YophrEJs331IbTwAU+3QRtonPCxQVORn6DQkZ2WPKnacGMDj6M+aX
MYs1VCdtsZrtIZGuVs2FmuFWTKHLcpK+77koqKWTxpzjB8RrFo72m4gH7uDVzw3oRLDx+tNZY16y
il0LmSDtn2mh7MskQUFjY6JyqTpv3m1JKFw3qb5Vd9xuGgzNYeFa5ZnpbsPZ4JGS9AxQ77+KwM6K
Ytbfj4U3IkkUCMslyQtzE/9PTsoOtRSe3zoZ6IkpiW3VxLyaVBUTk4m3ym9VezLU2NLMoSIOzd34
nCcCNiyrsxvEKFrEGgCex/I+5FKLM61kTe8ZrF3NikKd5X3H59aIIMlbowtti5Wkx15sLze/7b+p
Ri+lN3xAnAhtumRSFUSUgP+Ni9bRNglDoe/4a9PCWfEUwYa7olwZVEg1zHo2RF4k50yU3F6XpZUh
BblF/v7HHGl06+SrIeUVmcWxR7zNdLI9Imjs2NOqEEbVaQjzBd/olQ5S0zj846slmMiDR4J5Vm4Z
Q3VyA2uyPsae7UjPzfDBwATNj1NIR62Y9mpwyUwv9nSv9gDaEXS4wtTPwJcNoHeKSLVkhtQSmV7H
SdTVugS1MHuydX1ZYtguQqDsjPhAE+5RntC1zdFaOwFyLhHRKgl/KL/WRbqtJ/ij1ifmMu4+ZWn1
OPjPltmfzOsTkjq4Mn83OPmOXN8t6JfMQZp0yF2nVRK8+CCen8Dwl3rgdmMPxogUiBQkNvVVFEtc
gre7UJQMrXp46xjF/sqLKhG2o7TwAcmU9aT9ha3H//M441WEZYBCLj7ggxLFBW8i9cfVBxbqBCZ8
btnRTHy6eS425quy5nQxC2XDjSpT8J5A62P76QKO2t+E2s4Z9ghjICh3oc0zN5jl9n+pK0tc2k+H
FFia248adXBqfnV0unke9CEDrykuJqvxqMDrdxWnP/q5dYr5ODxdXjrYfado/1HnNgWjK2fwtIyA
hIM/HG6H4zUQgmg95/a6nmgZGtcL16DxRXaZLaoz6AMtGis7t8lFP+ZfLgl+BSU7OYci9y/StAca
7oXMJ8YI7mstWCEDahbHjyosGxoXyDbEcv756CFvUXh2vlDB+3ZmIzEpIpRl60LyTUPyBTlyVfgS
osKB2nxrYJHnA5nZ8iN/YcaUpdYQpUB5tUVXWFLf1AzXO+pZDqfvsPUfup1FN45r3L9fPBv+y122
NtowIV4K4bs2VXa+eoeFHFAT3J1SFPDgNougu2gBxmN2TJdmBIDEqOagtDHT3lAII+WnYzc1T8Ep
+c40viUT0V9YZ9fXFIVT4Ky5satNPWLVqAybHQQGbGxbMtstSgO2H0pLfQEiThup1M8+7tWLcI6Z
6rEgMaye9Qx4tOp5eRm7O8GjY3cBKyj3J5EbPEAnP8qpO6faWTbGhqJGyrCq1EXRsIB/GzfyX7Pd
lDAE9K7GdJQ9bW/fmoDcudcomYV+gBTlS8JMPZjuOiiiFd9UU87E9nTm+XpduVoxu/bhtq0u+XkS
Ham79HlfSwsWd8qgrnK9SYHy/U7IUeMTbH/O0fC1+FQfdG8t+gdeaHLECCv3t1lV7VV2uK5t9hAL
baAoJ2eOJOd9/+0vz7y7WviRpg5kd7DOax0IR6+8CRIxIAYgyRJURjYQrmcstmmrp2y5PaUO3IUX
uIf6UD6gSZ8zC+AbGzc6uJSu0pRtwLC9AL8mkuHf1QGTvU+nnkvWjP992nBqsVwXUBWSomW3RPDv
WeISwUuxXQLwEbgD0nc+244++mICFV4OptXYFpgOgOBP3iEtGgp1uIGlMotxfNzNV7mWjNkRJD1F
c/2cta/zl6CogKOyLSHulcsomvlRHSR9/vHg7ueW0Q9H9970W3k0uCwPPZGa2zFw2YUO+ElAhNpN
qUduYduXpa/gchVeFaCZ2p5fLrFksoe9ufap14+tlvleQ2Zaonqi0SwP0twH9PsVBQS4djAUV7G2
3AKMMIN6SRa72ZT/h4EL+N+t5pIpBJV50Bn5k0LO5scMPbS9hz44xHNXcz14Q+AIXU8QOrfR/aVq
TnS+p+ryjA6K2JxpAbQRRRFXiW41ve7SedkNUqJNBjReDGpCjRRQq70NTh+C8ezhRDhO4mNZYIXj
tgoTfqPECR/0wbWJ558+Jmf7lxq2eO9dCuSbu12QSp378uvJIXUc6NUIoKZ+d4+vclh/tBZWl1Qv
qD032L1g1TrMYnCnqm6qPxwLFjSCvyNvHfklObAJoA3LhXTbJhdQa/sQpZ0IL29Gddxfm5SHRZ5r
+2F+6P0oVmJZt2gaJN6MFTSckmWqqs9SoeY3CYToeiJdEHxEOrVLBeJL5YoafYJuktFMYO3nUs1s
nF7DKY+lUp6kWV4g+XuKhMC+RGqPQQzQNIG5Qyr+9tNV5X+p+Tkmtk2gly20rvDLDjPz/1tAjEhL
kqP+zaEUUnZVf7V8hvsGJc9sG7XssQuCymHb2bsXFPp4w+30dq2bv/JxjTnNNiaeKYsy/MosoMj/
pcPD76M0CtufCXsyb1oVJN8vzI2zSWpDxsqjaTm+39d6sr+vM5LSIqxJ/J+B+4P6ESkA83HNuEpF
elNMJHV1NocdSQv11zLZAmd8GoaBgjioci3PZ9g77AXFOMyuTXP04R7ptoOJjlfuzcrKUYaI6uAy
ZHa0GXFGlf9QgZK0RH9jqdGBswmbn21BCqX+VYEDcSRz819eklyJSE+/Ulz3oMAJr1JQSBTaLxLT
FSp0H8+jW3YwVhAdSNPfVWaZ02fls5K8igXw0VPcSJBdglKuQZyDTMbGn/9aVp1IZZVfZ9ykHeGo
8U5GM0t1BXZeCwn+f5xiKrzYCFMSAuIgiCoU6iKQRIm6grfrWGzqJsCXcl8gDgOmT/LeL5VM0YEq
CgjH2ZGhzKAbOu9Ax4yDu6+L/DkNq0R2GruyZIJUThZi67z/+5NDnRKu5kh4NnuFTXG62HzynsSZ
2fPmU5y0j3G+BR7GwrIOExpfWjVDr2xYWrUbYWoHypnspm1OdMWMmMtz7wXbNmR4N52JGwr0op2X
rP8ywD+c5OUesbqs2ELPoHrQKLh7JTWgfOEpkDDqAUJihCkJFdA8OXYDkkuGNaC3HeMTyp1RTgVE
BN5jhEsDgkX5vW+KChkRUuNHJmc8GSmxQcitu+TTwVVXO8V6QK+V8r+1bvs3Lc8Sa9/mfF9L8Lk0
55VaVWWhBBqVASgb5cFq4lZbATY3rlvA3+jxVqLnsqljNw9AhU2jZMlbj7OFzAGJN01pks7LQm4r
nccKD/sU2gn0o2nO9Vj9LxDLaqncpirECm1KBmDXnXgcM40DnOQb8gBsw7X6q2tB9jfAAtPCfSod
0LXY8aWcUgQUHQM/ZE3Mnv9BJ/azCGOtk79qVU/lnjylWFLrd178v0a6alYdTDye4EUpPqUVNzO8
Od2WMvXUPf5vmpNFNBrI1GZV6Xo6XcZEn+bMTfgcMSrGseIqnX9XIPlZglLZ2+N2msoy1krOBw8j
vap7WOXtNEw9r6xBDuKDX3F1FnqgpEOW9/5QW5hUdDkyRYYxtp12WivnnVny2BEQ0MV7Vy9NjSa1
ew6AJdrb3RZXctVwtGvasUxCilXEbuvCyQgEcJE1BzDh+MvBV3AgZprZf7JHYTWVDiGF1AeOc8Zd
ci1EG2rQeCafAra3c2c5x369KOF+uUIbvdUT2bjAdW3SIHuU0aB7/XnWdWXQjgtn17XfK1jwBj39
1c4ftM8LTQtkOXKt/6EobNS8m807fnDhq1BUnYyJj38IAu7wZen/ATZZ2COt23MHIoZ6CC/I7LoJ
S/dWQZgB70klFhABYf1eQWWDlWqVuP8vINAs59dyJgIB6s78SaU07LxM4CL9+T7Ipx4YCP7sXsjx
7OAjVRqAMwfNHTUd0MPbFd9FRYKimuaQkrgR4gVtTDoFInSom/XlHuz4by2rAmnkZ9TK57zleWGO
byAd3LSiEFE+4jwXZXArmPCd01xCTEkWpNRjYE7Ip2cZ04w9entARQK4LT26fmry0yhygMw387Nh
4QptVK+uplpsbQZtxRI0O2/Ah1VVwjATzSiJ5pZ4ZIcdAF19sgSoyoubQ4egdE2Of2VesaRGCgC/
U88ihwirJP1Shxjpa+dZ+LXSlzY3E5rOA3p+AJYYGd/jaHH+w/09AfakJMjGBSmyqT5o+zjWqibH
Jx+yJuhQJUHuatnPUe9FLLDNMhk477xxb0xW1W3s479Asp7UiE63VPosTqDRvwHVA1bwulKAMsjR
rxqapS6N8GTFQ57tpqWeGQB7lQ7WnZ4d+M5e8jYuAU+QU626Il8/gXQQXVj4IgMX1d97M8+wrpaR
7nFteS3x221cwOGmoglYPcSvq20Ruu0E2MLchkFhvwsBngiK2KKWQoGqoG67XI9sKp+w+UMiiXA5
vDiO3HtPFOSRSo4FyqVyu3WIBDYMefi2zNWFFaVbYyH4m9F9blE7I9PEPchVpqJR/Y8soGDtdP+J
kgkesDYcjhVZ9K7JGeSPavAqE6N0tYWey2t4/4CMDC04vdzXwGbYmeNesXA/8FKviYHoldVpvFKx
oBF1+tVg6v+Pigg9dGN/CbbUjEQxAtgnZq0zM2RROcwbFrfUVXgwIib4fGXLv8qabZ2boEPG1+sR
BLBIFhozlDR1ImJ9Y4m7esDN97+KYWBO62b6pJ3IebbX0xNvVNffw8ke0GNXYem/kK+VTGY2tBG7
CRuxip9Xlf6IGDLwg+00d0qUDP/jcxyNf/Feotfxv0qwvY59NZHRUqg5qnnSMBXR1v5A+n5cyn1Y
Eyb7xXLJqzK9L0hPomgCcXpZqGIL19+Yss1Ode+7coxxDHp2xZQ9pMaD08HpHBJjlrCrFmNLcUor
tbnj2kG1WlcVdCxe2KB+cwDipSR24IAorNhnlxpjbmGGM45zRY47hJY31RwqyEmseearqXRxz9Vw
QMAdEGinCQvnu1V9UaMztUoV9AgJT3+uZSRxZaO/wNsQZB/lXWEGidO2PNVlkRk5ddAZrjja0Hdk
klkT7zEUK03CT8TQI0A3LHEkM7QPXcX+7g5vh9BF1z234rBX7XxbxQg6UHWBxjcztTV9MoXNp6gV
0yHAXQYG9tDsVVgsHbgaQOH9RSUeZJJ5c3uL61pSiEDC5iySH9No2b2KWqho+/JEUMf57j9hurea
NP3e78M5HeXk8GC+UzqCq4q7WDsy5gsHHS1l9WGJ34OTygXZgyXFUZzK56kS9Qsz0pJGxY+M0aER
0toujiP11Y47ZRuiN0zr5fb1rga3Q6phmgcSZwY0YPJFDqvV1y/y2gvc9LsDHd5rOnK9iodmWXZm
SWF2HP11QoTLQJtg4aKDs2mFTmDlNMOFTbYjwksPkk7ywhh4JU0KYTRAZdPXWZTi5Xvjw80ZyPtZ
ZJxan0Mkr7CQnoXZuI865rfsJpRNMxFPK8QsQkp4QLTGC49zJS8IvtnWzgyYancxdfXA/gzeveQ/
pXSuQEiFVP3j9M1DRd8/N6IUTVCPLsP3Qc6Vc61X+lG9R4p6oSc55GJOabg59vhX95X0HjRQUg0r
n7+vIZfTuH/WMiurgSyiwumy3exzKNP5/1eMp0h+SYEQjtengjUDUSBp35nP2qjKrf653fKVtzlf
xMUEX8CQzSVvueSH40S6hchY0+FP1aXTUbfZhMYNkhD2rE7JncXfI2Z5htREphaUgmP7XwWRzSxS
A2uxD4usSFncSICkQ4fjbTJXrGSVIukzpaS1CyBvaXWBD+nP/8+EErbLr2ySSGmxxLegAwF7R6Lc
BwZf5KSAgfiQbZ+4hbOpVc99iyNnesQuE6bw/yNE7wWpI0Ej/60zPVn4fnc1yyFwLcT+a4D3s7N+
zNpdhPjJTEZD1HB8wiX3ex69Z+h3h62Wl2tMuy7iZa0LcvuvIpILyLXLMOxMZxHpB84JdpUs4Wbu
zHgPMXw3vZkV5GswjXEom1kNJbmydxnNxDgO4Lbs3mZsyBohmDpmJFsxFZFcFegsWxZcdjknMEi+
0msexM9Z17J9719uCp4K1w9l0eqOw8kJweZ2zsFbS+PvX4/fES+EobJL2CzKO5eFL0MAmNF3Nt9L
iOhqJbQfb0MvvrDMs4kOU4q2Ha950fv8kYXg9N7ijl88lysN7UgPDRpM8h2M0PTUiSv2MvV+7PwO
OHniujrTioGE81lTw/TUHfJdSxR8ImcPSpy4SWl0id2w4k28HkcmkNP51PzxpaBaI34x72aME4vk
sUZ2x2VcrQLzDygtyCAWthfnb7ir1aYlKr10ObsyNuXYnN6V7+In8hB8v2Ew8CllSEApluu9m1yT
SBCDQOnBCAWqZwiw/pgSS1ufEZzzWs1e02ni24YI/h52z1+8G/KcU2EUINZM0WnrrK3FoKDHlwTu
U2qbVl3IH00DFyn7brnyaYWpl3tfomEYRqsKwLMPlgCS3PZwxCbGDhIfOMJidkO0lBVhTovuFZrZ
CPv3pG/9b31CVsX+z5St6Y1nMp06rfdFojI4GY5EAQLrqhTTeUo1b/wxBslIEzE1k8o2pGlmQYo0
YJkJA9z3Yj7TUvNiXww/TuuEQZJzDiJjLtKMmEZoTdvjp8gdZMbtfXSHlyI6QOhElOwEs847a4hD
q622gZzq7t3XCToFX1aVTLCtCOIwn1DFxXXpxGI2OA4OXyeJA7PkUERLwhoefDDzUkGWwizZBCL4
OHek3uLsbQa7AvfC5DwtL0s1EnFyDejo7l/1jI+gFNQD/87iZHkC7yWOThZeAtM3Se0/1j2HbBGL
LHWX58BhMsMl7pMXDz3orVU8v7WbdOMM1ZrxF8igLm4jNwYA5XE8jZokBoIBSGYgxQtT/IvvtiSA
FmI9CNYMx0a0MV6CeNx1tWkdQH9982erwyfdTUhvsNPKyrSR47hLAlT2AC58vBOAy7rqhqoz/Ypg
Q1K8DJBTGWGOzKtx78ZL8CDrQgO2KG4WxwzqCWPR/tbkHZ4PeCnu/1o2xTiFh9jUaYHh3iCPo0Fc
pGD3BwMDHynrpAnqjQzcR8FoCR56hxWJmkm+mrtUX+5W3Jhx8nm9Peec6k/kKltn8B6Pxv2jSkCf
Ww4/gLY4Sp0GVxHth4TmsyIT8dmQ9VEKMD/dFUEPpLK/SLtajdTQOIo8Eh94N6tNeK7t2rQFjgPX
AKBunQZ3MWpjng8Ryfm44TbZVt8yP4o1KJCAZVKVHCi2pP7zrgMgqgNYwb52JAqORm6V3gVT7vZG
foTh1lK2lpWV91WjEQzhjJFt982sNZyLFCCUF1sNUSbQHfDlTxMIVocko0FouNmyB3A2qVsXTwkd
visZNXpawHiO4UQcRL3Fyq3tLYpvcDNUXmIy+cNjYuVJDrE4Lc94b27XXUg0nmcPx5zYzBKhyeU6
yApjYE2KlYVWQBUKUAJx69WRv5Zz3gdFpJf1X1MkUim8jnujxnjK3CO/dKeyG8x1TbdJcB6ry2c1
UqqmK6yqfHQJzUFy+ll44AydQlrv4ZSHh/am+up0qcVckbg8ObXwtdYXMQbWrGNAKT9RXYAEyCqF
OLjEz91FzdrMXDdXaSpfR1ibBi1LxBdSMEAbQy5IDP2ipOZsSUh9VO+ckB3C9/L2C52Xv5jBSD05
4qKDIkbYVUL144IWWX8YDTfHHugiM+VoGkBkS2D4uzrUYM4TLeLjJ5R4evPvhx23I0lJhQ8AdKzg
BRw0sN+gmnXeqUNsHaxzGgIVpsOJdlIJuUOsBQ9b3nOrxB6BtEbPni9HNeXrHsbgjmqW5OQIB67j
c95VeyPY1K/XC9pAik3gHr2l59loNWU2f8Vnx4yBIX/4K+WRZzerFdMJJXIGIS9bJOGBkoNDxpwg
yfW1WjC0F9czFWg+lSxQsprMLC4J30yQjBX6djqIeZg0IjNmHmKHSPN58O5ovinH6KlKZHzj2EfH
RD18DSibJfdDnar/tWkSkySQtQjT5ZqbFJ1mc10Ts++VdJtp2Wu//g9uE7O0deYA643qGMxuzLjl
QhLlhjfGHEYKMzV2o2MqEF5z8+xy7pRTzKEHyS7AcUWNDnu2/qFwO52rSMo2LR62rW0XljseE4nG
ygZiPPOs16AlefwjlutzNovEJRjOEIsv9o7C8BDD6+Ne//CN9YFAQyzOZOPVq9iN7kZE4RqV26a4
/LSlYLSzs0iHPphYD/siNi7PXndnAhTgUYnby5u7R1CF9flNr1VMBXUlGYEEIyhK4/n/Wlmo1oy1
3+w3EoAlophGz6D6yOFEdqCiKRqOr1LupCP9lWAjkJ/CJ4QElPQEzF9drQ0nSlNSfrgSli3PVEyx
BGK3TpBUvdS6JAf8pMBPOrdSjKG6MaPqBxypthH57CZVOo5UeaZtpG3ivBPw7DtassmmfkxUIuUb
19VGEYZD83FNEiHTS+Q72U3vH0KP9ZvlQ4gAgZ5WBZpV5ey3IvG/nDOdR0eTlH4LvMTnpm2XPyZ9
GW8067n/YvnBleZ+pmMv66+XWDmFgQgQ6LkfEuf3eXpMHXkwF1N8wH9kkKzS8ZXwrFeoUzsohuhT
+LnUZQaMxGsoFlUhD+Ew3Ybw9KAce6StPeGGCDsnO+DIY6FLJleDD0oNDgy9LZuNak4+Fyq+AFvs
VOxzCQ3TGzootWbZiZo10cviEt69TczBPVla1Um5ZUE7XyqknMVRQVFcjOARHtWkNbGhLjMMkNJf
EB2crE2kRnmfW0B/n8V14/lh8naf/ssCAaGygWW0BMqBsg4s3VrFfckVJ12jxsyX3Iw/KsXmPPqB
OZeaaBZS4RrkUImfTRFJ1HhmD/0ZAesQd9WyEQEAaTb6ujD3FxBVfh8o+9lqFMb0zF3EBWJY+4PM
DzHtETgLhs7IZASuwFtvuZK+z/qWGWpIbx5d8WzKuxcvuQSi0q9td+9ECcYIk0FWchnrvU86N3kH
9AcN3huy/+Ja2C9PGFIjT0OJWcZ3rHqb/KKtMrEFuf0Do8yJtlcF/HqSGbJnTLJ6Kdu5iWx7l61j
wHG1GOjY1fdDPJxWB8Guj0/hJV2FZ2jMRUaF8Ld7mRbc5NP0ibb3p0Ebg2mFuQ/01w9ba0wBoJ9k
Uu6ORED5apQbEkBdkkxmkbM4GzPN4y+nNkCM3jypOFhsEs3rJYe8hs0FdshEqRbiRryADKanY03z
owvvvmFjz/2BhqYyaf6AU4OBUVveFU9uGpLicJ5kMBH7kezx1URHiwhLV9go3IDmSo2cY4rKaCHB
yHqKn0iQ23xgBK0UuRBae80ZN5ZDcIV//ngwIcLy2Gk7t6DedBpbYKPcBnmHlANGkB24SLxsfdio
MM6L++N72qVWvWJwWH/QhqsqyEYlBG5VeeP/PgkNy0ibIuOYWDsf9mb6cCegvVk87gCKpS5pthp6
P2BuwGmyEnyapBaVCfb1zesaYs2kPXd/NNsielwm5mqBAbrv24IyPNfb2CQaEBzFR5FfMlshVdFh
eqO5ScdG0B+J8NHkfdqgjGmclw10va11lIHZYAmmC02DzSE1AFYEZeLsVR4Nrt5P71KgL5NxTHYB
Bxx2vV8YnRNumAwXjKwU32kCrehdr5mpHEejatFC5RyMNYO4+AarBfHwtjclkJmejNkxEfm2jmfj
IVkQNYt//5XpYvJ0c/YT7dD5eFfO+7Y/2lTVfAtq1KFH7yWQS3stMrOH3ugN69mpKS3xITVpOFhv
BBOckDZiirOMmUP9agmNqwvRmTvnL4B79feYmBLKi6Dsn7lIyeyfOnHOkOD/+KfLc9ZUhcWrnBRW
JNoY2AS+qKb9mBQoD0LbWILbQijvQS8kpDrlDrSpoRkeOS6RWzwBXXSdjbANQotLazGdq4NRMMc4
WfdmBSD3CjWekuNwAC5aXuxBvGk91rEa02IkFYhHTCDfulxya4fch0A2ROqCYoc+Dx1cbq6I0ExA
XVLCG6PhSgrh2NAlJUegqBoiPWOix9ly4+4QaPJ1ti5zZmkbSBGyRUk1EA8iCxIl9dETIgDKKmkh
NhOhQN7nGdDclMwJzVNqQH8qAq5+sYJ3yewAl1OzaXN3btiGN1Yf7Zdp2ADwK32nuXGOzj4Dj963
TtQEYlCKfex1/7jyWTk+HwGch4PrGhfgsfG6TJpio/J9gTZS1R3cqme2DVv5H2oD/Suxf2WpQS5E
8XAYlKMHhXoP9qv+O6WF+218k9VVxwC3/Ka2q+qR8qN6abX2HcipBAeDB5Ksi0WpYwkV4qDG457O
yHVoxJQzaS+waniwtu20zIfRoD3IxbVfs4w/aieMBdwAR/FKcbt4L2BO/o9PRgGunvkm1IenUOi4
EhgwBp0dnXARyH+pCdT0XBreEmVjnnIyMt0SKxVg5qZsxjiKOR3P7mTrxFCvJbq7Cp6FHVSTWPEB
PQbWA6PmLjY5uK8gZkh1HgH+W5luaQoOh04xp2UW7AKCZfG0wwr3WM/EXcPZG28tvbICU11CLeRe
wJYCktHr9S0oRBI7gNFyTV9Eu+0SMXcM8rtHz+em1jeTiaP3ESgfanbpKVEBG89XN2YAwh3jXZoq
nE9L8wCpQ9Zj8n/qmNB9y/vEFFVAfVlK+VPPj7xpeRvWv3WBPbLROJwK1buGZSnp80cYLCCgfPfg
Tt2igot+ekhGp9rcNd4M8ZngoBV3FwpVWfecA/i+kUABd8so22ENJFQ6f+bIx5EWeV/jGeNXIvb/
el256w3m4DOJ7151gZ61dCWw9wP+b/hNMJRs7U+6RqBpUXGd9GrQ9ulo/wdERYHhY83dLoJjJh1C
tAOaGucOyRcr+H52HOTDb2cMoubyaQZKpKiZ959TbQszfEgyc5hD+lHg1JdJnFpYKLmy1PSYvM8m
NgrsE+tLr6y3sp1Y9dDK+2kmn+i6+F2MJhwVvhkdDQhTXS4FVt0FlhRTVDJhtT23TopKPY9J/Vjs
LcjJIgb3o0ceb/6+idg6BmvGpLQ2gL0lYTfmwsst12wKM71Fl4H6Z7D4cVQ+QwVVkvMCAi8I3/nW
zDjBX12GofSJ0sOf0wMuvvM8HSfYjXEfBFL82KXFiERnvQJ4PcF7ekfgRW6GMe4TSIv8kVApt9su
qEf+c2G5RHiqUTNMDwAKiN+nJ2SrgjiWS7KYm81vQ75PfZnxjwBHav4K2ZaytfrU4uAvF43CgFQc
uWCU7uDTvKjJnm4ZEBpjqnC/uMXnbLy0QqgK6isWVjUIpy/uwe4iEE2UREm1P1CmC63xMbZaes2D
+fimpymudvbolYP0rmyllUwzNd63V0D87sjP3gMePdcjkCo/7bp4CWQaAoW//9lJiFx+Lcx9sPl8
/bbpyroGhCfSncQQVYUL1QFf2hLNcZqC9NFhnul/1eA8Fs0Y/YqDVN3KnLTAb6e9YuDHnkGn+w6A
XArYau61PT+JrFsI1H24lHwXCftUQC5qWiX0rwBK1fMLJJsJxER7FtXGx+gwT/fvdeQRxkdV0KTO
Z8nXl3Cb6yGgXuLmS1CKC8ZNa9mTnJT6UVs/3ExLndHPuq0j6XoPiNXwJMDdyq/8K9/T+cT3//cH
hbr+O6rZZnynSoyDJey6Xd4PKafC06tI8Brd8irZFDlPlWpvRZ4JJhMf0WVKPTGY5rNqe2veS6c0
7QQRxkKtgnKP5rVg3w1AHRxSXnwMzqNw8dmYUS78x8C9wNoMlyJ3BmJ832o4sWCtRPSkzDv8wZuE
fl2pPolDC9Y5/B6GH/K6ZyxBvpoDpnqkyvXtPNYdhb2H1B21jpyGlIxGR6zlCN8MslXdD9qOyf9w
tYwnfQV6gTRjDzykuMSnGx2haQXJ5j7FMGfOGC0EZVv1waPlBbehq3CG22ZAs5DDnQH2ZRZbM4SP
3YCctbXOMk49a5/oqtftjlRmgbHEh62TY0ASoseEZF1P15AfrYGUuFJTNoG5Gcrc2+es2vL91oqe
3sjYCXro0GmHm7uWdUbrYdGwgtpAnaYIgTtEXbHPA5UyZqi9rBA3Yls+b6hZFc2hOlsRVLCFGxU9
8WxFTLprWcb1T5KnCAKdBGRVPBV8+aCtNVrZdZqnvzOEQdRop3CXlPIEqBNCYTNXTLxsP2fZmw6i
LqtY+WyCO8zMi8bgenEVmWOcKMirjUtgYTe8Qf+WNlUg+912fM8ueoPvhKYUdOCuQtr9asN7Fbnr
DTfiBtQx00xZrvWvlKD2AMdpQOf+V9E43jVDGMi5Pun2w//8NRPCcb5TglRAL8QxYW9H2/QdOjkg
IiimbrZbnsbrteCEvBvG7kpGco4AEznA/aWMVe2/k4/U7uvR1xYjLjulK5yA/fu5l9XiwMhAo2Cg
LbpVBAaey7dwScmkMK2DpLwNN7AwpYBB/XUxufoAWe/tkK9RhXjkl5RVCj3t3NnuIJNqGL3qVdkj
rRgIXolujddoEwXUCVAMQJDXOkCyPOEbtWcMbOTLIBXZVcO7bv+71jjmnqiTjxq4qhYfxMl5CfQd
WpXqsGkVzCGoDTEaCgWlS3mCBTH8h7DfK4NF/t9FKt9B1q/uPioRkqiINAh7Pb9Iwu1u7dfl+Oh5
G7utILPUO4Rwm9qCcdR34d5+EylsLJTax2zvS5lhEGUtl/HOtHCmnHdJs/9hyngyVRFO2c+jGFGb
qiA0CnVdc1Td8UU8ok3tYQ4rGHFhQOnZOkff/d4ME83fvTZK4wOFUINP7vUsWM0vugwuIX7QYpvM
1V3yKBjST4yTgqtq9fWgtPDQL1a6ROSUF93xE9LelPtmkicbzPtfhewSpvM4rUCqDkZ2UP6DtLk5
lLjleImw5ITEZm+ln6fYalNq1h5cP4XX17rjirWPSNA4z7zlu5G0Vcu6EctU2s4fKdpkv4MmzxTB
1+w5rYwK+PKqM5k7VXwScjRSytugmrdOYHRMqPsLF0xnshnaTfmNip1WHAd7UQKNpw6jIplhac6H
fcI2IJyLk8may0yJjiz4wvvdaynPRSVnbvXwtGnKwc+85IBYk/xC819cYpHzRk87HTROzNyc4wLk
nH1cBSGMR79oJ1G25a63txinAYTEmjnD4erVGsY6mqnpD2Cv4WkvElNEtmXGf8xOBOROga2hkUG9
Gbil/HkqXcYEWifqRP+BRE7V2gbBpgHQkXZNspAnQffVGTfX2panAfQK6JQtX50i03BHei52jVYr
jUbBxQdmg+eQ+025djlk3dMhLY9w2pRmasqmEgCI2K7WGODjilXszgYkcJlMoO5z01XbbmaSIAGk
swqApT34/zPiV11Dvp5YXJgGnC3x/rSofIBVF6vqc/JJnLnUW0pRPEQwuOx782ivdxW0xWCU0XbQ
MYTX+tQh3PNFiwe9ExUKb5PcpQ7IGN4kDqQp8VjnbdJouKVgszGCqn7l0ERG7ScsIBojewYYERGt
CddlXfAlryOmQCZNyIlaa31xELXZu3HXo2JtQQA0ImEAuX1GA9raTx/+7+5AP3bL1OVgCHMFcQIC
1WdAct++2eVfPk6LHJFwQoLRYq0la8FkAo3pUotVRhihoD4IFkTfZHndyeFTNPjRO88igHZ6JTQG
jyDKXB4Hqir4rFlJWjvgN160eojuLXqNZWoXX7rB29v8pG4kPUVBM9GIeznkeaFUYbF1DEpotlHo
dnt4KFOPx9PilUPHou4rinxIxDvnxSZ07KLY7Fj1oIkfITAch+Hm0kdpnd/oEkg59CQgiXs9PmR6
APyIysMCHzqfCyamgiSE7knEou+YPL/wqqot6a20kQFrcplIcG531kITgvvtg1014Xq/plTAkEs3
9bf2+y9jm96SPF+bIbl6EazKohLEiZx+kYuVn6MutHGVgXjCGTEprLluw6W1/m53GVFvLF2USXfo
wUYDcP/Q+zyAkZocg6mqajdroDwpEnGWIndL4/cVaL6erc87VDuhSKNkz8eG31U0RNM76uzv41GC
8CSIuApkXvWE+SWGOfH0Mp/G59WE0zDrZ9DkipgGw5tX8DRihBlL/bzRzakrlKDZGYZS3HFgy2fy
V17O93nrF1p5eVI/3D5NKmfsM8ICGuRAslkFtOxNHuQ5X5AmBQyRMuNEOodU6cjddu9kJytlih/E
p6ntx/3FyvSF2VwSPJDT+RYvTimIu3uHNSMRr890qAcCN3KkmAcrbVfjgNAdV3/nkhS2LBLXx7+m
ARK5d7ijaqO3eokj2MVqP1jzo6Zv9RRqb+D95qJYX5WKMRO5s1SiKYspQhckAhy0ccfg0lfpfjHB
VndrG0nhwEPc9Uj+yCWJjZoAAChspqf8++6+3w+PydOB4nUcE+TLtKbHkqzl9KMp+7fBNLANWOnf
pj+EtdLrRmOs7+irn2Od76Y4lE3KdgSNvJUsIOmzw7rzopE17LTzYkf4W+y6w4jxiXbjaWPn1Kj4
CSAUPajT8z568tVYVQkDGLvB/MmCf64TCyyBWhGaqmEqCq2EyInSIoRhDp2IovtEUiuLEpJJhqD6
i+g0H4JogCe3WEFiHtqryxRJxvz9NFp0oalVUrNuUgrL3+nqmtuGmdfwtlDdWEWB9jvpTsa2Jdun
sJo6BEtyjCusxPHkivDySqGXTFXeVm3QUwV/FgHlZ54fyoobnfK0gl108QkyB3JxOXo5VCCn6mvh
bZ0lYfqD97QPaZl5iR1wSZrLpvtYv9ybfVRJbBj1y9+Y81hUpJzPqgGpYBFTcTke1i+7ZAjpbHXT
Ig4k9WmK/FXhqutnKyVv2/YsXH1ril39pLa7ApbVKI/+U3YmobYf+J8W4CtqfGnOEmyqSoqdOuix
TKQ6TCQUrXMp7tpXp+xSBLnieoXbrK3p08NuNdht/VwBA5HIlqr2CIgWg/LB9aTTMLMUKuVA1Igd
UvEs5tnUgazsCcL9PTNkGRwGFeyOe2xZ86az7XNLmUw3ylHkiz+DLR+4xkoTwiaIGjxSwZjgx6b7
GUnsr4vVGQyOnJttLrxvdzcfp8EelCe1yCxTKnieFkVhGqTOOah8yhgbejo1lakfs3V/trvrlJUz
863hr3Dz0H1bYIBnKUz9gJmNgFMzRvyDwoXj+gn2X9c4Uc4O/ghbXuqSRGFD61MYALesqS3wDDdp
qUEVddBEUWezsRJEZwI9gzYOShBUdBS5QjTNl9gKn+RGDSngJBw41AZrfj5WJzzvUZ4H9kpbXb5K
BMzprjV11l8dFLRioOgTyoLJp491fCVlQquDgPAe4VBUmeNeTHc2mhQLU+BsXIOkLLF5VmmOFh7B
7Tzz+n5ScWkc/eYrwDD1YMxK58bPek3uLTfpkf9rAPnNnNcJ3v9oFuWxCp3IKqelXN/Pec0jTPg3
XeXXDzJ1i3W/jwV78ekjPuDlNaDEMGL82jU/t9Svt8C5XBEACmTUiRNgK0SIxn4PGQem5e4TWUyp
WZI3zZITXNEYtUE6xHEWvQ7QbK2Ju2pz1+Qc5M3ZZMcmvdDQjMGL+udraIrAr2bpp8NQRR7SMoJs
2GIkPXOBHBK2htaf7VS2TQ3Pya2W4U3bAB0KWLV7mHmjvsFz2WwVqrZqw2dNhQkJjJue+cmJ0T6P
0akXbgZX0M2moZNMIRH6Ayo048aDDy6XF5P4nVflYwYPeXfF0EaNeQ5Ecx9B3LDU+VamOjp8nroo
RlX2Mi1IMbMfjaowIAK8iEPdjToPgwQ3R94yi+cX+kwCgnQbpVjdBM59vL8+BA3D5j8YavCNHcBl
WjWxBFwsVJBWi9ho7Mn4D4rmaBY4aeorNnWGOcVm1/igAun38QHETY0YZLfQWWKRffnARiGOE23w
Ku3rHLdg/gAKLGhlWpLH8u0vMjUpACKyP+GyAPybpCO3xpzLbjvIfQ+6t8RbCTuMaEZzZSRlP0Iv
4bq92Pt/SCIENKls53HOUzWvmTWhEzULG92Uf6TWyU9ayiX0eJkBFTJscDvQdElxW2e1I+cxQ1YV
FUIqDyE08fucIgkUPCeojOWKoJ+awRtS7z3N9b/KWcXCYpMRgAPPyK6nJhAsXjbpLx631TtHttL3
gFNo7+gdTtjMQBvSUSBbtQHP7oYrcqMzhyROgZDoqkMRDZ/Eu0LNoOSdyE0dTbZ2h3EAVpISspHu
Fp8JTxaIu+39qokwFMwejrI7OoMqkpxsBPnA7tzJ6W1akyatXeK+I/Nlz9E9OYETcr5Ils0Ws07p
RTqvjQUgzD5wZsWlCWqMRaeA0ccD2C8yR8w2hnPniMDEtzClJp/emMyX/SwLBd8LrfP98NHTC4tn
m7ZEJOvVajJwbteYTdyxfjuw55Zjkze4v/5jnrx0/wdjPU2aziZm/RzEPhdvXNVMa6WfsHla8snO
UGy1kuaHHJiUSseKiWAx/9CrsreA3Dihjshmc+P777lYFvwDWX2wWin5TSTaR6WOL2ZwpUQeOe99
GbjMRDheTml1W2v4WJRBBR3vLlPrOzkvVkcvUGN8a1Krnlk3Npsmi72NgeQit9Q7xi7VlSnvGGux
ABIsCdl+PP6QjGp3Dd5g2R6K96WGCyPR9vD6dG945hVuyamemKhiAa9NsLYA2PenZcAhJqmRh9Ql
ulxydgZ4QpM8Dr/1Vy4aiUPjBoTknZxZrHCcunA0PrlH310mDwolSk+Q8dBDYlw5oQKS4F+76tOK
lMJ6GVndtXZl7RI2PYHEwo3TH6gwo4eYhn6TvU3qw3KyAVOXjjyiOwsbNRwNWH09VpfNbeLPgcxh
IzMoV76lcqaC0wighnLOIqfy/SJO2XT/5Oq3g7jSBdIqJZ54SuTHKULGT0QGwKmQuG/ueSgmb9Ek
GZvEEpctqVjl+Osj9nenayA/x/v9v3bpwLdmohWiCassdKpAHZVOi0BYqR/0cWC/HBDTRGVQyb7u
E4SpCas7Mzpq0X/CmMWFDGKc4cAnsQk/VCX7Ed/SXfmCIsxCEFrNbIlp4lG/y6U1ygasFz6buyue
/Pw3QjhGSwW3tFMMVXgvxTrP83Fx9swOssMyN7M2Rel+AjQ4jltIyvrtwLqzHkwPVj65UKUqAO6B
77blZCQIVNkQ2YFM/RYN2BcxYHxTNyBmikysaf6I7tJqw0VsrLLjP5Y5eNsNH5Sme/LP01BCOB9/
CP8qZIJdhVFLafqee+U2wqUxS8I+37or/6oryeSlcjFF2lqVGLuaO98O2kFhe8D0rUjESJeBz3Mh
x4oL4piAc+rTvnfXY+89/Ai6kjy3VlbtRLvQCkdVxzmFHxgYIF/ZgliGlHymFcA2j1lCTt9iVNPA
ySkn0K5zkwMO6AXT2UWHQ4EOT54/CrCgxrBxjM8KWxtRdEueI/3dIZXIe1Dep5yJ7vV6vvsBuIHE
5CVNvDKqXFr436+vj/z9ei/1pGxDWt+yrbHOIfUvfakdNCD5zfAeVzithZzHawqXXwdMIzytN4RX
3ISDKcIwX1e9MYy87tJbqfebB7lQtJlbJiP95gK39BTv2jHiU7GTCkm1f1BkLzpmQgB1lZV3aasA
jdZ0shk4hmW6jz96e/Hrzv4s3BZrRPKQ6+icvoXlC7xOgy8PHHywpxDBrRa+QDDzV+BPeA7ogjsR
0EOMDXH9E6hNsW7DMzZLpFQfZZ+29G56u+3ncNA18XSq3K5AUne0JSoqDWiCOitSNc7OxoO9oPUz
dYjkRR/gCTGmJGfEMyZDX2s8v66dWxRa9PRDasDsWPkOgTPVJip4+45dB3/HzazkNVkiT197dzYM
trMhbHzi+hWhJCM9sKg7ZtsvfcmOQR0hWumSniz1nTHi0dB5tifGzchfkhBXQgKHEd+hmXE8y7e7
gBMxCVjdDGjqxRjRYIBTu0X973s1OgNvyQG63H7Ouz7kY0y+B17D8ly1bglaMLWJdD47A/YtGexj
SUaMkz+DYDpBY9jfCvxkat2pk6n5eBI+uT42MnLJBbCjzsOiI3CDymc4zcVvIflBytj7M0+dOscO
MTpOCWVQ03Z9MEqBcDUi9MZc5RADqgJICbyUUM/oZJGOh1S7ABIb7PejCaIRByPPMkzaQoy8eup6
3uwWf/ZVOODwpqyXEGCBEDnZT6RXBT8IfTeWl6b3q0Xbz6HkIl4huHUF7YJF7PT6Mo8RwkmOQjvo
GXhu6UG5Nh3P7zzMlJAaLtrcdNNSy7ZcQFx86dHdR2boP+rGTzZcaxvPqKBcYKtu+tKXhP+j3J9/
EZgVrSisinSlOBkxQoKb0H5cmqPY6l1jDty2EFyJxDGG1Du5vOdP75nA67PFhZgM0sqVZNCV0O3m
fX9EQ4I5pAQ3ty8xYiXbCIG/ll9ECqWhdupNs2TNXnA6lgqZwG8AsOMuK4qmkwjBjywwQw/hEMzC
h1ZeHaGt6rxGT2fPNZHXdSnABykYw1O+2LI+pxvIntgWgPzHbapjrJIpFjODTnYf1Jy84ZTDQ1Xp
5hEsZTLQWyKUS/a0iGiZYIdbkJfVQEXZR+zoBHMFu4dzLCk+WbydVAfrOsJEOlMzz4f2ggKP8JkD
WFpJ3DNGKNhzblXzUXgK80PB8sOfqdkTFSHLz1NyTaXYjZreKmXTxeOWInAc0Tli1ezZNrB5/MZ3
n2i2Ny6vkX2FjoVwxDZW6Db/aB2LklMo0iUOu2r4VRnMQ0UhdrNoXsPqbOIo1N5omaIgrPjS+ooR
F0MFgm+DiqMjgfguwuOn7XOMOQmw7w0uKZHI+lFkRmVrpWxmnd9UJuBPNUDne8WM8BwXMpdZayQi
d3kcMri9i1pCpUeRKW7NXnyIM+Asi5eYWpU+lE414x2nsEJRVk98NU/xUx7gd8DthXTGf69zDwc6
92J5c0/3uiB1w/aY3GxeA5B0wyJbMtH4P3t0yx/zD4n0v2Xmax8M4rt0HO2pGziIB0XsutO7pifs
Mefqj+hHZBp5SC0fYg4f8Y8p1q46RI7sDCsnlVHIXNlwqWz1MQgGs4Ak5JZxc6f4QErfTn8BibpH
ULuvacr7nUzbpFSH86IR6+8/NqYJTTmpZKXACzTVvVeg8HEkOxKwIMHIOhYhLNX6Kdv1n6VaHppc
oARgGN8pqdVa19dCzFclocnthqeSQm5loNyJbb6aPKzT6v8Gr3wjbQvdd5C2UaXIzKFqHjC++v1P
M5pGSHlW/SIrj+kSQtiziET2x1D07bALFCUmpy1N0GQvKDA0b1RjDyeRSXl6qClFWXNLgC2wfXNf
4jhGhft3c1DEHyYZUb/W2/5UQoS2xtFCn2H2Ol6qoqAUnQ1/BwR+T+3UUs82NssP8hznsahe7iLG
JYrDQJSAv/CaVgJfstxOfXZaoUqwaBvO4ffTwV8+5mmMEsuaaRxQgkmNhrMiS6sqUty762JKNzz5
hNLRa7NmS++6s+LCs2TZRri8J3Nf1CPnEb/i1fIDfPPaBVJoyUEY6hJIP9MyNGjtAC6TevGCIIZ+
LxFHNMJlKD0iamnraV4qxtd3fxeOa65fuR/TqvOuphc2/lPOFvERCXQ1lTHlVJsyaZssVC+wyJUR
Xhu05SjxDuSieOh2V0tNyRyCdGShZuQKiBioW9hS7MTYR+sF2rrqNDbYjfMiOnypKdQO9GpQ54pp
DVjzUyyyvrIPGU+iIq8UysM4TzXtb4FHMOd/RzdCacJG6pvrN8ONIGXVFn7R46gKf6PNyz6vYPG7
6ndSCqH3mM4Mge4HfQawlfSKwSWcw+7ZYlkFEWS1DzcHcPWDJ0BVNlXJNNWc0+N/x4X6WCLDQ4Xe
wj04lQnJehcwIbXEXdnWrNnlF7kcBdzL40z6E85vwZ20A/6mNW8Sfo9a+Zssd7JpBtwsH6NSqljd
4vp7PsnvGwNGZ8SR6OuZh5/02gQVLcK9sDbzZ9jCCSFeyRcML59lkYiHEOX8H8+HS1M0doXnFbSx
TSYVlHinesjdaoy8NccZiqsBA+c0XA7ykZh6neMiLn7+7g6845YkV3HXN1puUKPmSwWPIMAReS3y
YZm807l+nQIw1i9ibkRzrh9f1vox68tUq0PeRbZMKVNebHJ/RNIiHdR7+aJC2/bH2ymD7i72n/aS
rzzgusGJh83vyKQvNFdkmzaN3qbeDTs9PE3CgXCUOXeI9el1qNWb2+/wC57D/KDhvJHqT9m4C/IV
X7joIXgaFmhj6yRdBsiNXZaHrgCUtSAuizY9EWDp2I5leindt379jMFmDC7aspVsvhhIBvT0QeiL
7NTpOP/C2uggakAqqMcmwlWE15TDAMPmOJzks4p/8c6pliGtEE5d/8Jec/cQgS7CF9fawSvvb2vT
nbL9f8R0iiymJX8mrLYFBmkOyssM57WxSiscN7j2IoL29YQgnX6EIVJCyzJvZjkFULRc6msSvsKE
NDS8pwEpPe/IAk3Lq4FPj+b5j2mRnMWqXSytMuhJlFvatPckj1F9UxmQAG9stEw5JMnU63rmk7H5
x/o2qBnLhnAzXcypDy0sfA7yIw5MoBy6i8wz3QkEhsioVlF+QFJ6YfPFX1G1BWlhwrlUkIcfhLE8
LzEc2DAuj4YFbgBRZ+CpsbypL79OObalbytMkMP98h7RHlop9lmZFBijgMXoFIIhsk/k7BcTbBGF
EtV74RsTMnDtea+Zd6sbn7U6jR2MC3KjYt2Z1+eLjGQKUTdRC0dL2M3Emqy73hz/PuCeWiz5RwaQ
lfcy3J9k8J8Y/M6MmwE5/SXEvlPbqaCDoP/o1YKAeC/w0h3hOlOHmUbkRHulukUeFB/k+V/yVHtd
gUaAy52LCx+IHqGEIM/NapN3m6lzhBkF3Ff/9c/jidXX0rL1P6vVcRI3K0qcY7uSXyqs6RZfjfxR
mMJ5Luui/EXHgWJHvrnc4c0Lil234Tihi8rRjHkmvH6/Da4SS+An+MjVa5xB0ez4yGQ81Wk4+i2V
UNFGXGx+4LP4+tk6viNypit+Jf+XZ/jX8HK/fyy9uHV2GuNJJr0N0eaXTKFjfhLODjEThF64w+yd
BFaX5yUw6gB4wIiiYB88v76IopX32ZZXhV+yd3S0x12+M39nzUNosYuRHvmfiZTPSWslYzZMj/zd
TWXT9i92S3pA9px7gWN1O9VN6q9091mvfdLvaZkcHs0HjWyG7zJi5kq59Ue3W5j01TohWa1n38f2
sn2+woqsF0QdapvvA0L2aZERWGdVG+VW571HT3k1O5NteXQ1dPC8bek/qLuRuq6tRC+FJqqa5ztH
SDVr8vjJxe/ZObnjIIpq/CUOOecEU7onrT4OmaotV6RJk3nabEZSbAoMLb9TZJCyLNNktkzlY8sq
esfDKrDRxVIpjH73DBq3NG7km/PbhCZIe56VtXhRFHoFEcVxu4rN/VE6LaR60fu9l0DtL/iXG7R9
TFHiqQdAAgjQ0CI/OR2SWXT6Q+qG6EdwPstrLt3rYTMJ+afo3aW+oOWS4gtyfIaZbeTontgqZtDW
G8vi/uF78nCiK8+d7AmlY6ogBNJogwXeDMtQGtNa+ajMPxQxxLnOqqIgixyXE0wNa3xefioo8p0N
coLdaU6opZwbaxyV/Jza1d82WaXrTpYkAhr8IAuyCl9Gr5p1HMfIySutapOBGp78hFetuhnBLP76
aRmd9OFipywOEqdn8scfc7xG6sdEFNbQIJtE34J7Z5LDpfP8+d4agEPm31cNvmstfB4qlUzD4QVj
58AejH6WTtfTA5XRr6i4jyxy2x00tX4/fyIc4w/SUuQLYGhMY23EWWx/z9g9T2lM8SAicwhp1hiA
iI5y/pMwHkIVpJ92EC2OHLejSZy7UPgKJ456fnDo+cHXVzZAk6IM9pDfE3lWIluGxLHKd2NKfblV
y5oBZINlGo43P2WEaxt7pJj1N9C+XOK/KmOOkbt3DBFNoqRwnePujofyDyQfBxSanZDGqGvQvDao
6t6cv/ywkSdDKACotB4RJhuPVSx6AorinqC5f7uC6/bVr71uOvmhk3XKZbM40eqglhsDzwAZpKH8
ADL5GCwdpUuNvffIfkjiMwqwoBmcnZnAwly1FsU11IT2FDNriBTneDFTFOV5kcqbUa4e++EwoAfP
MVM81962ZLyLtA4owTxb3UVR6XK+mhu/t7QL7YX5YSV9zS3Y9bi5Npyg02oeD00k8X6beDOglO24
+G/DhmyTjoXPDUkJsJHUhDZMEBldjkKfYH5j2cGMjNyKg06X9UcEe2ff6ZwSLq+odYJFnNE88anw
frNG1YZaMsij58vClLi5VTPLJVHfbJQwtzezelgmlNDo7CwVszuXSEDnexEWAFxmNhXJQSx7rX1M
NN/Nkhv1cuoZtf150oM9nB5BZrfUvQWqs6m+5yXv4bXIWtBoM03F/UKTVs5No9qS6sCgvKSoR7t3
pjsB22dGMypU7nKMluQayW3HHQNiltvEgd0V6rCegTgsBKktdZKyWde+z5Idv4w/RlXpUSPmumY2
8APqvSHdRxBM6rcrayTVX0aUzi4JzkYNChVCPwiEqp+zLGqMP6HaG65lNjW/RjbGiJd0Cwi+s6sl
5r/JknPonrVoLSNLjRgdSlA8vrtUICO0v+JILO/pv3cSiV+hOtFVMcbcGNvl58rhYZ5I3he/G4Sn
adnzwDWaSNDKdqZWVkFELuDeNQ9JGucVYSr2oNnmEY3o+UZrx14+QIGk1fBLD3L/Vtz6hpmDA8VB
ZWvsqNeJmAJSq9FJtG0lA/orKQkv34b0/TAtiw8Q7CwjaczVGYCvubopY5NCETrRShtK+UGscyBt
TpjfmPu99a2tR4lu6Uf2NkfVP+Z5IfVXxsYMQqO7Gl/JTvIbg/flurvokvkH3lMXvmnQe7HPpv3m
eyNmo8QvgPnNhLc32TnzJTgbRK+vfPd05J7WvHNNRWxJd4L4GXBBrizZVBatp2Qk0TMMlGt4UrWZ
GKQg9PciVoXzQTBJKwuYR1z6waD7OLzjjDL4lhRhIhBfWekT5uEZ5WAc0p+jBB1nzW7MMhf3tFps
0YRI4GH0uaPmJzqoiPjPPTZlNUappeLO910uIjj43I/Ph60nhHRuvRWgTZ/4QZdfIN+VQwV1mA4B
Ubf9FTPXdJC+0VaMuCW9FGntl47grBB5FplNYODMZ6lq/h+xZNuBDV9l+cTCmYXWDDVZwNP37JYA
iogNWW52alVEuZcAeoccpdn1C4moclvUBv5ZH8IT9PJmRxqpQ+PV84QlhuOVbzwXiXokf8d+F8xQ
vZMmB68I7ragh0NjGEwxfBQ56uxegqQORrX3+9qK3DBlrBahUxKQMLjqwH9eLD8bN6d5Z6yDjnSP
tjY8H6Dtl394hKMma/0m42z9jPyWO4o73j3qeZdj7/oicHDLHvpBAZxcw3fk5+oE0ZLOszY0HX0M
xT9CbGUYCtkHuAL5BQOP+gxVa/QJsQoZ2hHGI0Cv45roDFP2gdFGTHhYQDbbUJ+3qCMHGnS+qgKz
STmu+wKdEixWlTE7Jktqryf9g8VF8KnYGzD0IqU11r3OXrKqxC+OKlqXh0KyTc1YD4kKW2eaFb1x
26XLQ3ldIGCOMThBX76sr5iCaof1WmuXYWatvBucDNjzoSJTdhLVkMt6e+fP/TREO0S69Mxqx7I9
ilFtFLKbXNnpzUCLyOFNsVjshGZlg6YLCnttjlN0/yNk7WbYHJ3PgNr1fqRGUMgiex6cnwrskKzm
IOAouiWsNuXvG98+PTFIJBzhgEEjt8AbfJ+TUN8uf80OfPwZnkNPgOuw9vfiLCXnq/0RZUsS3lFW
D2Eu2LBs3hbDgsc9C+AYiP6ctRxIhZPYQ/KCEpg/TxEVAh24z7Bu9777rzLpw8VcrQgwzYRC5GB3
cNZuMBv+mW/crT746/Hfh8pu1SxePug7SeRhFxK+v5jVH/XGFDSpDuCfXspUot0hTIu/igEBFbn8
Xq+qIj/4q7Lavc2S0YT+IvxR6d495pBHiqpIOvyZAH/+UDa1/OojJhwCyNI4w+OvmK8QzHX1qJ5z
AUTrDjuKV2ZxXmLCE3kUkrTXm7p0DT7Gf28tQMmA5NKZIBkQP9dneTXjZF4LRgdyTXXvIC/UgEQA
AElW2cGAXxxuiKf+42hW16DvYPVheSAdZq69p7vXwcuo9fsfr+XxoTmkkRZJt+92GiglFilTVv6Y
qj+xKuL6u7Xe4JoN4+QwMJv/CRtHSGiejUuoCmMXoifCHJtMpUFrC1qstWSHuEgBm8ZyjYjZNlmc
mymRGfuShBMyc2hJoKOHpOArEEpNUHu4s2QNU2AU4v1jZy7dn5NyK5mNLAeUt7TmxERAFxWXzYOg
JoOKwToVKhSEQWSfP9o98KJDD+kVy22nUCzkWJvWkZe2PiroQRlljVt0W/1OVwpsi2NcR7ZNbppq
ArGVdcaGaogin1vf5kxsdRsFJn6DAOgBiIDJQvhbo8EaYTnqVbTxWmCux1G+jRh7QCr1kF1Vf1KW
hbnCzewdTuPcXyH6J7hmWwFetfdpnkigPA3/OY1QQjunZGtmy4ynqnHH/0fcF39MlkJ4gCeLVuNU
p9WKbcvhvuE23lBIHUJ0iZZIP/osM2wgIDcFvEPdIV8wVl+YC1ZlQREq3wnb2XQc1cFHQsCfArsK
OPb+veQzNb4RjXVTbrEyz8X4hOQQUaqW6j1JLQEppakzP8x6MoYtJQcDlK4sUokkkEobkTRD/Zq+
qu4pBKZawvTPdcXblxUB92EZwFUk3o1XO8GYSMTGBgjVv4lXViRzX1Yn00KE12O2y4hfMthgrCiG
B0YFDIfPMUw8HiIkQCWBAU5FXTX8TQtMSSH231m0eraK5iS8zqNOKKaGrnUGQ6w0Gq46UPJIHBAt
29ikbbSAqDqPs+1dAVeB0ICFb55SdfYzx2/NYp22lKTWWZRm0RXAKBPk5LCg6jrcym5U6g+ENk6n
jZhR3emEOcRYvLeWtcisd2J+psuWcHoENcmcAFIUaYsC31ZVF+1r/bwOfTewTHUbnzdBJJFYGj1L
+VR6/+u1j4S8AC5IVs8BOysohNQBkDvpbWXjrCNgkDQelYvtkzQRfBl/8UlMEEEGgfbYgFODVwjQ
eUjxJAeGhN6i2q6d3eUYzKnRK8f6TOWzsnHMmeg20Y5ze6BS99ipBAkjCRluyu15TU13hePhpH6N
Ze0c8ozt7pakxGAxuIxT6/oy3ozWq1VKi/LkD/vNEPcHqOUFXGL1m/rTYci0k3MqvLkL38ixClVA
sqe1FokAx0RVntTaY8b3zlZ2phDTCwYvSlDhFfmwk+PLRmKUlh2Yr5S7/lDEh3CV2g2KxRUszz3E
rundPX0xiAkVXktvnYIzYFFp2I1fMJLli/Wi6MB3ycogjN1pq/5unaEs/KCIO5T2WjXJIHckA0nw
pmhIPoaBKq7YZsknwiEuUEzcM/eIQvbKIW7+kwCdKM2zOs8M+7PXZIJm8KIabArD3jgxYf8HGoI2
gDNSPZ0SYZAOkKXuVv+CMXsuAWiS5P1H9jcsXS39QB1IYDgsL2piT0+5Zggw+KhALUfRVlrV07uN
C63WHeLTF02pXZ1J7lmb7d+7Iwl9dcWwVpUrSUdDr16dOfC5SKfPN9Qn8PTcaGz3Kk15dKtvtwby
6NKecGZcl8aNSthMFOtBBq4+4KxLDiAJOxVuciqTnroaxC/X95aRJ9mRFd6u1aWuu8320O86kR3S
5yswZFWn8LvuICHuvdo8UxonPkg8F1wz9y9C8g+aq7wQW+UC1QHe6wax2T40xzYTW06mE5PTBeH9
FAhUDu/uQ4up0LAqVw04NDDTcxEliJbgXLrpbcZ2eYPxdvRFREPdRja/D9ljmFVopbo7VbKY22W7
yIQU1B3qeRRcS5qvjyWmDAe69+JsQGZ4SMeJDSSSErwHqaUx6cYvhb8H2UsPADxlH1s31fb5uTUk
HFSHyADjg8Xo4SfzRq454dlz+QD4NVHsp3RcLPRd8iMIXwHtkK0C4uFGPjN17pQ7X+HRBxT8lR0m
Lys8UjJ3776TgcNVn2EXHAucm432KPERewQ0+hwX2tLYLO0IAaBmKMbxYBrqaNL4edOtuI+5IBvA
ReWI1tCkujdLXMOLIDlLdx3I3tpj96/dII9dyjwjlRvPSR8Nu2tFojSX99k9ifRi7PtKxgpFyRFY
RIiEiS47W6Oxqc6MGwzT5YTKfPAX0yVDGbMZCFTnawHnSG7fEArHr3otvLGDXm+0Ib6bqfDBMJCg
B3fJ/1iCwpq6NFcA7Rhp73bwG733M5I39TuysUfmATyhIVN4r2iR0GnCUMqv9EuUmRxs4pJzey2M
G5r8w5V8VSlNLisnY6N5JoCo55RGyg6q3gVsrDMzceyCvSwpIDoMm62gr4Ng7rAXtcOP2sTI/5jZ
dRW52QF1vlcRUSl86EbhDI8Z1DE4ZB6rJw88WVVhkFsr4bwquQBPRQWlEKXkBOsTG2/fL7YtRpwd
OVtHGL4dV4h+JeodwcFRmsC54bIBaEVv5z4bNqztIwh+gBI+6VvLNQz2/5y4YNBKghbyQtXplVPM
ILFE9fOVHLHEFfMftbg1aorvagbgBwBriMR0+HMz21ILVJE6f4TOQEUpRtX7SX/xF+PgOon0U0bL
g1QJIKTqCfAXQhHYWC66h6JcqCi3PBFn9DsjadalizVFwqYOJ2y4nw49XwZGC6bSB2dkQRREaxj4
gPMST/wFAfT0sz1iJwNh0DbddqpPpjM2LljeI7fW5QNgIW1QOJLBai6Pa0dYHRnJ1OIgU9aNDWqo
E7ctKPxt0RjKfO31L10TVhm/ee238qIz2GYZ4VPRlVDsnximrsYomOOWbLxC+waoRTdqYG5dBGyM
xdlSkVNad7xg9YhLZAQT+WzMOaor+9k57guUFBKYqNpb3GfxIx5JkaoHSMuAGtrns0Zmqu5Cq2dq
I6deuwGbhWiBpzTjnPb1GnhwNvbpL1c4Usvb2FCfGrfOiBNnKIL5nw5pdFgVNn7N7uyO4lmDivcC
OHgKFBNmw6NLb0OsqoC6thowmDgcKzEcuZO+dVKeiS6LW0zpUWGyncOj8+cAwh9Du71xsYWbpinK
2sngmK1nxqHDz+QfXiyVWWlM8HsK5mi23VQHGJu/WQbXOsgPfpBRHn4INzmFIHVspMaYmCpAvgbK
G7kHSL/SLHnbVbc8YYMaPktIo/QFrPKNmEsMiDNWWiTW/cOcZ/8nTLv7OI6nxWqWg413sFAyQ32c
8v8MkJv/BjuopqyHs02hvGxC2G+UugPtDUf6p6mJcl2tr+CYHwSdUOXLcVU5hgLiEqqbCptlq6xa
EzUB4AoCYwO0E1Eu9BkprHbqS40BElRPNvMOF+mrCzdHXZ0D0Fl6y7sdxnEWSe/DpWp+q2MdfYc5
2LEXU6aPKY4kH2QQ6es8m6JZEuhPSG+zNbuxNx1fUyaQqVo2U2/87MYao/nO/YAwBDcqdlryqBMD
jDJ8LrGzpjzKKCxk6CKVChzNMko6UI5hQS/kaiB5CBSH1nehU7P6xR504HCljR1UHKzYm69g3QOH
g7MJT0aRjTLqWpJqcQyqFNWSEP/uOcuV1++16b5EMy/xSmP9nTfYLUXLbiC0Zfxe4rq3AcrfjKPJ
RfOX86Gg5bF6kApjPUgznsxvKv984BnG/wsPXakK5JyLnXam6tKcGJlA+inmEMG1JzEhLiFGBLxC
YKkWO/kc0e4k1XK7A6dIJsuPY+2XtZezI9TTs8f9bzGT0ljQ/+JZ1A0HcnK7BXUXgcrwRfeg8xFP
hjQTHtGdJWcwwuTeJJ6UgdzpxJtxVdwex6XMMFkpfisfMs5Tc+wRsH2X9K0Nr1ZT3cJ5CwTuQnV4
sKQTp3WKV3kMFGj8/aBlZ3tQWBm4o+pTbJyZ4pls6n2YsqeSzwYfu/e9LYTXalK4/1UFwTzxo6EE
1+4sYfPkYbrtkg8wUZm5ZOxPyv+qxsUipDGsNgnzZfl4AMS0Z0eTfmX7z+hRNoRKoOum7QYK4bNF
+33xbnZnIdJDUUiKnI5SSYGZo0migf8rIV03dkNCKSzJhS9nNyA30NmQaN/FOKQVc7BCYpct9YkC
N47BZAlsIOJYlViygOISmLM5ngfXXSUQM4twNSYshEZmyTnKaNZ7M79AEqT6a2X5/6QdgNSOtbGd
87CJqCZVRpEo1isjvEkANcnr64Ar+1IApXc9WRs6+O7A6hI5PwfvcJDCypoy+nwkCt0Y+Bqj65mZ
tRZVesBHeLTckgxh1PTokJ3Bx1VxEKo1di7pZGxULCGhHV91QiXRDXlDjLp18v5TFcwnlqOJiJ9M
rOkutv3DDI8ETbxLQx+pNeKH5ls/DH1rFZQF5vV6adcgwwFf2MeZI5oAZeOuovetqjmmF70huhQQ
QO5xkLVDnLc0oRR3hhkAUumwVL3V/8Ev0sMARy9wcK1wlnG4fQHHn12TrbaPrO9Ts5PWhfT6ls8q
renCvhbLhCsG+KsQcoD2kyTK4CMFEiSmN3nHnLUx7iAw3llUbtvpUJFFYwN2dy876DR9PVMGEiWt
CeH4DsT6J9Waexo/jzfEUZwWcdk7YPot2nzuuIKkAm6zaD6i8t9vk5upfKjLtbHxPEPB1mr3lhx1
Cpc5dIFbhLCh6/dfq2WK/wDU1Lj/g80Rf9zUdhUIRkqpKidQk0hDYKo8n0x6nKgALux62E4kXj2d
F6/NRKvnReuqJ/3dTqS3brbKHN4IvVcrgzPxY59EqSFy096oFM31EB+rJhdEcpiJhFR7VyzTr9O7
zLbx4qVG3ZkeAWHC6B7C/9ZroYHbL6zqorRgLA66RcygiUpe2CcMNln51ziqdou/zogEzP2sUu7i
klimga0EqSz438ObP9Q/kxD7EBn3Twq8SSBav4842/ljDGuN/osLzhe+T3ZF5NCiHnpKZNxKRwdR
pU6S6tpBCky1MO8jE41wFw5i5U1ip2lXRBCtnWDc45yQC1TUdvua2Ly2yRTPTSqBmehM0UA68ILw
L7kRP+lLWgS0akVmPTD1PPIx1UjJx2uaawcbedCBwcldOkF4Xf4Qh5CFlvs0hiyHLckbHNJ4+xUW
fTH/f3xxvAiphW7A+/jMdH0gRBFNTmgA/4etDv8Z04QdAHXKr9ivmh6y9ntoEovYyZOHcVWkqXdX
OU0316+cXs6/GBt9KEOso4HABTmf1L6HzUtAcu0blJZ5Z8chnfdZNDmrWPkbK1ombFsKv1ZyWjyq
N041t6EyKUPYYnLVkKeozQBY4eqmrWB22c2JLl/OnVwACRNX3/+zgypDf6Go0eoL5F/ZRDge7QLw
ht2P4JiKCtEOuvpX6UFKCR0bpIBdAXBP48e0gFJeYSYdO8zOWcXjVEe3oEE89LD/T8v0WGJ/WM/k
IcGgfM3ryfr62i6iJJCp+TDh8ATA3a19zBKeWHFGAYI5wa5F2R3IbGgap4LcZ5sO1JuuJ1e5sKk/
PNoihKV3I5ah3tXokSW4h6Rxhyb0XICUJsk5Dc7YkygMZ/zLcUP5GoQpMPQ+Bzi5+7wlWC5kT4E/
e3srwASD6L5aa7dDlOKunz5bcPuhdnn/iuR8x/cBMNo81zGHfrs6zhgESbhPBgkIw9ROtCUMhYHX
32DiJuHJa5sqBC6yDFwVv3eMAtEB90dmX9Detkl1Bi2KLjJnPUMfiiYJQ3LL/GaCtpxolno9hkW4
thiqWmbcMg28TCtXNuMH/+byFBOFSFEYi4d/skeeBlgtdWanZOCPGNseLtse6Zxut5h4RPdL1Jcp
f46j7ORT5sC9EfoH7QEiGgqQBZmQsf4egxMQAOaybdnfMwB9CHIzIcQDckQYSpSXchKe3DDpiIxt
Lo1C7NkmPWL6yyCnEqRh4WTtysyNHETCZb+O9P/swjYQcRtPY4jHeI+tiuTjUyugYLHBJkvH6Uv9
Eo4rShXyiP1tZu4SmCKRbBw57S/3fobCxszxdoNYP5y6Pcny/8aGbofEpfIzCLwpphYz1kUgNNEo
eqaxMMDIG28vTY5/7Gju0ZU83wycAm0OOWv0uHP5Hvp+hEbC8dmFSlgYgfyuMWHPzuEh8oJfEGeQ
xwYNtaVJ1HUHC/YtF4C+r+no5P/n9d/LoBykxLmsPF6zSkJ3qYKL2mQNlGZemfrb8UR3Gc41uLqD
O1NQuPHKcy1rYlY/CWMa7Lp1PaeeZwZgm5iS1NH6AIaXLOdkmQK2fRjNfJzEvtQkEDRIyifb90H2
TB6mRdv5YQJ3L9Iljz/p31OOU5WxkgKmB3mQPXLOZwoCRM2Ysg8fGyT/Xn26CJUohbvhyA6lTkOm
WMwp4/fdPC06lcml6gPP/7yCR4iieIJW4NGHhWMRHrcESbXdn22bQJ+r7MNGW0uxfIlRQHTeJLgR
41f8mRYpRRJedgtL6dIAlFN/m7DzuM2kCxHlOLpYKXtYuXuhFQttgDLxnL8W0EgFtegLQsg/VNWR
O+t+QB77qz5P5AbobU8Ua00iWn/gmsvZDpD0idCTNmpCYbjxYnwsRw/Doj6+YjFSzubUE4+UVFvA
b74EFBMFsfGFq69WtY8cG7jBhLrywiE8jdgARJTkVyHKy/K6ezUfDoilMXn2YvsXMD78Jrhr3l71
HT7BolsEgSA9OholEQJcRO2mq8ALcpJBrAOWYfGwNa9LMZZe8KWVCmBF5ENZ0gH/V+qIrINTcUc8
+bXsoiBlsI+xtDVbOHKWBD+GoDZJryU8t8Cw71MvXopfjifr1LTNWqVRflxV1H0OxNzWGRcgcTGu
CT2nHpI2zOsN8qKkOgzeA3F5h7b2a+MNlxX47PufWy4QEqcdWJ61VQFVt1N7rmDz1rvsG6dkz+Pz
4i9JhoezLy1SaYo23JptA2e4p3+YZOvQoBfTcssqjkaXoV+TQCUC+pHz1e8kmkiBebilxEwqbqh9
KpL03osRgxg4q5ca570GiUiGWF9D6PJeijTyqZ6SnQIR7He1QxcydzzTZtLctYkFt0ipE3VpsdlX
FIH7S4sNkxhaLi4cwLfDq6VwfK7X669qx7omfk3DkvNWG+vx6uzmpChxxavJNYssCHFjZmVd2nFg
qXtpAnezYJ64NySGXx1MjLS5ds07h1OrNP7cHe6GqoikEdEwtjBRXxMlIuIIhMV+9EPqtRPQfg0e
cEjAsyq/JkYNbJ+tk6NJagzWK9kVD6meFqGnlqHqoS0WyKulEQRI2JbClUVMbs4fDDwQlo07n2un
o0kKDIkXf911NySa3ClRA5KEOPU8Z30wGM0UlEzsI4QKLPvlRiANVHHVvQ4fAAej6xPeYYUwqYOs
dUmKrPKU2UthH2xUQ0JyXqeY9a+oN9nInusGr5sRs18N6DPYO8TTC5l8Qahru/68E+6LDttWYFWj
JzSpvHshHHmUkJ9mG3LzsB0/2YaAZlRkRKo3fOk1FvWpxl9cDSWnkTuGafxru3iwokZRI/AMUCaV
8rpr0LbYRF6yluUhupKtRqNgY8Yygt6WZHnGgJKr9O3eHIf9S/mnn5JXTLyQftpS1koeSEGAPTIZ
AJUovoPczgfk9XMmQhfozU+Q9baAnMALJVNJ3vlhajWpKA8r3joCbnOojyrZb4aJeONP4/oTJv/i
ZP+yQHqZjcYAWHKg/fyxH8eGRu5BGt8244xpp3Rzi1rQBUPjH4cjCm77CxGvjHkjdiv+0R5/dTO+
/pOpU/vKphomjCKrkHDYzFbGeP2F2uo6ijNq01KbxERgZrl+giabWMqxffTZwJHBa7v3e4Fcr2q7
pZU5jruvjCSbbZMhqIUvzahbgJnJGIYvxYx9knkkqWeYi1aDnh3czZywfqCCxiqW8jmSU7aZvuSL
YH6miunwnrTfWq2TGHp8zLR8udAYKrmQHCuqjOMqwBsuq8KZbnSGqQ47g9msV2WgpcBe5/oMwJBu
x/TWRxUmjPiVZVOCshx/1GU76RLcje4QveBpvEkNVXKn+R+PqEsE9bt62ipH36LySHmSwI2ECQDW
7y8Qohe8RcUEAZC/YjIfSEgMTIdvKafKfwN4HAqvnUIcYOSAaKpTm2gqUToq9g0QeYBoJyMtnYsV
Rg+XgdGRd10q80V0dBsEw15IMI/47j5OiB+gaCAMHGFASSHpcJL2YLHH6RrVL+qjKXXmlfmHT5Sp
I+K7ydiAWhuU3KQvK3kXq+7rRAiTA/FrGywrKJD5euQnkQWCeZJVnonyhJGyFZs+4IYCJliaaNSL
OkEB1rlPu0i+rggyq9BKmzR/6R4qFJt0qku8xSIqWMuU7sWPkEnqnrUvnM9YidB76zisFTPdJwE2
QfY2suOK75wuL1yGttq4uyoor/Noc84mfQUPn7bN+N/Fnd+NvRjCnoFQYfLSYsZ9S0g+RlgDZAbv
vJ48qrW0hed8IpJQXvuNFvh7a5ap6dvqaiVYpZiRH4BtSJspikYA41Sijqmfl5YiBf50CxSVQr/C
NsjqfPJdhrScR/FigT34SxdnCLNdyGlsT9rJBwkLtsBtLUpD9yGgx4bY/cuSnTdI29ClGOzyEzuc
HVdg9XdaXuvvqR2ZrXVV1Po6tixPGdXYH8jZRI4RxD1JRSEvs/5ShoVvBpIQr9SU9jZ0ZXJ1mSjb
FnKC/ocbaem269ObAbK5cOw+wdDzU+IzSW1WoKuOCG0DoltSUlLD9CPxCnYMn4ld47p6aEbR43Wz
Pe79IjojRwYgNO8+Vm/UufxNjGnr5nhQFrdMESxWS9XRBKPaArlWw+xjVAh5ZgkiJEkx8LP4Go0y
+NKcOxoWOse6QXElWkwF95pdetDQqIA1F96Ho3OCssvUoDXRCMzL9sNZGDoM+gJqdnk557MBcAqm
5KmCvQE/0Ata2ah9gPgUs0yW8iciUHcYMtqaEr05JNRburcGddfb4xNb/fq4NZCAhr39XStuoKgO
HRf0hCsqk8Vj8b13lxvgtKfEF/HjK/us8OInzc3xyRPVc3xOYKKI7ctWFH7DPTFjTp02sXAA+nkD
2sogn3wUzbESLLjDbWjZImWDL5uf1JxPed545LrsOvEd7oC3mDETGw/OzO6IdXwuz089Gfbs68WZ
1QQSzACOueFfEtnJ7CSMEvowpB4wl3Y+ay9ITTRJZVmRHelySkRuDNkUugpdwXEZjmUqi+nS1YMd
MX4qrIelWr4Xi8zyDYjeVK5c3UGlkggkShmd3qFDQb3Y38bAmp5g4hfVgnyH4ZC7Nji+uy7o78AV
KSpNTcGPf0Sis1O3L+kqCW9dcd5PskDtu+zqsyKoNieyDk3ef0UUhrNp42ym1QCQOw4xrfYgBIGI
8Dec8m+zZHg23e6A7zeqFTIycZPEFh9Rosy9zwanN7LtkjO+9XY9ZpI6Oiw4zk1U6zYBwewJJ0ZT
55uZWndVu2o95YfLoyiSCjZZe6VkiA8K7+uhUV5sywg/q99a6OBPMUeuBxjRoFPAGopZ/0GhSBrw
wkLqYuHurXNzmXRECr/Jqhu/sU961yhQH/4tzkY+qYqVBCY6OWNIjT5y+d8ifmlLkCiTsGnEXd7v
1Kk8zC8NUOK6IcNF8QnujxqcQxGiuRH0s+p2AAmrrfjchzux4+PMeLFDuQGibAskf4H/oh30LwRq
DERHC1uvqhzxK72q3Y68QL1tBLP/v8Srmreqa4hknuZ5yCaa7eSkcBAnzfUtP19qdMzIGO6sZP1l
YgMcJ0pl4RKpoX4otEsPuu5fgd0TdngLHz009LZr8lV/lslaBxbPiTiR24gMPaz/NjmuE54TrbdU
snemDCQNPbOCwqBCSsKZ4fnnR5UmnxAugRFCSADEVsILcFMuWHUpQxcLvvQU5XZiUVK6q0ApKFnL
MxKnavf2+MnnvrgA+ZExhCZlS7SAmTbHlOmr8VIwhLRHc/wooljzgtD8TZBo6P3Gh0HVpMxyDDrV
fKao+vBxG2hPh7KBl90YvVePkwbu04vbVZaYVo2jCqNJlKivhTV8jKewGnh9mBbmMtqf/YMzJUv8
FXdvxjsJcOwLX9q/n3csSv/VJ3NoYn+HbY4bCHwaA5zcr8DqUV7bJv03TZmnelTnL3CFD/lzSszv
XO8Ysu5JDDg6epC8QwZvn1TFhMhqpHanCGNll24tbJveCVcfcF+XQrNX/E+UNNLlu4i5FOETZ+GZ
ivY3lPs7DRFpMmd+94n2ncMcZ27Y51448ntwQt7gdPbbXXXfwSh6UiM1uPEosEC+UUYp+Hwh2+fP
hnt7IjMKKxSTfrrO1FMib1/IU2M2Od5urvFEO6PAWrO3gM0JxeDkEFoMM5Jk8n940eEngUfEq75E
uOJO//4gA5sw7BfECbxvfOBt3LFsbUYVm2KONkNMwx3JL8t634Fb3QMykP+cciQvboVdnnL1E1bU
bPE+y3GTrVD0PKGi4V1svKNyv351J7XReyoC5/kvzQHHUEaCQF52F23Fg7Mm9eZDz35Ev+kyiASa
+gmW/XXQPzI85qWrUn5H9NY89HCA0G7Ek8X5MpbBPOvT70m7HpXBWys6RK1AFhtEZFZOx7akQVom
XTodAebFuvjD/m1d6NbErZLH/UualYl6nfszEgpyY58Hm4vvINEZw6Y6LKhGVESnjvTYIosPfZ5h
QSCMQgCCDL7pljPuFPyWLcydWwr1GSsgtpNo8vi9LJsOM0ybav0nfSG3EndhLoZztbKL/t5m/dq2
jTQ941H1TTYtKf18ldXkwtfxULgvsfvfKEnLJuHFYKzVRYPNxhO3txl5xCNnf8Zadvz1mCD57EMR
hV4iJXbmXnY9SC8R9n4SgEblTRuTBfEyEU8yIIjnl9QQ6AmVNfrEXine6Pr98P/427ba+zuZXbNk
Q4txMoCvDOR34AF5QubzpmHC5j1c8mV5q35q4g2+KGBS8AAgjEe4kwNNO1emv0+vIzWP5VAszCq1
WaZ5taHMAA/KxImAfuAwPV8WNOVDoXlBcy9AR8pyD7NGWOwQ+NohJYB8pPpWU6AUPRFwj+slIgji
nUmXjZ3HGxWhvwVsKFUvL59dfNm4NAB2S0zjlYn4aN/2URIM5MsP8P3oZCdqltYMKZhsd17aAS02
sAliD2dxNf/Gleg498sSY6R38LF54uAYWh45cXhn1+udP0JyuFVyXhLvrV2sycMYrdYixn8sGSDd
a2l6+ymO70siBUa0MiHQ4El6vJVmuA/plaE+k+Q4ElYGgzJbxDl9HEQD00YM0orQW37qCm/M5yAD
v+hzTZwYanqFNrwe6TJRjhgF6x1TCRGFEbVpKjtLmwjMs0fmnxocgUOPhu7TCHiOAncKLcPmMXbP
a4BjA7YhKWDWewZfq6U9PmGk+I4mOIy8Wgz4J8J6iovQmvUNjOujh/tUvecp/xRi0UDEACEXZXO/
3gseqesqA71qihSBtacGkbuCdHeFNhAS1lmOudbB7PVNafFD29jqGvEA7oscXstGlP2bwkCrmnU4
mttqlPnCAbinsZ/h4nQo5SNOj9q0gUi2Fzgu1fZQb4PFoBWBBzVE2tCk2LCCC1j2dmEHDUE722Wg
fP1TlEJMPmH+q6C9G2Br1wt7kJPZT7mtX+f+7kVjWkjDo0LD+BMDhvVOY90MyA4ECxl9rRsunwxS
s0LD3hx+Ii8uuyl3dxxNL6usK9SuMhDqcnSSauNA0za3ATbCFm3ZPmgIjtFZQyRvbbZzu783sGuR
dNM6KcQ/+QNBRNcH0WP8UTWyAUv1V3LQ5iuS82VXBqNJRe5PrBEGZHTFqTUClhvQYEooi1jKcefq
Xtdm2rtvtwPMt1wEyJj/v+bs/Ms2fL1JTqVZ6ZqSoX4KaXSyXem8r0Ug62f4hUdCM/jMxdRqspfy
inHKYax5zOBlVReQDGU4y6yH0vOG/utL1oZAI3FU1ffcuP2zrwunbtmXGAuLMqKqsEudhbEbF8fh
T9wK9AeJkpowZifocSGqGTgMFf7j9t8woAbo45rDlTBdon8wFztzMrR++Cc5m2gr7LJNb7Rq8Whb
Eh9P1EXWbto3+OJnnRRqlc5d1Sz2hqISFwpTHNPTbm5U4gJ4rMkLWlBTW/tKpaXAwa7IvAXbA0s8
4f4/53FHUv7yaaUoI/oYIcnBhg0nu6IutJdOkZwCKh9yo1/E/sc2n7+tjwPr8KSWxMCxgZk90tCt
NpjTSNn6i2rOOtpeurJTj35G0oZWtV2PtRNTaH5jhZjOt4D7uAFTYyTGBfKyPIuPMFGBPSnudFo3
ej6jqKyd9jYlF9adWuL4unfbsUJCuLjb1JNNC/0pUxFBx4ds6Fr03I1eZsvabtbCVx/0kr7oYFFE
MvC5xv5k114G6ble+sUkf5s0Fya4GqcgQsscG0TO7MWCK9Xg/w2OldARIOtdQPc+z0PSXGY2qOGN
F4Y87yVxg+IMB7DN+ZHDj98tq/RDUlBUUEvvvIMcSLIIQDuJA5nw3BIbrczVgGXDOFoZEt93VMFB
5ZXSLrQGSQiz3DG5EKCRNCRK/3PumvdLMiB2UatlzEnrZcEexKTSad5RkzI5PGI52Qy9D6P4ouzB
V3rZx9x1Bajq7T98kb3OCA8MXqKtobBNw/7Vw38pS3I1FvoLwbIXzaL7hrMmG7Bwpw+r1HXV7NJB
19vpEfOlJsNwpkrY7LLbPkimtjs9z0llrmf18RWpBvJjycgFecABK7LelnRk1GFwNhnnIAJw6kTW
6Qd4W8HTKjCs2eDUkb70UPOaVfg1+Xv7G6/jabKahdGI5s17bxBJf3pmTPBxzf9Y2WlWKNkZCQE3
X+o03qGwJsS9zXs9iIwluMNAw1Qw+6KSb8GPzpdMLBaIyNE4pHE8oatjV7W064Nxy/APhxcbX/Ny
t8I7rlqX1ir8yV5wkPWVwyJZyZSVVb0zWJS0x4QwEckHfZQU2hk5YVNaIvREeVSBIPglMSWhuJUz
xqR9botIYnz3dddtcJTZF+/NMS+umSgDwEdlcIBw+Dl9XxtSPz4sPl6hxLcu6e1YkU0Ju+LKiCZE
2d6X0PymlmQFDd2uVy1ISkGSF4fV5Yi7GiS0Ci4eM/lrd9vU6kIADq7BYE39q6LcjgjbL5yOXwfn
BIIcqhCnzOX0EpXsLJuS1hL7fSh3CBGm4ztQOVmKLU85CXzKd32RKZvgQy1cnlkSGdW4bnS7yr3w
aVW6JmlcC3sJQE5+0cPH/tfZvHksZt6h5aWuu3V37rs2/nnd+YwCeaLZQGJ59KMwGzvUrTCgr3l1
kBdkfAT+wjQzr8X8aEADcP4sdojGT/fhwkU0giX03+U09VmWy/1FuW6JsrtjKZk5+wtc4KLN5c8h
0gFB+KQ8KjdmUhl4ymWerYOtEF/yB2cMTUGv0Bf893FWDLoXqYRnQAcx6rza0HYbWTxfr+9CVp1S
kN42A3TXlb2ZFQxcz1KqM0zR4Uk62oYnADF2JzDFij6Jh7lS7dOj8wLeUNsnjt7WVF5dunBbexZi
wX7rBqaAcd4/lD9IjZLfH3zDffGVu1OBBTz9mgSblgKVgF/ZjNumiDHaFQdHLCHFWkczCIOn4cOc
T/dv6hFWU4eZSrDv9uOuW3tTuLBzIlXMmS1Xig8AsAuXLi5wL8j0GpRxcLDl2tz6flmw9jNRc7n9
09eJfXYCF/iDkt4s+j2vuZjLETnnyYTO6mDex8ScFRzp7KkRcIKyX67vlKjDc0uv+A0s8YXgT9zL
6lQFoA+y5QJFwWVIEpRic8/lcusYm2E8OldtNIp535zOhfNkqQDFTjuRG6yi8d42vL87ZbbAodxw
WMWZoymE9fkDHgToiqoKsQPzT3O5aL3866T4R+7oOdFIYuUV6QkUh2TrH9D1E9I7nzkkYT89/MYV
vaDZKKw+OquhVTf3s25mCjKIhts+CmhW7ygpAAYXxFeBk5MHkuRqZh/qsUt9mE/dP/9s8wf/6Qd3
w14iSHjpF1KcUowTW6BLomcg+agleMCS1/2or3Ny5OtbiobApsjusknq2usrTwku1QHNUtWV3q0P
RbJlquKF6ObB6fXXCxn5NrOELYdcyG5TcinWOHpdm+LQ4YhoG73iQocw23XnM8nw5zN8nM3zueZw
H5SrxImZlfc3jVrJDq2qdf6Qgq17NIwiJVcckOcUjaVzBCl10aR6pzLZJyfkeaqrVbX1VLjK0n5+
X/PlSoMJp3mA5T2XDBr8OPRc0NyfTzY0+mAOFWglixPHQL19sz/5kYm69ccwe+FzUgv3DIZ1kVjy
Uur57aUWd6MhFJIs3W3/bzPfnTS192JbfxUMSWzZdBNZfhtyUN/9z6GAsqStnv4xTm8KnrJxP0Jv
hFjTwueQMBOJk37pMOY34gQdgxl5AYIUTV4G4L5rTkBJVpYQwRZQ1FGFF1oi0br9hIajueXhoxlz
6B9jyd1nCu2QzHvrB50eI5UOzOTcGpb9pVHuKSAHpq2w+FYq+gaVyN57rFhmyC1aN6UdrLawEqbN
PrXdLnXnMASSPleMlydS2nh0L8MQAzSNUJLmumR73o27n9a80C7/hgksl/QG6J4Rp6qh0P/yHFBa
fLwYPyvLjtRtBmIClbs/+R4rX4N794Tj0u2L5RUH9bD71/u6bX5W/9gLrWt8U49tcEnP5Ma+xz3G
5PK5Vb/73xtpCotxnylCv2e/zFX1XdQIMnp1yeGuzF8eYRS8NbzMYyeR6zE+aBmaz+O/IaClutVL
2KwuSmTo9PisD96CpYRI+yP8fuXy7ygV5mZkzbCIQuvPuk4yYaaVduhSUTAVjuE0J4xosNhslSGO
eBS39DeM4ieuKiTWDS/pNW6w3j5aHBNlCdFoWBw0sxOM8jGN8qhoJE1nzyrRUOOtzd4CSGwZF6ci
QiniFub1rQvXJAH5uLwW8PClMrFyfI50oHqPDNrvBdDdJveYv2ADqamPOhq2PlIUWCrMyBX/Pq3q
izvqQ07VwGEf7DVL71p/DNQoecR9gcI8de+qKT4PpGzNMBeOfzkTnp+woW7fDyCttTGlyi3PpND8
4KaN0ZmUAreFK6q2OJX/AHyP+/jp3X7e03IH83g56MDism/aIdjnaXkeDIU/vyoshPTgTNPYmXdh
xV0ulJkDd9RB8/LC9I1W8+GriWtmyIC2Ox7VkCzD07N2Gjjq1sQ6tfhoQRDRsfrCBVrfJGsFTvlf
hFVzUW4KlL/HpCOE9vG4z8TyUKwwyWqSVAOetouySI3nmmpKZDtJ6AqJxckq6fNy/JoP9x0MKxZ+
SSfHnUkSzoXV0TnXmkHhP1gdpj2F+0Eh1XmOjK/+EVFVERXUyq7D7/2y9rvhTckjveeuKCyf/gcw
YbhBV74M1m+ub9xOQak3wuqOtnMt85og4PrUh5IYmpOWRzPgjM+yK2xSljMBXlfEET/g/DbSqxSG
7M730efqvwnU0EKGpQFxeSktYKXIG8zJmFpVkmZRaMJyeM5tA8Y9u2ddod8osDGo49QwljWSn5GN
FJyKMEGzfuZIy63L07KYPmNjFU1yN2vj/ZEuSxCckAcruNDoxZYrhNlh1ZxOotR3v9x6vPoyzJEN
ET2/C7eTGhZRNUz/17qBiH79Tqw8RVP5fgcN1pN+BnHSz/mhEHxC03MsqhAzSgWTkLQSqlFz+KRt
w+8Z5qdc+DUVGyPIFN/IRlIAGH4+eV0gpy62Rf+kOsdZupu/SKLnWBm9Epa6VVUZYI+RkYG9LwbE
UeAO1AgXiV9SF9mhl2Joilis3h2s1wzyaeczMsYkXTFdatiA+JOukbcCmaTJ4DhbUDs4KDX8oeQU
wpquf5OriW7f3zbt+48Jhoissjn7bPwSTcBBznu+8S1UiuzzILu3ZeGemaHhNh9PkZYPhI4ZKRzZ
WtmtHFDUnH76kTtG6aqNIBO1nviqLjUR2xO7vuNALfFtGRtJCULNcDMWciQGCFIXnu+i7hrDSxv3
ptkbcRTOHK3ymCp4s7CD74ziSvJIb4e6bemSJ+mlApXAMj3zh06t+n22YmjWbtWVzgkNC+GcIkGl
uf+s56BrMG7ttk9PwtO3YiliK6LTRlPwjUqzWe+7go35o5lb1AbkvWTJTCviXosld5czSAHT4kMH
BQZByR1Q1DvsQux7EiirDxPzxnJmg4S8XMEJ9hjpX+66FtJLqHyOMQ2CNuI4NMgSsYEVBbU1toqP
p3AJD2xQNfM4dFVeHyUDFjQwIFPEPrzDF05eVtYmpKDqsfXMkcmZW4RS/1dVM76pNzhQeaQ4osfW
ofD+xuVl/JdvHefglt8vOjt24b53pLOpZ8sboHxZ7DUDcyoTEcjuWToK6gvgMcjbs6p7AvvUmhhu
9S6Sj2pS7xaS4AnPyHKwneFYugVnKyGeUnkLia+gkVkAmv2KoNyU8p0dGFHTLDMrXgBhI0ol4pwV
RD9x6QOUy6eMYafHChkuz803XFnNvzJOzJG4Cx288brOPgmOPqKLrTlzG7CDp8O4fgpeHbRPfR56
E1ILwbo0Re1Ebs7LpcNf9ehJytpwii7gBk7gpCPkO7zjXXiOHPLBGD+7nCduDRFqt6Pv8jDQZU3l
2IcbEoUy4rXpMX0CMI90xZWIgFMj4lriR2nIAg4eCrhAdwNEmC2Cp5V1ruB4b6XeI/HBn5+0gUM8
WHwva5eBLCTUuKkGGip8COxUGTxzWQECMbUjlFbwtGzDZmkH7QGEIKZ52A3sHW2l+xbxgg7GJCWW
LuMXVyMD8zzF3tE3EFE4C4QFA/AcTaflEaV/omwo9wau6w9S0F3WrGeMoqyZrFjJZn2gCnPq8cfS
IfnfTGsA5wZLSTHYrPE1tFTaGVLmSPfd/dtsMvgleSqHyzisrUpaC85aaJzUd3mtEV5NLwvzCX++
1AY2hsyVuy6Jl6uFR7f3WNqynDk4s7C9SMgWcHcj5QZ/DXjvmbZSkASSAZ5pIEG+1AAtviVrv4//
rHe+XDTA1K37nHmMTh5Z+eJZKSbMsz8MzNpMUp7VbwdwUNd7j2UGJxrmwANlAqKLXmGR5/oVOPhT
ORXd+TJSJaOBQMnRR/zngeUyU7+jdHTwZ4m3xinlqHwzOHc/pBlsLSZE7ZrZg3fW6kWswmlqh+U+
xkD+5K1GJrjI9iW4F7t5ZA91tg3aj1lFyEPJ6gITZnROL4afW86+h1kmIq/acf5ulRSL/k+Xmy+P
6+uUZzwtERmOGxu8Yqx/WS81DBUMA56J8x+XNaEQ8F6OWxkHF6CXpM6vfnCbe/odHPR0jx+gtVHK
HTZfJf7HY/7OosF1kUwVXm25UT8/CC6HNMS2BDNXAPfxHcpE+Wq7I4O/brvQR6qXqwSHzYgKlr6I
YGgMZa1b5CZgs7P2vaT+RVXjyo/Un5YEqpq5BHMKGMbk0XcIt6uCYPAjB7Y3/itj3WbgOFiYFRzg
lfyPfh7NZLgoWqoh89fBuvs+75VekfzFvKynjWMKmrgZ2zvkCM59k96OU3/NWt5d5AL+t+w1/F3T
e807wzM/vwFMmgzozAR/6tLnKtWATgEn5s26Eqn3q2tzwu1/E3bO92Gb4seeR0dm5y44CA2MQH9/
XNXqsxrehH9L4rpvuKU1Fe6+QSo3g7v/NLezxVgPudiY1VGcy64kvmT0A+7fauYrpjUqvw0QKwhW
CIc08EbezpAUQiLCyq4xqKbelVFUP+VSjkdeNT6SGTMCrtcQrRsvrmNeYUb8U9GbalU5vrqx5+bL
0Fgx+YUArwrZEtYg0vj4sDFVYMh/KUsn4vakCdHnuyD1lUxYCJdGdzu28Ga8vE/qO5ImyLfrt33s
BEpSNUrCTt9p3i++KhhUj/Foi8o5i54eOLpupXROrGS3OipmOLSxAJPav3j1bMKabyuLy+yTp3vL
swZ7KsiVZwd5+HEbZm9W+hk3sCkA+DlYpP/lUmCpGk4Jj0ktUBWrPnp8SKQ8m5hV9tbBESjtxRZ5
0UydBXFRPLWScAkuQHLTcQFNSNsXA/g/rzeMKzn/ivyN02j/YVd5blNgKj3j54OZzuMS6ZEzXsSr
zsKQpnRsGgU/22MuMf1l0NdZEHcLR8gh5uUrmqnECqjUmZe+Tg0A7H3wHQvNAGmMiVjTMxyhHGNX
O001W/3eps3uHx8/tpJD1t9uphudwh/Og/z/ed+TxunmFip3P+/oVtEAV0iIovBGuBblkoNC/HPS
Rgh7G2Ar8XwsAAz9cQOvcS2RoQkGRXmBzLVlPgCKPLYqco41Iy/5lYgfZtY8FI8fr+7DaGyTgIUZ
HFOaxmvB9KMuEggoF//vPy4CdNYME6DtKEq8oE7ahQrG9tDzSh+nmc6CrbJOP8/d0D+nDW5AWUN+
RU6/aLCVGkVPPDS3twg1LVrITua2Ir0+mogNjmYcQmWN/vi+livJ67s6+yzu+cWZFlZJRZdJPwwu
x4DWtOWwAAAHFH4ItUhwLPdwY2D3RzFvyD00ThqxxHHXaylXFHmLbhdAJzLJF8Tfbf1slBxTyWbV
1hgCFzOeJr7WxP0GFWfIVhDd1g43zacrT2/GYbIiPyJZt2lG2KNgrMj6SfLpz4I8FFcGYK7DH5m1
pFnlHM3pAx9Y1WJWJy21HIYXEGHr1wAGaLzS/2hf5OlZIgqagLsqB81T8HjWqc3+Q9d+YiEJTG6a
FhRGbl+9xu0yPEZ/RUS9aqvgxHG+GZDxUwJJiKsAd86SnFV+FN2iDBe0Sdv/JeVLwWE4qexRrZVv
0RbSBZ2LgqrGoP6AMuOYAEUR1MQDLciIggsGC5fmtvQUsXqWunDREai3L2b0njIFeBNUpJdKLtQ0
jW8Iw5Gei2VcbsR5XNLumDTGk/OJzqITPk3lRnG2/zPf1XLMrjvU8vxFasMK6wUqGLkxw/ZDkPBu
ossxUzkNDK58bhjEil1T0sd/Qwb6lCTcqzF8nwisej90X0CO266Huns+EhrqMbawqy+/sL3dIuKP
aq1M39dajPYKSe6SGX3g2Ukmav9IgdwlDu1k8+rX7nSHzU8XwW+7wDjoSsiGylCYhYqFKNe7Idbp
bt2/43TL2H6Blg/xbQeYTLEBedIrJucPzlXGNi7gUBzMvwnBBrfRxnHG+EPgxNK6oBcFyx6DCsfr
BI9p4tmJqb8JdJlC15LnMWrYBFPmIrbFh5SNT2dNzfGZJY+bkL8TCT1CxSvwS5dphdQF03z+ewj5
bNowRfSJTflikYI5PfbofifnDs+9ZSTvcsNfBK6eArgDmEyspG55uwvjpDiW1DUQYsrrT2R3qYea
SPH32W+QvG05IOi9ABURuHl4guExpC/hZ15f23Znz0/K1KhBz5PGdk6us4F6QlAbYngoA40IP482
av8QZiYMYlvN7lf1KUl0KDQ5Oxp7JMdg2F1ZEhP0YmDaEpvvT7xycJWLT+vgWErjl2XN1V0NmrmY
Wg8Ig+FDY1i9Pvn4O90yDhpYyMh6OmQifILJ0W/SsqM22AnG5/JWieDDI3v1OuHS8M0wfD9eAV0P
oU04a+eQI7ue+HoPv3xny3Pb6p15SafhBdpdcC7d8hV3r7VwURrwpKGc/ct/KHPnmiz5aYhAGJ8T
tChVA67n8zYxMQXnmHDObX2siIMCaaFWZAApn8w1URixW7xS1DcUNgGo668shPT0G4XXjxZI34Zs
eF6FB3RxRw6Hm59RLTlNcKPUvt3okuHNbfMvrLPc+xthfV6NMdNuEfbRWb9GudyHzt32jYQ4wc0z
IjBH+X/Xd1ZebrUKnCe1wH7UsxuyjTCktTRvtg6b9gzWc9OMRjC8sOr8OTEYvKyp4EzHfbjmSMJD
YsJV9KVEwV28Va7PyFIyx4mu/F+hPyVrdMXerNxJ90S2vXPubHx998A3wVVbZku4R2bmcR0lucyh
V3rEh5GtWrNRPHmy/6RH490NNgnrFptpyY8E9Z9bGU/2VZhz7MJMieZ0BEYghQSCYLOHvsilTZ8q
tqF1jq9VhzBOqMnBSZRzXnHE/+ff7S5hld5gDbn/jB5vbtJgE2I6aBHjm1BQ3UAB0YtqkOhhT8KD
MS3zswR7ZXt+lrrlEoDKr57mSTFaDH4cnEu9SKDrS324sfMi8Bv20C4zdrP21Vs0P1POAeWq4RdY
lTV3WLT0uPGLVOsQLV43oykY3vlKMxHPCSec/MVw/rrInMCdZCbxYOoAH2Z+PLqD5SYDOpTV7Nqh
j1E1N7KQrdJPy43OovIGLi1FrJ8Mv53a9FCMb0TUQpUH7c7dzBoueHvbuN8JjksCForlrMqUsFmm
p2VFRVUqm6Wc+kNjtPjCxRjqJPC5dY83qS9pyTD+uDuI0uWVD6WrbHtuQTaFgR9Ep/FbIsRLigf8
eTLy9GUHcXgQ2hEkc/OWd4x4Fc2HTdwDS+Kf2ukloY03tGK0pkjS02oZLxtfpgk5EGI6SjJ09GBP
ZulYHn5HueJU65sa3xRjJYlQELi44jXVSu7/t+5FbZEyc2ptbCpjGTa1N0o2nSbYZpUYxJ5y2c5c
o7Xcu6o+AMQhsGglsgSU8NGRCZukOAtRhX/Du4QJCJeOjmwbRGUOssAa8CAonXsjdHFWmYCpeonQ
DMslK60PzobNTd/OKYcqnEaib0WCURqdv7vTEziMdRGhIAx0FeXksG9DZ7q79yQhC1bv7/Q6GMsh
ZUTPB5/F4tYBsMz7vNWCiJR4jwzaHD+oo9V81lDPsuBtVbZdtfmxvZFKdfFHs6UmmJ5ZnmnhUmMI
Rkx3tLscIwt8OjCTG48U7WmFR9qSv1K1kdUT500b8EeJ02WmompT2mQqkwcn3GIrzIcDGxMcnSJW
clVZHFk4yx3A9QvOqiDcdXqlAaQLVpsFTvLS7dLqabLE5ykn5YU0wJZR3kgd9rYfyJwoevMn9aR8
ew9c6o9MCPZHYIHVMAmM9pLcfOtkUAW4lXI2/VoWLn3GCAkfhf0I1xkJB9/Su1yJBcgZ0pATxPSH
ie3UbI9v7oOnGmWc3nHAdM6kFIF2xZDywHtxpI7oHjUsPn4TSUqSPRYLV8ZMBR3QdpQD6v1UU0Gj
SAImXtjCBq4wrp1DEFspDnP8rjpTr3swUoHZE55FoxTRRblDk5vjlefPpThBdjDe019DnRzCIzgO
mvUNhHyFkA35ACm3MeV5Nt1wCvmZpUjye0H48MVAy/i/N+xQQuxSH0QRLy+aAiXBjtlWppgIBIq+
jDT/eK29RXu1PIgk7Rk0+SqVKEBDpa9HXXKYDFzct6id1fB3EfT203dt8gDnFC7GUZTqXz6nbfPh
aZs+l0eWxg7YKO/rPAiZPLd312BTzVVIwjQJ+utWOtO4NgXqWpbjF3dbOJAs7dyuRpj7FxkEvfdw
oNq0w7pw+K0PQMwZ9si3EX5cgZxZn4F0H9kJe+vjlUKdTLjj/dKmFJGteSiDQ4xnWcvpbxs2Tpuh
jT8BaC/8yQ2xBAKIzVxYf/LZ83Z3RSI8T6sGym9Qpz6GvzSBgXk15Mx7lXz6pjCX7CiPxMjjNs1v
iOqCV5LFVJzXVFtYTulq/FqETl7Qo7D6+Z8lbZNMbRovdkfUb8PCWDoT1TuxM8Q3g8KoRwr4Ja0r
uCkqJb9L2KoWBM/dv5/tlGfoGHWE0l5yqq0wZdgOS3UEnolJ0x21VcqYXDvXwjxsjXv1xuyewR0+
mNpafQQXOZpW8pisWiLH1M8h52/SRP7h1tsoQQRQjWkPgddDuydLxSr7SKKalxJ1csBKcpSi6xhJ
oyJ82bUNOoeovX9V7KFZEncf35QJL20HrI/NBmeL3qXS9W6MNAfxR9Z7lClgxYM86DxMv6nKVa3H
CBl8mKM6RF8QO8/GgZw+Bs906MAHgkTNTy8T/iAWRYP/61fq0DDxIT5ZhhQOptOwl+gbPjJYldKz
nGE0B+BkMHV4uRoILmITQ6ucmNpZLrFTJ+fKQ22pMgNca2fGqFbaWwHbNu/CQjZXYTpe/UCe/WAq
Y1M9AJJ8eH8pjH6hWPXRVfrfnKn8f3KA5EPM8sJh1F73QtP9IIIZQG0K2np4WbGPMjXrWU6+JMZP
BWiMM6CMbsmgzu7ex6anXfIpWsG9iecVBg0EM4gZUzK9OFnibvc9JgT0/i3PvGVjrWBvQqjufDNd
wm6ixjDosTV21MDop5XOTka9Fm13BCZCOnEY7JC98TtqXwN5OUt6cJapGN4iGLD77HntMcLHSU/p
7kmuqskzpuIfd2+Df/V3+hyQB02+sAuevcHxgrXLQVmxySKEi79JOad0t+Zit7cLAcVcHjxV2qNH
AFoiySPwb+rQKwtBO5ta2DctsRdnOW2vwbsQHuwYp60Nk5fP86VOG2XAPQwAG1dF5L8zyvgqx3zZ
aY/1j1F6/Acv48xhcA3tPsm3VBLLg1LdByj+y5Gn0yfGDoJg86DkTLPczQLBWeyZLbjKBS72z9I6
lDfLM7KOf6eEX9C3SHeLq34qOjDBovz2Kgfic6a4qFJBOD19B58/9klZ0TAlndZpOeA5CLiX5ADh
azJO3Iw/VhEahcOlgMRcyPfRSoA0Tujg+HQpgd22U/87xjRO2AA4akEwPpdkalk5ICiM64BOJtxp
bum4deJ3nFYip/n13dni+lEDd7PQSCEuQxYIj/n4qGlvndrsnzPj2HBzzwqO9BU6YIPx7ZWXDjXl
mWd8PgW3K10AyxOPlTqbGGaT3kxXFCqm4hFMp6Q2fyBymt2IB0RpsnfVusP14DHr4l1QBbLrupNk
xNt6rnu6SrVtUh2d3Dq5RD7FKKnGY6iDfIPzOuRPmEC3ov3CTCKY7C46QNnHVx62vjcyt7FrjUIc
Eq0+z1W7QIumE/IqeEXZC8E++T8EnV7DFXqiWIZmF3DoGf/G6stUNXLR9XjUTW1Ndo/o+Guil2FZ
myCScY+wqNT+Xxz5hG7IF++Dsf6PZNDn78KEIi8E2zKV3gJ3twgzuefcOU8klip1gfuFE00DkQEb
DR27mv/rmnfBmlVcF/wXUlHXedPq7lPDFqJnszmMZvX+UfNxOikSpEQfyE+ExT9PGM2cZpv7+/fk
waz7bHtZGMplhux3FobPgkmTto8m+Xg5p1taiFeaim2QeE+SHFbDWoJcQFa5tyqLLFNjuF3xFdrx
v9wGHuym94yeixYn1TjIMz6V9wxiG75OafxmiYjfbzxsk1uFgCOLc9pkHcw1i6ZihFk3GcPFZA+S
UlcUBIkhL9KgPJF/4yAFg80tlfsyC8v73W6xf6z7MqiKZOtYZrNDNoiP6+wUEGLF9UDZ2s86fbif
JimSn1y21yyY6pTWgEdVEMny3UwolhBsFDp4k3HSqDmGltjpijVv7OR/1Q4+X+z6mmlZr7QRvDo4
19hAGQyDWC0ppyWBDW0GzvEDoQKmtLDeSYAbFb1GTRM/90rUbDv1AZVqwv+Z4vCGfh4cRhEqrZwJ
ac9/YrBhGlU4rxzRwNQhcOvLXLUuzG5PSc/babvt7smAl4fkytdzWFH9fcjjPFMxwPDBomqWMh4N
XghuRgfXcPbQ7jrX/YKmVoZh/TJkOUKMkm2uaeho2rmQrpD2fYiqOafJNrwtSY5BHR9hbepME+YX
psqpbCs3e6QhcyvchniQaLmYN/eBV1Za4/1DP62wzcCfgY473fuaItC5kcJoR23hcaWUCaJKMHNB
MtBmqfj1l9n9WTQBQ3g+oLhs8iAoAK0Wux+vk6Ab57J1HzLpnsfI6rFod9+S0oZ16yulNDcwPa2n
5N2LkARsBwLqj50mDFlrl10S6eC2R2WmmGsSbEPu4257We6Z1PTA+avAet4DydslFUsrFFKeoQAT
VHxDX4oBgefUxllethtm7TUr0+nPS7OBYF98FU7nTTmAG7V/CD2n2qt+/mVUF1J3utwr5DRvIImV
nSsX/xaRjXvBQ1qs5kPrBK2Ss3yphw2Hugedn1Isrqw+wkMSuZoxUfWMLZvCO8DryyudxAEG5Mru
EcxRdC7uN3P9m54jEk5zK8fEX40M41/FHyOM6MniPfQpgZxy2oXge1Z6aV62SMJZDTgLlnJZkgWh
E2VwirLLhna2dFITy+AxIWQy1WjMUCeh3zWtGNduuUfKBoDN+fEmvfiPxN1ACCrBVACubAwT8W2o
3bwcY1FSXuCTv2HhmE/jo4LlP0Aw9tFCcsu/cZo/DjRVw95s5c6Z9GEMXw0M/i8sCBLFCaJuzaLG
Ap3gd4+iAR3O/8/5vJsLBXcprNlrBfLSDHV2ut7VbeBkR06XaLbaF8VZTLIBsJLp0pvBd+P9sCMm
32JYIaOh8SCHzheAocRSkvLQZtS5UoIDdy7C97G1rnr+Usjd2s1kIP81bQPrwIh9eoSL8tCHPqn8
W/34B3wyDggjq7HUG2H1YA8hdjPwnMUxuBhCt8lrOaSrT/kupi84Rl4WsmvXxb4g6GsVB8DshIK7
8ClMmrfvL3SRUEw67K440p4ryQv9iAxGx9RZ2YP2APTpWXjy4mSMBWEPnwNKvjAW/LTJ0gz3SadX
WzeCmHOE8/YjfdIR1U1X8TLPggOwSGVSvlvG6nzVoUzfrsk2akHOQj9kJBtWF41+o3mcM0y1OBqB
0sJg8+lVoLUIjrjht1Q1tFPhTXxgarvrrHTPSjLQZTKLo6XoT7guyGz1R3sf1MfCnSloJ3y5t7Z7
cyJ4ewwzMR2EU0qYWwv8ulWN+Zydccflw0t1RBlk++DaMAfvYp6/kApI5c2linDpxe54CfCt4lDU
ljYw7U/y2heDxH98wdRRuEp537zU7oNNlcbgdUb1QoEe+YeLwmhgfhhoEK7vpzLZq5jdZRJ5cGbr
xYQN9gTaq2URYE0NE1vJQNTWR9cIlV4Zt4pMqZN+2y/tbLc4goMvgTMep29TtFO47i7mpYk9ye5f
tPz7WpW95C1/87eW03pAr9gTKS7QnoKFZ45W3y0DdsqlaWqBN862hWWxLe3V7aY6r/eMbV3a75H5
/sKhNKfOjUA+gf0CkneBuefb05z9gZZH/AeL8aFOrOgUSLYHEE8ceV5xp3Euf32dg5nYz2Dcd9/Q
c82bRE/2CLYE7xNLgRVHT10L02udQas0Urs/KKdRhqiOiKkWURchtUm2qaJrX+e50oBb12JDuF9C
aGpq4I57uvqqLEIeAu0biZzeFa1lf0yGl2LUDqwk/v8JgqTbpNcQABABZsQraFLdmqlp4y4r5Z3z
zqGB3vl8JobWMVJPjXL9+/vxZuCt6/wVHbqP858ZOVUXRYtcoNWV2GtS1t2F3X7WL6KWN2pf7SYN
59IW8nMPYcPfS4k20kLcNHmZiqkSsQoKRyeCq+EyOuGwLksOwUYqzq3geQcSUu7BPDhE0q6uzYoZ
OeTkiWuvtgxEIRlqNYK51Boea18IYZbzPxRASvzTHMffhqNoq/ewb4bfSjWwU4akJp91kp5IbPbQ
pJTbqQK50icmcxeQwBvv4EeBAfEx7OkdGItQ8++duKPGADCExcQkeQ7SCCnFgG3FLYXOwNexdEjx
5sR18rLJctd6TZob9q2Nex3ZQxliwMMJ8dNHOsJp+TJ0ln/7mWJKDX8mmUGm/mvyyPxniaxJv/JA
jW+I7RNaAdoPcSBdtBJ18sM+PFrJghBz5xb6UDnnr2CYzD21YHIOVPgZZD8lp7u2ReGmZaGOFUzR
1RO4Nrh++zQarUxKTUYL/XmtxZVTugOHRkwIqeHvUn7Q/S7lO5uIFT4bhzX3cRuHajc0478bQMr4
SW5Nn5CtqcnrjjTXtsXqzjmS5l/TGJbsr9g/3nKyZVr1BnxNJ0lZkD3w47r5tbU3NmQXrZR56+dm
292MIBQ5wNnGIa7dMlL8ukHr13FdV2zEkxghpuLkgmTT4dTHrt0WnqLqA1FmOaX1XVbsABKXJ5B+
1ODO2ujT0I5dTNgTs2o6h0DoCi37FTgYosnqX/CXrDdFXPg2plBgH7HQ95+1zbZstz7jpP7GUXJ8
bNFloj7hO6+G+jg/K+F6kcCV4ZxiE9wvi8UImPzkePI4dC6QJXY35aPuFH8TgkyWHQy9xjuGYOjE
BI0nwggivSGmHyvn+NFYNTHSiHbQQoWno3qgwvVOtYpcbc1zjfiHnRqL/4hxKPkXooBU4mN5Zohy
jUmQiu1E+/Fbqda472Io+aZoOvsxyNikQvMbG9uc5oiNLFq9Dd4JaIoNhNOKN6Qbcy+CUzg/071Z
/XR4lrxnif5fYqpgf2n8Ns0tDyXoC1gqQCfOmhlo/VbGlb+VXPMt44a5/ysX36SwW+F0AXXZw241
HaLGjgwdpcO/PeRNVOM5dhrgE5EFYIN/HsdPwjZMUyJdA8N0jnQhlBR2OfvrwVYB7e+j9L0zboo0
Ocgmq9U+9I8AetiLCuCK7jRhDz8v+RodeRcQVBSizPjy+zsz3j34gVlM4SxyM2vWW2gWUlHWvxa9
6QYBsg/kyROXARpyOpCmMCEFSTD1dvY50q+oddWrtg/HroAmaFHyImoWITrOQa3625B0a70agtXs
GWndqHlEpQExx4DRBzCsekNs/+4uZeyE0/np8Tag+VP98868YFFueDdznzLcCru8RXz1GTBz0evG
WsJ/rGblz4nLJX8EAWWDZR9cGWp8MDrmoyn1jrxm7/rm6qCS3cR4YtQaaXV3f+ckXKOJhCTrabkx
9Zsdik6/4hyvNA7aZ4CEeVf9WPj5wCdClBTZFqP+QxE9S9MuLm1teT34qlXsrlvWDfj1l7zpZKJU
+obfiljlfl3HtNBVp9r+mMeY9TVcEyLeInHwQqaFaIty+Xw/XU5RA2QJKSseiuEew5w3v/9sUesO
ocSCv4vH6Qbnsxhgmd5uevAP25uVqB4vMaYtliiIKAvSEjgQEegdPgIiUN4IvqFsUHnbNnIN0Zrs
FHnlitV38zE9XwJS2tVwfNx4eTf8lyw4RLlPp7pIdGYN4UEl3z2TkcFI+UZfrzPKy02N11pXmLwa
juRQkFgyFpYpCG1ysFtbnzbNhM7m6t2mm8nPTbffvozMdzd+fEKlBsXS0EmklAYET452ZnBUfR+y
nIdtks3KeBfRLmp1JNWQw4aktTCKat4yURBHjovy6kCsOtwEmnURFFz21Q1YhVTvU5b9vgBdRUB2
jy4rdm1xaFqmhwVExmh8nUHGBcGRbfvc9Nw6rcjN4F0V8rDry+qzqX99Lv25j3++wVy6VevMy4iU
0OHSCFNEpNDa4WvRcFPtcKYuTv83BykhsDFlflCIh8G+URHHgqYwaibHwDCLKY42dnralViK+jP7
XxPurqOP0/psuAVvsouB1uhEDk/lIC60WFu1JamhptBKLnTl/rSuC9sFltJM2owm7GX3OzEo9hDd
vmsALGgBognxix9XswwQb2A5vPWR4AAmYpHeDtJ79Wd657bJYKVHudK65QTjsnoQs9h4IROgn7Pr
ZhBlKZ0UjqTPAsbylgj4QVZ/qjDRGs/b58xs5XpVXJBBgg1Yx4hvxuni4E9Bv32NoR7qgCAlpgkY
GmEMt2+mCtSe3gfJRpQiKuUOf1TysPnI2cgeaW8wwzH665ErHvQmOgYrHBo7Brx9YzTXk98QThUj
QIyY42TeNkEXtYRHbMimyz2+dC8P7hu1edc+if3gPRMKWAooCcc2Lgqv6d0a6JKmodTgOqrSR/kJ
Ykn2b69/dIZCHBK6oYShy5zQI4Wew6+Oaxg0eDfYU0o1qbFQWkk0qlISrUWL+kOtghPQ67yyIS2m
mngZFhagzd6iWz43lGpEtF6Hr4FlKNrWLuh/u+tP80bawM/yOyc6fUy+h1yFVt82yS7JNSl0ckVR
cwdWwhKDWYLl7foSNbanin+hgWOzHR5WKGkcRph2DKjcpcEUPZgqXiN8zw/VfuxVVSoaYNFJt8mZ
K4/2BJf0jbfac3nQMyrTb1hYZjrL/PYqp22LkzkoRdGR2+A4AzZZXxtFaAgWvfkU/BHuLdTIVYL+
e/XhXlb1I52EFAAWcjleYcjLm0bIAgQo4MbRTQQg1Y1UlWjE8pkPOzefg2rbbvIsXyPnVjDXFKn1
ut5jmlLagTFW2Qbujou6/m/27cAKXL3h79/zV2+3j73wYQZqId75u3p1IGcXayqhfBhRx1Oy2BlS
yLE+eB1XR6uqelsLab8qifP93DepIphEMQUiDAMmMsilXLxVSJ448Df2NaQZjaebFStbvY0P2/r7
d1QuZkbHb80nP+cByRonmnc0REKYZAeU84+fyUkcT9PB2DWkwdSGq4ye1G5lyDRpOG+gKQetDATF
d7P0nN7IReHQq5Q8RbOh3+yuqgeakJCQVtJH1tqEJDtSJCpRv6Xm4Xdjv11erHK4esd25Flo9+/0
UpM39rxseSSbztFN3DmCzWp1qQMtHlD/h4N2SNFYKX6mx4drbWIzOVZUbR2Po3b2VtXZeuQ3hNhR
qMixqq6xEO0rkO+OafNpdN9Qjrz8ttEENPlCoMw3TobmROl3ldrzWlM2q7QvL2PnythTYznkb26S
Iks9SjwHhOk+YyNicXqJvr92hyOZThGjcHY8KsvdP/N0VglmJFTIRg2ZckpLSHZVrpAqjkf5N7l6
kYb629s/3zUOvy9mfmZeG3smZum6o+fuTrTP0wq8Dp3sMaUjZUc6p2UsFbW9xS5zBAwjbyNO86a2
Y3s+q/oFQU4LeT0kgZOom+IAHRisxl+y86hesBUqTAZBtXoLNVEJnW98pAIUF5+J1+L4ZRscmrYa
ClwsOyht1JOho9mDU1673IMWShOhlYTZEiEPkFm5/Pz+P5h/koMz1QzJBAQnrp3hRoTNfh8yfEks
rtmnmKSAsGsYjdOV/EFAkIkfeHwQkcM1Iv/gRZorVoxwe/SvXRSu+TKOoQe4GDXAC7d5GdLNy/k0
fc/UKjkOrjvS+XUF3yGbuFl86ZT4Fgj5oSofxU87BxLjNcBMTqRNI/94G3rVJM0ZoXd/H/5yy+Mb
7D4btGVTqDtcCFBmL408shiXDuGNmz0539y8oSa8G5RmdTZTzySRC1UUuoD+RL3WXbjH+P+gBk5c
CIxOH1j4Z6J0V3aGZxbjA85Bpjdk8zaBmB4XvE/xk1hW7TF7vCNbYOBZIS9yKvuv4gPgLWQTAKpC
9t86tZ7EQOu8gHqtqzp1DICeM0WWMit+piphQ18idXMjS7i/sS5Lm9bp3Q4mnOKjHgwAfLjgrH1f
b5HPfqHeYCUzZITKbTMWzY2nC1dimoyWrP8eAl0AHIpa5KlaM+9e1XdO+un6AuXjx5A1dyzx1Mq8
qRjX6v+H4qru6J2r/R0ItHSWNqIRCxQTpW6/ZaBQHrin3hbSFeRogbSbQWTcLbcZ5Ni6qjfCfgIy
DWGFNqezLmcOFLPcL/ZSHFtiyk0NVQDS8XwgeAlIAMpaQNUvp8Xm9blg4lNRLiOyctBfZ9DQ+dBe
xDezpek8LZvJSzhbJzf3vKjsCcZxBneD4ucNgbuvmEVyko5oqMh77qbb0gOjBtv9W7k4MNfDdrbw
uHkoNBcdqZH7CujZMghIBNLCODRAC6ltlK+ETGYdsUbv8zgnLbibfAdklmFBBCcpDpMHgFqacilK
Em+hW4cBZcuNOrnV9cxEwc4M0EmoQQKH5rodPPDZgMbklDczDUvPBNYYtZGhqQoY0pVAF4/Kyt25
oIB1Gdh1XBSa2O866m0IsAfhFrGA09dyqGREJXaHs0AVvhQs7k3ltfVr01HABc3xdgJ3I1nP0h3q
tVZiOukZ8mI2HRlDoaWQ0VL4sF1QzKgmcjYxSKFA+9hXYrB7Sq1lgsf7LCMTPeD/v5/lkiXY+SDo
UBSwDfKY1lekrUq+PfxiHsoZ0Yu9ZR54g1lqeUj8jnkXQ8Scy+Mvvr/w/jNz97NNKfrkIOxjgexd
igfpijioDaWk+pQluOy12kt1WqaHx3wKOT9/mku7/+7h9JbcbWHUTQPsqc32nhhthKc34PYQ+LFQ
pfZ7pqwhom7Pz4non0qzg+v15IlChwAD10VLNxBx09NWHlpVWu6pKm07c08oauWxJgtmf8QWCWja
Rp115rWSiea/5nQLAAiaprshtZ22GNq6PFs+qAbwm00HtptUzmUpnSzIDqoD8E6C0YvoyzEsn3Gw
qKovA4oRSUgS34fQ8C2ZEt5QDjXUkrbV7KWAbyswMk7dZgbnykxrGi0TvuQeWCmLYmo+D3UvELx9
dSi2f67HEaIfdZq4u5PUDNkWMdWcpsT/zjREuH54SJI06iUB1WCuTAOhC1OXhb4YSj6oHvR/xcaY
llEVJA8IXbYBgp4VQgqrmFev6suN8UUrMHDe5ZCpQ7VnVSTpoPl4BE7qshjttfSJIb1ikBiWBrJ4
A00UNNqg9NC8ksvzeTESCSGB64b38UpFEZiEUf7x/iFh+l8FuheW7F2qu7O8xa1q4wa2igkoCWXV
PdHtcGgJ/w05YD7vC9QqAJlrXFlpqsyvFcaMvGidJCukkctZ+D2gJp+trxyxAuceNvN5uZ8ZmFtI
u44ImLLvc6aQrKYGR2ucAgqJqxQTESKPRVJH9YgApYJ1+r8t7vlZM333gJB/AspK+HEnc4Nzu2Um
yZIWFVLhHruOf1htHCo2l+GfQ/LIwTH4xRuMjtsBzoB5NIUcuuH9TzKahFA5/hcWl5qWSdO/g53l
oOJVW6VGqdLJQDjbtEyRNpSCz+LKcS4916KSWdyYqkSTDE35hpD5LrCIGVplQoIjJJ9ALkv0i0pd
IwPRQ9qwU3MfADDgYuXHVQzgUimXP1OkcAgkfYqydvSpRc58KeuTRlHLjQmSXuK7rpW4ztKUSWW3
zo05390FK0D1lKMNa1LTkutg+a0+/fR3WxX3AHH632ptNLt24P6/6nt6jRxiueyVtSXe27xLK/y7
7r9dz+lbwrvMJRD1amO+DGo0Y3eYfaOMZEFEHr3e7J0rAaN3GxCMJCbdJbHrQ//6WQLI+PyCWaRt
D1vpayN19ET5DmPVZBFCHait/bqAkQh+6scHO3oLGnsee14lyFb0ClnQQAMmeUre40cWzBo13SEv
tr346NS/av4Ouz+phDVwueYK1/cREhZepx2OsCEFjo87G9xZDiweRberLvxlWHKTQ0en3YAQMQRi
AGa7nU3IFUJWV/B86I/eoM9HbVDE+JP66jYjYE3JJN3aOlpOga5qMXRzUh8DkokaeUQp1OOZODOe
LSpBioG56rFtVl+SvVwM9i4S9x0iyIS0RfJu3Ftg2PeH71UL7Da5zPmCllxTxDece3gnqrZUKjAf
1rUYu7VCS9GKD2bFheczN+TCjVCfpc1/sjGzu4c+S9R447Dg9vngJMZjgcTImWlgGTSq9Lch04jM
VjDueIvgxdottLx/L0xFT9KuX81k4uVIQsFX1dqp8s/iQjuIPKVnAp1HUeTCzzGPU/uMvyGYDSGA
gDzBNTGWP1//Q+2oBt+8yKkOoMemQPXJplB5ZCZm9g9n2dOQa7VgPFjXc0DcTNkNHnShMF9iFYu+
sfoUftSiQoJnSLH8J+3ZhPNhgZM9DHaLyu7avr6nRY7MkPS317p0aHfrtDF/m+f8dQCYfstiYtZC
vXP/rH3hbP6A9fci2ZubMETiFKN4GSU7QRHnlOUv2hADUjpR0tf/GTL7plrT2dnwl/cRWihfal7P
P6e3cKvkjcAzs02B9wC4NyvAs/F3YTxTC/m6du1xZKweJDL3zU26dftjj3XSjdjr0Y38TKEFg7q8
iyidHKI5hdM9oSK3kMlr4RBgkEeCkaYpOcaZ3oe4vN6DfVDf/Y/dqVawE43jlYz2lBs1JreearAw
9RbzGzIgAtjtYNWtbyslD98Y+HDgompMJgxpf5SO3dMibeof0h/HfkE5RgZHMFoc5xqaAEB59QtY
UvItvTkvXPEVEdHy6mhLlS4Yl3+i571g692fhGzwuZ+V2PFmtDO0lCCSKqnBTxT9Cl4vq2MVfSy7
XXLg/o5i3tI+180j6s+9WOD32MxX/1Dh5jN1zGyOZGpnwzKE+rnRXhQ2KFKie3pBTDovDq7Iu4Xj
ofvYI8qseK5HSk//tHMYLcIGXs2+IIiJ1O5ZikGM1o0RWM70oyRaq4AzFqVbFUePgKmxJ4cYpLDD
0ztXQKdZm5ZsSnfXStp1KQk9rBnu0Q/ho/4LsvGA7Pq2+GWT4Y/QfZ6dvHn4oMzu7uv/tEuGOm/M
shrL9uNa/wH/OsfsPRIu5yHSKVtSOjoPT8BhbmPlxvB35RkvU6DDtS4Ec+zIk36uctaCruiRgLz2
uWTagTfjxLqde2kMxOi+yf71FaI6FYqUOVhZGuoWW0bXcs1y1rzl+fUM/y1dc+UoTbXc8Op1j5Xy
IEXlLFINvwaC585MrRnANiblRiU8Ra2CMfmXANMnKad4M1YJ75x8G2iMfnJOpHT50/8VeKWAaaLX
SCTqCJNhDE+BXceGS2yCO7/S4aE5zenw1WrjcopeZaKFvCnTBQkLNHtMA6NinnkaKRE8EywzZvW2
R30iz1ts5toTnTU4gmijQDZKy3ru3aB57fTkRBvp2NGLYKR7+tZN+Nm10DSERqnsTmB8vzdHAMh9
TOG/j9c8M2E8y/0hxddOZ+IP3DsZrL++R1Hd8MXFcV6JBOXu/d1ksDxOdfE9+zcnxg2igUMtrdhr
XfkfshSEvIA4xzhqOa/Z/flCISoqlyvKu5PNhhuUtT736UKwBlEWRW7M0XRE0km6EtBalkQH6+r+
8wHBHXs1yymexPNe0qGydMkuv4sdUsgyROf8yILzlGm5PfganHEQPZ1xgoK+ynuS1ijx0uBWoWuZ
54Jp/Gt2axMjyK5TFgjpurpNTex1hNAfTbL63Ge8fsYdBPufhy8NhuGZoo2xa8ooAUsdoFbDjnVO
AjGkgf5JU8JQAIXA8BZBQtlNsOF4r81SD74tt4tWZT4DMF9i40Q/s+UkA1MlTzi6/By/YDwFhhK1
esmvhfDlGPA9o5JEILXHgULH3pVNaZ7ZUwp2DM1SKTzUgDEpvUzXXa2fI9+uf5dt8u4B4ccPrk43
FLr6MXn+o10smWgJiUv7wvqkFOYTP3Fg0HMIkjn3zCTa4vUm5PLciMS+LcvBAlUW+74nsXcdGPJX
zuGSoxF6RmHKHCMCaPGbR3nVxieTRq4DTUvaw7Yc0BECUKjRgzG/5KTWHCkcWmOUWgGWwKvtgVxX
ThbFlLp9J4rujp39VzWpJM8ytTGAGfmhRImq+c4J4OuZANv/BQL7zH9PIIg9u3pGhJWAAIt2N8lr
U/YAyetieaBBCdY02Gh1GCN7PvUSVdHi2Pkxwbhrkg58ZVwWF8Qez2L9gymSUm7QoFk+POxiOBP8
eMyN762Tfns0IAzQ2jYfs60tCAsWm/w6qWPXW2+4cVzhI0xFIm70zkYGa4J89G4o6OVITeO5PlVJ
dnVBKoney7Y0QrSfacjHmTQSqXX1s4gSnRS4Un2E1zziCx21SLE8pNWC9ccIM1udZThdY6NzhwS9
MJJw5OT9LpBgI4D3frWO83M1AR7hUcOvfvyDBbPl1uNHH9y/feGAL3B4LhgNtm3sd5hms81gpilK
qUN61//bU0WRODSR3AeNTMblVTDQVnrh4Z9WQg58eymbQkinfB4JVjJssAv3ljw+hYvaCbQQyIAU
WQiLKGvMNWY1i4XhJ4HESLI0RiFOBEQBHGX6SxZBeTt9EarzUOfoze8Z+x/BU4XwaB2MFUPKMXw7
rQdwrh2j714NBXizGfoe223j+d6T7Cai+Y+HrgL69Rey6EgqU0eKvvXnCGguI76lPfibpT+zsqw7
9cjdPJWt4POJSLQCYLDgOq/ow69xM5r+7GlwgqnEPYlb7dhq0z9OZXFC81g6ldIAo3ZU+tWdoqPE
zTMmxhaCqHKk71nGtQAUnB60m/3DERQF6wbY3BmUf5eSwnn7hJDG1mSqf/VPI8MzFX+nNCUbbjUZ
3AkA/zOQxN1pXJJzftlS9MuZtubKgkixjwd5wkmL+T1qOwwjE8ILAbWt2nI88cfBVPiUUgKcMrWx
IZpuQLFPeEPW9r7I/4rRvFZWCXhlxHoUZX0PGlw2kQB2fu2KGmhA28XcqQmppmomSw3xeXeqXYe9
hNLa2aY+SN3WMTa+Zrk01m82vCBPBqgfhBlOtRgSC0bMvRGUqxRaa56UPLnqA0vGsBZeEFB/Q//N
3E8Bmgy4Eq8aKIPJW9XWHG1rk5c/R/rLac9SoteGtzwtgg9TAJkpVRzIdVVLGt8q0zgluXza/LKL
NKuM9b4T4Oh8rOGX6EP35CcEvNagNjb9k1Dceo0UYJ9bF4Hmo7FJ3DFP6/hwQ2L0qf8147MEpyev
xGZ97YCJqNNj85cZ8w/lvr3z5bJKrkB9RJ3Yt25WpqyFpxYo9O9CS8wLzYJvwryRmkjbDiv4x0RX
peKThzubwVh9wxpko3uR3wBkxkuc0RPMys+cwhN0PXiMMgSre4J6GZmF6V1AGIMRZOkwfYrNe16J
PmFXJq+qjXPXBdatGeK7ThDG60nacefi2jQMk91m0ZeCdAVpjKcccohQZvBiVe/egneuGyHHlIq3
GHL/fkQuvjAkrIu5mJakBgtdmzZPhU3P/1aJ5aIqlQlulVxraq6q/3+kRqLBF3MdpHEwAT96L7DQ
wccoQ7jkVX3T6lsRWeG+rkGunT/CvBYi/Nc5UtuttQMdXa3UU7Iq/RolJQCOOZTltyJA4Re5d1Cz
ye8RgfuJ8rfK0s8pHg/FlUBQM0UdV70wKhb1yPQ78DNl7mswKInjYhAACF0tePXz8jDFATyu5Ipb
zdLyCg6AQIZ/nj5PRxA96BmRZbTIMmZYly/+FRfiJSz/B+xiA6jD96Q2Uo1pDpPkIZPbLN1dPHhs
ce98CScZd+KMPlpK8BdyZnkITVWGyMwFLrU27LB/oLvYHobJWbgiJn6Os18dUYWO6mARRgSM3egk
T/BRl0x4K+w2gPbj8802YzA87JboQ0vg8XHcEm0JHCu+4fwdA9F/xvHLP0qUc7HZpW+XnXwcBJcg
ep1eCTmBmUEiQ16vGMjVbcxQQ22zXlsfW4EHd5Lz2NThTW/2L0gZU5o5qLK8A7EiCWjMic2/88cx
ooML8jjOOg2k11U+qOIIknfEFTjVsGNglJRn2vQK25Wa2U6peJOw++WiA5On3lt33GxyuwzydmB1
sGAGpqJOHnOaTAZpZCJsS+1vtnKc+kmDU9UEiAs0+CDDoScaFeX866t72KXdO0ZbACN4LSOfY8b9
/Spnet2CQ7MeqFhMkFjSB/BIxFp4Ncz6Pg8lzrFV9QBqJvQDQnLSNYC+GCMN2bRO9US963pxfSRj
zf4cCC+oQcD/dSS4yZ7pzTyW8ijNCzCND3VdNb04pfC0Dv/JTkiyaQrnwuTcQnV/wZUZn1NZvxuA
zY8bUUNCCx5gQwp5/qQLg7Pl5u8KUn/KGxsCMpeFnlHP7Ao8yIjzIJz19vsKG+lS5e8aCyFFdsWy
gAP6rF4RHuPjX0eQ58mrj9w0mouJ2s5rkJRmYyHY7DCg5c55JKVklYo8laeo02xylfyq14PZK9st
qhAVnZ4CTI2Q5tIfKgriJBTW4VxnN9Tm2npAoA1tbiateEYM/X+H26EB3JmTwPnWevJEVQcy7+Sb
gSCstGAxFfWBhVdrbWOBI6ceBOo4ZJbcBeqWC5pitWcT+5FNZgLB+mElqRQ2zB+oJhq7GaP+wwd2
hRIn7P1hkr0vmgATfKHgPqC1vLL2VJp656f7/rCRDzThuy3uKAf8MbC6d5XXfTk4J8JmVa4ZHZw9
AASb95AzgQkes2QQfdjQc2xgXqFHkaGmXOTw/h15yDhf4QS+5WDBTYzD5XhKfuLmnuGqNTnpEvN1
piDx1EhwwtHxCd7DGUybQEC+tGoKFB17gcJ3XwjP0qBEkFqwff9KiuY2seXEfcPPrGpWv3EsQWc2
n2nI/5wW9h8jsXAlB4nhtRUPCicKs7TRznepV7NLwG0gb27Hc7tI1saKwetxcwgarlyOObNB/s6q
9u2rtNcbVTF0NoHL0Br4E/Jmosrghds+WfCQRvlNDkdIRCEDMgIQzqZz63zKylGatzcsNwU7llA5
uxM8crs4vvjb8HNv6oX7rNbjMUAAMnF35MHym2HGbvtE+8nw4a4VhBl27ZZqnp6+ITMeqKNwxjIO
K4+lgoNpML04wsNgCOGmsZRxFrnSm/LVXAJNQ0Tbka5ij/9V5FR/KthFe91no40ssTLA8eyuVizK
f8YojF/BzLrqPHQJoo8PCITTEamWXFqnLrK43/Ck7oXYsNVmLGnwERNE3TqQa96pyuVfqsmZghV5
xe7KlSaJciBEA+kO7tjojqeHyAGSS3bTHeLkssi0DUgOwHA4+9OcdpFtYOTcSUr+OiE3ZPe8FZrw
Wb4EZBbgvcSS+FzjODmW2+d/3Y5VtCB26I6Q6H47T3RJlAy69SLmN3OBZlvGujSAW5HNhZYjin4h
CIsfdzPkHCd5+MEbuivwA6sGKVi0WcFQFW/SZDd0bBeq1d9XvQAIxLGf9V0bJziMqlaXNg7vzSaf
q8jOKbVg8epjr4d1Dp7r1bCtpud1mlscwels9rDtbkfiag+OxMOxfACru5nZCQAmt5E0e4i+nrCH
hrLSkoIxfqX7+Fc7V8S4LJBEENRgCe0dZIbch8tYfyBAGTLabh2iHvtSRmdHKwxpvX7ZniGW0LWl
NUBLoow0Z7Y4UG/eR3aQjUZiV8j9GGbRZg9aWT0bliWvGfsLRCLBI27JDGIwY8UCzWC1LqT+P6p9
r9CX3pgC4KW6kR8Ys6Ca+M1WoSOHnwErosFPd8Ur0bhNFbzQDU7VsnRBkayFJzS01b8iQOLnsjf2
yyXhyo1/xAGiVzscs+WJIOWltrT3Rc8dOE85xvH9r6VVeKTIgqbX+jWrX4cteCZoGf8oriZhuls7
ts1hOTuVluEx32atCxm1MwjEiQ5wMS47gx+1H5qA51jqWzszFL6xvuEvVTyxqxNaVIK7FnCqCbph
TO/9KnkSIK2H4wZA5miLei2OQ4NPWmtRh+OXbepo8I+2jBlT1v2lHc0pvV4MdCPY3oktQMHzjtnD
iRm0LtbIuKEAfnPruYbj9mhBHVMHYTx9bh81xAGjfpyL6WzMJsRUcyBayfol3eHsVdoiinDkK/kd
n9+/wt4ed2rb3sakE5AzKH6TCTERddY50X1YVR7/a7l6OHyXYaqULK5X2/PKdHnfSOK++I/VQdBE
S22IuL4URDNRpBKesEEwgt0MGjRNl8lVyylWqpH/P/Y2r+Nm+Z4rBlvgN9EL5261EzYP4i7Yb+Jb
lsxEdbUcp6pmZw85FzvJsqT4TnMVA88ghjTci4UPe4An1zE0At9N1tawD6ZaStQY3/KUwXwpOPil
719rX8H34nv6ip4bcJ6Gdzg2WG+z36eEWT5rSjhigvl8FVnrtkWnkLCKW7DN5Pzhpj5Vy0XovHag
FH9g9qPwd0l4IofGxXuhfoj/Ux1YYqHgk1ZyytOWqtR0qsIsKvvmaXh5Xbzci+QTMO9qvxY2eYcy
O7cZZJrW6T+qenGV9jhRQDdPywAoEd3DBxluYqqH6YSJgF+jwI1y2mYZRYydvHTxuV3rAs5QxpKc
xsAds1JhQ0Gva6VlngJWolW7irO/58hJpO4eDE2uOBUX8s3pzI1g+aWZd+4pgYLg+IIgCQs+p+3u
oDWsi/HN7xg00S8Q652ZEddcxyMAIcXSfnrWy7wK7UXRNmTPJlohNh7dxhLZ25F4WLb57VVrlosc
Hz4rZ80cXZNPGTHoTHYaA0jdgcJ3BHLgMHOAClqvHzGwvMd7fF+MMBo2/9H+sx19/zVKksnSoaj7
oKRjjtZpS5yqy+NHoAMiFYPbH3Pud8gwnNCxv6L+9Ae/deu/HUPcy+8otz8sUAN8G4QJ1PRFxTGw
TlKWaUVZWIvfiIwE3KOexiZ/pdXTYAJuG+aAzO7EmR7fJUb8BoCMvJjOpkz3ISVV+XeUFSNJhO6A
IySVkx5rUxYwJSlIA5iIyum8qv7hRaJbETG+Xdk3Otgbf98Vd66ZgYP0f8fxyFcsiX1UZs27kXo6
RGtPk/Kz2Wax/foco2ozoGoz7RO4kfB/fysY80Y6faF57mhaaD+4h1DwFTUh8z4DiMfetNAJlmWz
0Crtqo87AcptBVCk4JMLMvHwSSKdFrNwV18TpuHDkEbAyAlL8L1qNUCpMlmKsCyZh023vxm0Z1Cm
FjHBF3zXpr/w471GtghdGm6yqZCw7/0CGpg10Ddh4W0M3wDJDANyE6iudOWbOYGH+yhl5V73trpm
J5xmD8pE6KYp1PzL9D92Xgg+sNenhy13hS0mQuox6aTvtziRiTf6Wno0vPcqAiXwov8nVT3gA2EQ
9c59WqHuXdBuwNMOgztwx7bCpMxNfvFXeQn6C5KbGM3Fi+Ys71D6yYAf/uK2H+GiueZmflDk+jgd
/BAtpcGK3gKWgk8srC7WKy89+JbaA5TJS1XJtZajO+wFOkpQiZXAI3v6Cb8bUlF84WjuYhSpT2SS
uQpvtqI/HtMrM5RSq/XOdpuitJtQBUabhV6IjsUMJnzWqWcxb09pC+PxA/jHSRRRaL7xv5d+KCt+
g+YKRYMOSxOYrSZfQrC2klKJ7GzqkuB8K0U3edTjlOxoazj3cYCOuIXuqgMTTYb8qotv/bSXEL3a
2CeJTIm8Bl04VhbWn74quar4mlBxz7/HPdkm2H4OThtPvPYU4YpDNMSHzdjJWwLm3PEIMZHfPESv
MhHgoarSfbWHqQCX75GREDW6HYkBN3Bx4C9G3jmKzMF37V+SEAYbzNT5t5WUATvWmNLwgWRBxZC3
hlX7LRGpLgmZ0AWmGunyeMOasw4EsO4obFCWflez5ju26YNCkNfSw9SYBO1Mr+7YaSWKPfiFIjWa
jSbvhQoGCjAA3cJ0BUYsKgAT8NEYmw1UaJKp9HQjhHdCukqMDfIg+qkqXZ8U53XqUQUgaxkTXv6E
TPcOnUjMcbB7X0DGGtIiq81xfOd8f+YvbEMxG3YpitrqzabS8Q9m0ZJiigS+1kYSSeI0hBp50uzV
8ryhHeefTyNUXTn5Bw92Kh0aGp4o/XutL75brS9+1fjEV7SlX0lMmcjXo425XzV/aO6Zhk3yeXWr
PQO3z+5kebW12l2CNe9K2Zm9tFzP9laQ0qsGFnl+x6ZdL3BDERMC6brakuQNFNO1qoMkC+TTAja5
j9d3Fi1Ig9WtZrhgFITbvZcCjsX65zhb45bbFW1OurM7VgU9wKn9MQeSj5OzPhpQEZwMvsZOHSiT
mrQ2w9HMP6WcxlfTs5E8vnLLKK4fcKGCMrFjhZk+ljInDlhvYNa0Z5fOSDjb+Fa5Ia1ghd7JkPXv
UxavaZbl5sk6ZUme7yO833zZF1ObiqS9acFQTEl3oLkVgamBP+IfS5lrbqRLSYtkH/7RoL6HNvhY
hWnWUxozBIrBN8gmEdVLpgMDsVUh/m9PMwuCnLKaEiEeFsfVvs3Ta0G8UOQKCC8M/E9HmZA1/zSH
fOOjFkegxL3W5baaTWqyVvjla39UV0LafLzIrb2J+7H09/gUCS937krwmyJB23yocgZESMUJXYtQ
hT1oZLvTegzMxfNzUYx16TPqe8lYc1arVs+zY0dQ7l2I7RWCLIa7P+RY6gdKU5Pid7XqqQ2JIZmI
UWbnlbULphcM9ZGqiz1R+IPqoDrSwxYBvQT+MbsbCYhFtPAG+iaie2mU3a2Gry+qkXujoLye+JsD
wFJ4Fff9YAUCM0THCAY0JAaNY2jpVwurEsZLQF7ifllRjeIzbnFVTJ+sygFa45VwbD+oDDllKR8u
CPazVh+y87crVQpBmQGLoDW0hGko+s0c8JzOR5iC/to98nc0AjdcaBOLUqVUlj5N2JcdmHNU4p9T
L40smcAFLIF2+cLBuYbAsCTSG7b3OauONXdTovZQogeDZ0ZrdtKsbOnIFRxmjzaHaOePjiWIdz3B
YuvCEluHDxlPbzcPu/g4lgoDT/lds0lm+KKfwL8FzsD9/md8XnYx0XKJbIE2+y16Nzjc3iXlj+UW
ei3N9pff6nvSWecjdr8SaqzdHFoB2J1NwxuPmrxzmY/DT4Q+U9I7jviXaozuWLBOp/dlSY7lDiDy
TeUczvIY26jaUmrgZd4LfpOHGLOw+XzabxwXkG9tMlUCzU75TUgfO/LPThNd34cqdENHXUqY7FMv
z0ms6Gj5wPjRK036WzyTVsFe3tg3pejqNeRHjQbMLKcmP43ce+zHTuuvBzeo/AjvqtnmVgHd+gnO
p3HOIqCR0GBLhy3gMWbHzPyd+yt37zE2w9U3nJv6pDeN6ftAOqkqIlqdwk6zzoNtp0SH74pkXTHd
zsKZfnjNjsZlI65y7xrMRUJ7muP3AVW+IIbP+dNi3fMXXAU+NN/Iezd3fvXo6XFilIavj/OKYuhn
+zc1yjUT4cMwlUM7X3XAw5KxL01jm5X2Cpq3jejlwcFBQTKMCVR28zoxVavkNnjnubcn2kV7kZbV
ZEF3AFuhnVc1GTMLQNfFes0ChjQk9ccmnm2DbbjA87T11NnFazcKbHynrvNCrAklBSEb7P85eU+r
oIOhmn2JXEwscFbDBQbjo9x6sefzmV6RsON9BCDUyOced63OyAxTvglZNiWVRCOs9/kb6CG95elf
wX77aCH/7P8U0xfmUICDqnrnqs/M4ymFmM8sdJjG7vTu4mp/lD8p9nRKV838SI601H9IH/G5sJ8r
Wluq4JXcB0/Ha1MD/4rfdeWDNzwkkuZwtWNot1vLiOnWMb85QOkSNgNxvz0tUu6FhLP2IZwxpGYT
xk/A51VVjszmFLO0UAJCVcvXDTdNt6U3EESaKsxEFHChQJmpuvh1LfTx9MjHkRGrUJpfUiuJsmmD
xXHem1+Q1vZiDLLHMvgkBqC2rgvyP+UHUykVzcA9l9B9Z1hH7/fE3p19+Xa7djpvNGx+0r2ipjqw
+HPnz/e61ZDPSlyGol0JFQKlGCXyB6VeuFC1Q6QwjKaqy3opbajf+61bGujP8GlsMHmp4gUJ8XWa
Q9wORc1pIHszo3qWVALUBRkG7mBD6bsHaGwOrgGprlIczqLY+0Mk99DtMS58A64pH1eoPGaz5l2q
kbXGcySsK/PKn0WOyadkAwc0tPzDYsdxcR/LaXZj4EvuLzthbJpmakG1Bp8SUbMTelfq6aGRQ4y7
wQWhWK6cWLCB6pl1HZng+JcxY+RI+n1KN9qcL3jZCSMeTjywU0MGGtEw0rAMau0Flzth6pGlDOLk
siYjEuL1qlYsFJtPcUMmkMNo7cjUbY6DLPmQ4ehm+MHDZTvo0Z5/IlzTzVRqA5TmTgT0UMtRTwLg
ipMQ6GiSpiMYTugl5nzCTwqTYg4MDVOadEZ1wgnlVw6IgWPo4QQswAU9RL/gkTWdS1zkVQup1OCv
2ZEe3yH+QbRqpxEdlqwNfWzYYN3GQwR0v/Vrb14UhZsnkIErOagPKqRa3roJuud48Yu/1ium0+IR
fAdy6wyYhOS0YJdMUd8FAp1UUnpCPfDouVUcpIyVYQUUZcjlzl/onoLYWS3q5enfUSP++IlnNh+x
nZqbmryZpDLSXV+YqOqLa3C5U9aMprpnXoqZdH4y9EVA4GetiWTosJpndm5KQ2HRzBjE2emIQqiq
ZhdoxlzyuNMCEb1ZTT5oHPfzaFh8b9CBjgP45SL4Blg40rWMVV06tRYDYI586F3PANTl+HcB2zLk
KmdZasftM/qhm7QaECs5pfU/fBfQZDjHESltgHk/BI7B9ZpQ3cfPaVggsT4f0j7iPy/fCWsOPf2R
doVnTiwvWj0hfisdC10vnXDqm+PtO8Za7i6uWdRQRb05Y61PciLFWtzpNCHsUSNuAUhMypzA1Sh4
F7ECBHuuRmjXSB/tB95MQJngCCesCmlrn4gKnMO+BIR1YRK70oeq08xZOo7Tsfh8r+XSAh5YHVjG
Bmyj0dZybGeL6AurzhxAWxqjwt804Zr34hHXYeHy4uu7AJTLflcYlrOVoPtc9qGyRelkvA5+aYnS
tMqSGS+UcmkFUgpgZKnWx7SFNqpbhDp+Y22ZZBPM+ldBlXSIhT0fDS+s70YfzMwzxWvlaP1+/8Gf
v4ySxp8vIBq7WXQvpWcPfBomQHnfe2yOnDozK0htvvBRm9l7Wjip2P2yaeSDW0F2Sf0UANEC2oPx
R9d5O+56I3/QlYkQpNzarIAkX/dHMSRCqpNRffr2JM7fd3Xy8oYhErw8DZ1glVWg/MeWe12BZpmt
1LAx+Zpr5bPDilZXHiBI+5/VcMdciOSd5jms005256dszBb1L7L0Mtwfj1BeRl5NV6tCQBW/NQJO
apbtA6rIMncAqrqEv2NMTTXCi1IIo6otb7u5m9tH0MVPfe/O/cisDv1uorclmJ2c9u7VEt8vVvzK
J/wSm7vVfWj6KQlshYKmIzSopJ6+VrA2eGbwpNX0pIlIRkAh9YmNOxtXPpnWmP22CLUY1kdZ5O2j
0puuWEhoLCC6egNX3VWmbPP6OaQtEvBl2jdpUtlIvtc0hmFnerIIr9uQ/C8z15V1hdySaJ5n30Ht
CQi1kiBNRGwJoDUiyFmLpuY641RtoEvUlsAyPi/6iFxVwIYfYg6oN1jveODeB16uE5FvY/3zRwss
QbsP5uQYGfM1/7ZnP6riDNXUUjdlDVh3EOCVUBUSU+26cb5++Hj6dpHaHJ9QY6bCoY3yBM6ONyLb
DR4VUft/byR3F9QXO5awE8AW6AR1FTgZYXjoq0icSfjukZ6w0ml/wi0OXhL0Ca4rwcYVDGW13Ply
obx9dcWQVqBZPrIV9V+Mo/CWaR3Pk4MI2CN0SRDR9VUGB2x8fANo7RnAWI/b02XfcnThhDzn6Ng1
9VjFelh0QcGmM9JOeAZJGm5fHk3IfWUZkuZU2PDdTAnVpfezJUdnSilCfBjWK/1XI7TjoTXbDNY/
S+/a9w1SgTKB7rxOrUogzQwBJx0jnM3KIXirzhfk76HHKdxCgVJ3jaCDRvK6v65/iHw3LxAO5r6e
hameMc83J498G7SIx+nZK8XbW6h07fCo+MZ86oC1gkPgqUP6rC06apjzuKqpMCo1nuk1yi9xm9e0
aP9Yck430fuKIGiveEwVylR84Yw8Wf4/v7diFxFEf7aBdwvqQoDS3ByV7wLuP+Ni9OvSX3m1Xe1p
5wWQg0pcnsgXPsfehoK1Cbcqs+zrLUXGKP1CqS7TfsuIBLQEAF8NJqegV18lxAQS1KNiOxAFNK30
SiVAOVgLP9KsQvGN5O5/IiuDWRP/LH9Mksd5R2O8GyP2IuD9JXEXPgv0wEDgZzDyxBh3TQ+TcemC
rqYTh9b6QSOcGYqub2rNXKrqgB3djTXdrEvuI5Z2klTRzfjVXSIRe7pqWqYXL0VUy4h4dsUMUI+f
cwAT9ttKKFIeVZy5CnzCXW+jWVp6ObAI1+lhP/oHQ/EV5tfINb0JWNyxfQX4SLjLpY2iYjRTlrA/
THHG7cX+xcxXmeGLWGdPtyEeuJhq2NeJg3TgCPanAfoaau63S8YUQolIMns1cRWM90jnMbgI5t/E
1KkBdCDmn0JmXnEUFoWJ3a4fdm4AIINr0QrjZ4S24SZgzD7PKY0c7P5AYqEk9WuvZyO4FsF2svby
UoRo1MeXYUgnKCz7GFUwTZ/4uEVcQNOVp6Bfd1/yn/xj3amGjHg3dfEgtqqtS1yV3SOJxT8X3Kan
Q/AIG/YY/fdU6UT1A7SudRUo4hOFcEwigYW40tXKEUxtalC+c6zLaF/sdRbIiekAgeuYSUaKqBQF
n57Q1fGq3815btlRvlYqMOiW7iVVk6VmInF9XbQP72F/4Hc9Kf6ismgRh/Vub6V9pc22fB/hdozI
/e1hELY6stjfmnhIBasKbzrdNY5rM9vuPQ7vMPoHk8T0Qc80SZDbnhJsBBh1+cS0x9tmpnSF7xEB
WkJQDpCFFlWykuAdzBSeKw2N5bM6IDCKDDqm10ioQ7N01WUWAGgGcYJTy51CMi8Dub6FLtqC8p3m
m1U68NlR+BylBsccJyo0Lxjxj/cb5iHBz/tv+zn3Fau6PHjW4LyKfOAIjKoWPysUE2jyXqRFVY8j
loiKR8hWNgRckdTPxCp7xsw5nto23U1x+a111vSPIAwhkFJl4Omb5Wg+lAtYwMw1Efpsoue8MtFE
ap5hfWg6PcVk2qkOT4Y0gAxMULXQBca4PJIQfKjb/0mTz7Gst+bTk6bCNC2UadHFAaXdp34y84Iu
E7jGkPN0cNS+1+q7AGjrx+NjvbiP0ZGVx1h9Wk9tXqlQurQQR6259JBaVC5eaZOwp/MN9Ps1PvTK
M9fT7Cl8h/vtgHRAESM5+8czStjSt0JPDhF9Ry36xvuCbTm5pdUS5OQgLmm9z1LPcOmmiuI/Wl34
RANf170k8IPy1uSqkFYT2OIJqhvD7QNwoXNbyKB3yFtlm3RfPESeDLEUHrEwOy3CAsnm+9RMRpjb
3x7SmMyof7WWAbFanfHI3DteJCwGVCny8W/k+WI7kZzRf3S1T0n+jIRbW6o7frpdgZFMk8yC7LM6
E8GfsPwfWfVywIj+tHYau8eQpD1GNDBPYptKQ1dI1XknjR/ZU9n36f4CHbpC6O0e1FYWMGleaH5W
6eXfpHV80Sk90KY2+ood8/DT89Mzjf+PsrgmgjaszQysXSym+7Tls0jXIo4F+b4kKmUowgZlWV1p
FpkcTKy4c902k5vqocuH+DQe0H3bFvhTMWAZx4HHCRUlHBuJGEI/B4U8b9WHpYK7b9Z9HXvgArpN
lM+7HDsNvq3Ywa4St1MXnlDs7oARxkULwmPTDDMMZTP4wjnxa/RbcivCr2Fd0ENexbRXZQ+7Cf4L
w4vcCwqtSa3+x62zI4qtzDhcErwaviCuDLthOvOKQo9kAAZeSyegl/boB6u81LoCW6/KIandOA8I
k67F42eCs4nzzxb8SSuPwan0TZt6xD/QfZirvDqG+Wz2MK0Oo8qWsjvl0W7m34CAsEHPF9DAO6M8
s8cKn+3KVY1fKzxvpGXkm1C6pwN2CnuLhnf2mAGbTbZ8SBHEJ2ZgEgpZ7Fn7rk6DC+qPYNqbLZTE
93szDDJAvhwqd1kZh4TwXLYYj3NGm0sqa8JahK9UuTYRPUil5tnDriFPQGje3SJ403nrfJQZaZh2
ZYTAWaWqiNkC8Z45GiZtAwyT0vSjlYtkMycW2EDcvDW6OWwdkGBUAvySC3g4h5hAVd9e0P7eNSQ9
zWdcvvCMx+Q+kes+3NKLH8Q/DV0yKTTxCLsEKNw82l2av63kDlnzu+8tCbxMinPzQYMHHRkWVhTV
19BLt/abLYNeuiJCtLn5HJfr6LooKsaAmBvtAj5qbXWp/iRoFCu6eyA7+uy0vrksjM88f14fnSZ5
DeZ6UoghoQcR+1RCb7zhOyd8uKC78vzeXUYR7AU8Eli1Sxdt7KTsYyuFDx/DUcNz9Q2meWjJIVwP
AJ5tysgPVY8anoltBZevZ0IsH+Iu3mldY7WXofOOxgOPWCY+8pd3EcTsHfbYkh3MDmCRlKYSK1fQ
uTeOK7kMA6sRaWb6QFe9BX9/jlap69bdzr6WtvK8kjz9aUcZtItix82xhQLruCEn+WNBzz8Qc9UF
vZ8ATjlg79BaRqxg3VyYpeu19YptQUzgCd9oYJJGbXWVuCpsLXmGTvFNkpTixJCDiwBO2Xule/sV
L1MuXFi+F91n99DRsXbqtug7D7IbWaxFwn325l2hoDwrRzNqp38RB/EF08VHVuBX0K2KD0rbyFNP
sCp5oRH7yvrC0oQiQXh+uR0AVA13++UB/GzgB+FD7TuN7AK4P20qxshxHgu1BL8ASfNIgbsbrmEn
J1u+slijR61wU0OO8AOKoMKuOWcUQifkgm0ZAbQ/3PVR6mVB6zWxBm0MHENJrLNwrhZPv7j7+c9z
mZSnjsbfzqh+xPxQ32c5oee6dtfiqZf7vttCas1I9ib7EH2wYE6BZX2Fumax2VxxsR3MsF5s7yAG
u5JZrwcDM9+EopIQTyk5FSy3ZNnaqZXh/TYuCHlpk07sA1s/iBiCK2JZk7RmVlsNlgx6pOCwBGcT
x5xkEpOOYpQdl4G5wsbXGHhRyCjxCXJ/3WqQnU5uoQ7AqxvwajSRjlyyXe62yL128x0WiQLX9gwh
SRd1Bq22Nj7O2ICVFPe7z6vz5lYUXQC+IcdHEg1c0171sxsnxWfTZ/ukHskylyobxdYdFbctcVmQ
iYj7wiR9hNmt4CWy9gl9YNizz9oekyjTP3SaWVf8718JQhpV52E65NkwCfrwDVq+/mQB0FCcaLbF
pCV9qfhhFoqn1GzKKUJzALQbyX6LFcHYjyc+/a9YFKklPeYU05Kv1JRkJaW44ogqNysSl0bDrYjR
58pjHwDzFWEtaelkEPQOJ8UKTczqMJ2hdzZTbaVCTqg8yo00wU1h552zbA4JDE+zoDHi54n84Qki
hu1GpH7OvTjbZTCd4keGyqKi6B6KtnZX5kmSfq7sTsRz8fpPQ83bKghQfnnOH2r3REAI7XeF868a
XIUxWMVaeMBG3aY98914uDz9ZNErSqTBXYr/xw3UQK4zLJHFxnq5wwU40PW7GCsPMe09otCPzDkT
wQ3WynnWJPZ2r4cHI0bIKTvpf59S/6vWvOMu0AYcdMkHJkC+M13wwbvMX42QOEM11DgPj5u6Eo/G
khyAGaPd8vkoLtZr1hCjaKcGt9k1xIUT0pf3eOgQjLgULdE6+NLOOyLG63YOpUx6a06ZXuESkJif
Q/QRtAWS8UB0DzlvIdylI/SkJ3LbLOKGeaVUeY3Ye1CXtVyO15GFveB4RwvPG8IQe0ATg/mV81pu
QUV1vsq7/LienuGASl0jDDoovDxxKmzor/LPNGCCw1T3dhHHPd4ziFPiCtNoLnXaRX22uVpFgRYt
h9QhW6YdAtXDjQ+Ke5fVappMU91lRJ4F6XcZokyPJDtBof+EhAgXfCXIrBW2ZrEAmp9BUmtNtr7l
Wd/uLgPXb1Rrvp3jgPiJfKRnumfZakithRvvIJlh4Pabbq5TSXcE+irgDtXphlpBFQosrE3AD9sd
gyH0gyV/IYmktPAEDgY9BCmLwWJrGWv+Q3sHi3JF+mOS5GZOWkCvrEBNaDAcBndefGXEPz+Xxjdg
sDRF0EWkWipmZ0PNty52xVzq0eFZuWNOp3jg960ja3SJ5p9FYTb9P/wnVhC5oLlSjYhBVygCKCVC
91fzVSv/DxL1KmzOcUcKukLPAr51fm5tnjpDq5pkAemkH1g3b9tbHF0K/t5eMlNnFTm4yy2uIzHE
eN0XtO0JvOY1VwVBa2AvtlWh5MnjX3J2dsPWBo0i9VkvZC49W8ldblRGjEptLGXWD+R5MqG0Ogzq
iYLXBqhJCKLzkmW8ABB9AZ6VstO+OEoSf3FA97to8hteN1ss/ka4CNnCjO7SeVAw3HwaHEEBSU7X
WC+M0k+Y/e6Z0eioh/kvHqwGCjat7ACQr7oCLwIWlvJR+6HehQ9aQEQlndvMtifj5BTouip9jvcj
dUctZEPO5gIfRc/wKewPQ0FXeSTiBAn+u/qMVpSOlGkTHmIcxlgbf/iqZw5w6D6gjCLFPvoZPk1J
rMJmP4KQ3qSabgt2LZBBAe+hKC3oNf/IDGfAfd0M6C08hd3/UJkBx8viS+ffjh0jF8GwcYT7XURa
DLeAX58Id84HmSHgrjizjKQ6gPy4f+hBg31x5XI/mvVMlbgBf3Rd2kp1UxE5VYfcRbfipETX97Qz
vgsXCTMQnKyy0LrnGa1lv+BF+FlyZ9exH3mAb2PSfJk2o7vlTolsNDln498z5ByN1SgtQ8WUXiZH
tlZReYF1VoxOrKtKvSmiQ2Fjh+KLodD/Pw6UucnZCK9P9vrTS+0xdS5yaIQNiGhJIis4NXFJEPDn
IFCz6vnCYaI7Mfs7ion46Nww0ixyiy3XkfyapuPj22RzN2XVsE7p+8MBVbhdmwrKEXQx5reCG8TS
1C8NhfeBeB85D1KHssNU38Zitzzd9zcQRtXgg2oAUUn1/CkTiCUQKUR02m1OxQcQM0lslcW+KSiz
BmklZ6+/K6paz/OVDeruZ0veWY7Fc6O+7WQRWSczNkp4BN7fVhgMW8vWFmx2FDPj53Evz7f0INnM
VYcpbcDzAWEfMZ1Y3grQ6NSNLoQd+2OQoF2FzkFYtz1YNXaQ6XL2tlk05kMwnfAKx6/1pO+8HKLP
lEA5EUQDLcE/jBL+/0VBKgmloKutJ1yIy59QRrTAlcBRxBsIcBSmloK0iSYpFJN85X+i4LmBN9xu
k1b9D4sliNTJ18Jwuoaob4qo5+KWkO1RTgCp905n3LGUSCvyetWsXCXQ0AASWp9msWpDpb48uXHu
fKMGemwmmDar11TWt/jSaRLW+MwQtpanb74QoQJJT4IhLHDI2zKqJXdKYEK07p57Q8yXV2pTimX1
PakGe3z0GdliYKVElTJeflpzewWcidyR3ldjDnIvRs8gGHlZImbC5S9z/pYD8oCB4EwRlE9hzGnD
QVSWo/bnU4K1/SIKFQ5EhI2OjSVHzjhYztpXf48cm4ZYnm+msZxM1eUyc+/CPoZwEXl0JgYpzFfl
8UY7yiLtnor1BX7z41o6/MsBak9uKYYUdysO7fNV8tv20Npau9CnDSN4ciqpZkuU4UML0Lmh9X9T
UKSGjD86pkIaMqE2bvOg45Gn8p6eYEiDEUNFRIYqhIRKPHL6Tu2oET1rVc3cYMQ1Ph3WmeW0OG4X
/L5V11FlUQNmYf7DPVuXusZoN1OQlq/R+/MzeCy092H6r0UEDejrODFrJNb55rPN2SUSJcKp64b3
7zmrVrN/AgM5Y39VCIEUYITpJNSNRhkYcp6gLL7RfFZDffKh/n5wck0zJUv9JzmNersP7m5AECyq
p6iujVabOaE98bP/HzJFzl5iLEGBWbXNnYyp1A5zUzHRpwFf78G5ugE6HSFFOUEmArlc0S1aadeK
WlCGb7oRU73/1Y2xWfwlll1WPVNASMS/nU0NBpwJLxGZMZZ0k26Vyupu4k257izFHSfEHsdXmJZp
d7scBjEXbhwHi/7kxw8NFxEW8YpL87pXJ15EMLbyvVieaAzqMkCjBmy7WPLBoBCHuknVR1MwROVR
BXVTANEPWCeOuW/myAMb6LzKCxEMu0V/bMXx74njM8U/ur295SSsck2hocwSS/FgfLBNiYd/JkWy
aSZblVpO+XI8mafu7dAEUZtdp5DeIcXX3RN30JwlGr2ICaL+duwUJYnxYOByDUUFQ0RglTRb8QEc
NaHA9WqwZMbzvQJdNmyj5iaNssqdUMm1JpeoeaFIptu3SU3sC6bQXnxKyvowM/azGjh4Cj/ZKx0Q
xOEIxAwAtpUrMiZ3IMBbgKU79nr+BItsxq/U2EIK4jpJz/jkX1CZwpxVkxbYLS3ZHfVInvC76hVP
geYt1o0E0tNZe/ygrdrKTQjCIflCAguDRmcBdJ0sXc364wCKfsl1rdEsbzsHtzUkhjdNtVyzpxz9
RLQjzIxDNDPSrUVXjJAb1SYSyHe+LA9OXftYxZvlNGIpO7jI01x7eo4XyQVqmVn1WW74pL7pzpW6
FGcCwDsjMZDL4pB3kxcYzt0qKblDF0SPg6oyKWB/wtz3l9HF1SPxZByghCx+oaUZS9unLRIOOjBQ
WXHmDBqVurVKM+g9KvHIFmRwKW2wfHvAaqVhxl752eX+C9fBiwLQt98qdmtPLofBhViRJHOsMjF8
LfxmOFc/A4a2HmWfzggxp0rmoOUV5/w2v4K9Yh/hZjsrjSOW7Ihqf1D9VeKAu+5Rc8ACJRGC2NsB
/evZkJWuNjBr6B7NF1I0vUDsRKwinqAIDb7Bq8+FNVqVQlyzWN8hGs9LJACxBWBXCnUh4fkzth06
7CC9R/XthOiSvtGt0ZlmUDr2MDBp8jp+LTDg+ZTbWzSYrHxfYAq1LBbCZ8Fvh/3P3mBv+qhgKFhI
hSluylpcfEqWUbcWkhuImfpYnbferl43MzFElyef+WFYBb6GTtow7B6U0vfd817hv6t5bw0QPoza
CtGGSPjWw2tGOalG+1jwAlSv3JbMIiDZeQBWGFh6E6A0EUYHz4fvX3dHb9XFqkTscaSSnPbBN5lB
r7W9Pa9WwBs1jI0HNqL/Yfwbq3q3wHvKTy9mZevvwZ13HgyIjLs4yjRgx8QyJi36IhBURyl5N693
4tp6Quv9W6CVGxUOEzeyC8ar3DcXuzWXCpHZLGDKqSQDFNR3T1QY68Gt3yS8vl1L9Cg75T5bQx5W
nF7yt0DDte9eRUmILyA0lX9ZpIAPiV+Mo9mVrlcQ9i1xxFwRdZLyLZmlozMLZD2QEHtmM0IMYDe7
aYOBydDdcf7D45My0a/yr8H2Az7bfT/Re9zAr0fuutRgJy8Vn+pg0UJJkqNvxLF6T3qAJ3d9h91X
jcho95UiErlSeWPdQ52pY2hsKPFBwTmOmV4OGGizVf2qgI4+5Sa/mj+KduJnnUR636D9LG2h4qAO
uOhz3hz5Nb4KXv7ykQC0yc3tpuTATz4/ZCQ9e2F8vMLGdpsdeAO4L3XW6UlLZI0bpVqhYabklRu6
8/pWRGFwUUAApp+gl/JFK/nB44TypshRBM20ySp6sWBWYAXpL5L21IebnGJjJWFSJpGczRxKkLF1
JLLNq/wKxCSYQmhoSsY1XRGFkD4MM14qax2m+B5HTcxvoMEcy0fVychkc1WVBOVvH59hySXfRfE+
/8EC+50kvjq5BGe+65HLF2aEaYVdUT3UwbfsMVQApcgX7P7BJtY0PD0HCFiqjP+52HVv7Qoa+wtN
JQ4v9tUdIR1rvU1Z7xaULzuxMoWoszG4H4WzuzxvlKCbd0Eg9zYJqi86KoZkJ8noR7KgUTeNZl+p
r5aqiPAGeQ1c/HL3eKsF8gwReRvtiYIMuROdWXCrlv2C8XB8ybB8IrbZLwrXxJgr2ToG7ZiOkbYt
w49MpOZn1kXwC0y+P5CAOxwfJHOh4I6GmdZhejrEtbvSR0MmGN7nHi+RL7QSNIseqULZXytz5ANR
iaK32aON65iONxyagWC9p5lnppwa9EEfCL5f9nhtyPx4LaKijs963f+ao0/Zdu/J2qJgOwVBY9tH
EYjUq2zJ4YbO0n+Yng6o6sYUb5IZbf8/SX+oUJ4Gg04XR2pTsrc9dyGZurXyDSJ8wfHMB9BwvNxh
AwoFpHGuQxB0N2uXReslj4pglzJhT0FX3KZd9qGhjnivdwWGRsG6/S64IiylP2SMThV7OPeiK9M9
1b94MuzcJ1dbEVwhYenRpWLUJyKgH48sHJ9Xz6uIRdKElocREA/N9Qs0UTuJp0f33g0eIdLN241P
Rbj/KMGGbv9E00mExlEuTK3H1MYmqNN8jrhJ7yT5tczdQjTQt6QD3yCtkpqix33HxwT8BziZCKXl
9fcDZ9Dba5wV2NMj1qWJle4nP+1P+Wt2R/In0MFou8JDJEkoa7M5jc1ClERztZNW73AacZN9Y/Nj
ddaPHfOcR8Dv6D51b1muOsngaIa3AXJHcaQo/0yWJoQsxwm6Kt6kJdVuX9E1IUTXd+v10dW5AOBA
SlRGPDZ4TgnUTVuWLVbZPS5KXy/zo2892jfxP4dXuNyJr6zMPbsR0Oh9PcyFGcj7xI1OHVDKcHaz
uh2rSS/ukp2gCj8gChxqWRG+kYhqgqRR5Z8V/1nzn4HOBDe2j1LHf9mZ7DMZR4UlFjaMT2Vlk3JI
CuMFeVVnGxAedXAnxh5LVEAJ70s/+jyD/yWpt6hehurRkNtXPJ6SdF72GHP3RjwFB3+gJM2Gu/kp
hG7hjrRZ2ZfU0B5n1ELz+Kfp2GsOY2eYjp+0Dc5GU7om+8GRrpZiUd1dBXbbUGT0ocKmaZTUVZK7
U2Ytq+nP36SRHOoF/ow3dNNTGDeJtZM56iA9eziXJ/3ayobjGigvQB9z41XEppWysw38hm7XEzcL
EPEsAaG5yjhwswxNeiAHoCmsVjg9ENYyV30gOlHQjAQIqrNiTrG1G3jb/XEV3hyXZ2boZ4bNct1w
aDWiZgcAE/BDhoX1pV0cE+0+nO1/XfXifhgpILLFhx3SVpoLymoO9TaUgZMM5mOUWf9PClnx/iue
yDDs6RiLXjdKiNbAtnB4ObVYljXxKzC6oRhh/apQNqGu8TPfkPQ936R6cjfyoKeKboKS87kInqmj
tdRJMd9QPcCgVsFZPtDux1u31z5lyaHhWfeMSnpQ63UNYXn/CzEmg2s+lkXdbf7HsY7M/y/VYWJ1
2vjA0COcvKSmbBCuJczUF2p+l8o2Or/U13nCLiAlLQ03T/H4LQugktARSPIWdwEITQKzd7a+0NVW
ZSnJgWVKV8phi035UHBW3ircOTY/LdAZ95Inrk3GE88d+M87msJYy3gwH5PPLcpfzF/KUFHKkQB3
50ZjdW1nBOx/Bi5b+vQ87xB20y5obTUdQym5N0l4KnRLcOtg1C53eSjnNgGQBZ0mS4tV65i0rTEW
aZqi13Wv2/Dpi/wSCQnh+O97AnR5wWnLWHPe4igbjHWMk7hGj7hJ8iZxfdAw5gavMkYGY8duwvGu
i53hnEqwYWMMVmqCtZWJJTpBNjesSeUDZ7VAJGfhNEQlrVFfNr7Hz8f+6mXb54qwLCCbwafwMzRD
Rm+ENW51TRhKqw8Rc53UcKKGe6nGpjedu01Td9lmCpLDqsXEOjPlGXvU2c6szrvtrKLTSrBO+f6K
/kOzsv5U0gTI83S1G7X/tlDrbKSkFYwP2pYs1mq68HlSjhOrCOal7hPYlD/zypd6Jb+p3V7MEL/h
0ZMLxGOsv+RL51SEwH/RIQLkWJp1RjC42eosYDeTwJivPyNPHbyDjwiKQcqh5i8DtsMnSEFaPym/
7c7ouSbR/npVyhNuV4ZLHjlMghj/pr9lFqKUaiX6kxmKQFQu8LgtGIj5e7VprRrywb4+IAVANfjk
hBPx4PdzPlsBOplRtl1W+3QLg/UIbwoqMVGi66H847tgsq9yK56Kr8ZA9newFyiBiEjwcjw6/Cof
RJ/7ofkBv4yP10cBchr93dLPEwyXh9lrJBPt5U6/7djYrCF12SEphuZ2HzKmxXMzqms8iI7bl36o
aWObgDu1vPgx04FfPDmumN1rE3NYXiydGgl0Q+MrvVWg2/BKpuSsPvuz6lSXzVYBesv2pXnIlESK
OjfRDHpoiuprGeiA1JehTGsuGiFaH8E93N71e1Pfn9g7MEsrNDerR+rHkZTmAWDelgTnToSws5Zl
lGNkhE9PYmOLfpNEqYMfZJfzTTnIOLKRNansDYgBvjRsUlHI+G6zBUjjDJ6w/E0dycybjfhCHUfI
gdDI8yNqlVB3tb0MRJfdAVb/Q2M5YuSjzVOOK7hl+hquK7IIoOuejYi8bKS5OK3PioRxhFskF7tg
phHXeTPIt+qqRTERx6qwVdKL5XVTN41kVe+NZR3c4ijbAW6K4s0VZf+XZSzVrW/i9eNwFc19P5lW
MIF1HJ9lmn7WW0sUyTudLdIGBHHqDWzDfSAeWbri+8P0pqB0Yg9bY6+ZFEQAxYxRXTuF4qWrN65p
kxNVvfAlbxONDG8dDh+PXKsr2JvVQ3Itk3fMmdrAMEQpIhxM+vPCv//j/ab5j47ZXZ1wRMzdpaf8
JoM5qqhH/CAozjzgeWHP1lBNIHho74XSgECSYgJFlmIHNG8+Yn2iLTF2KZwfKwXK1DhXNQL8i+hb
gi66Aoux0XUctXATSQ3H13+yJjIHBb4mHj0zeEoIt0tKV0/roGcMMdur9a0VgpjzrJ3jJ53H9fAf
xECwfvjGHNo09+idWzIQR+RyjymnDTrNm7jPzsT3xZp5aBam2UsfBNqwMvwDNmzhQK6YWB/wkiGY
AoRB2JAEdgPKtFBY5htvNkiHSivtuqpIpRFo1deZSysGkC/ZpnKzuJ0EDP5Jwbbv5hO0Ty29+yd8
CnXmi+9x8dRX4uhko7098fgTHQOUDaA0DjP+okWSrSeq/D3qSqXohZAHcdZF5L3f/SPQ99dFyJb0
0spZUiVb4ZepFZoGRV2nIjVgVFhHqzgwp53W/4YD844XG2FBrgpMv6tCDwkXRWBmrM+DuLp24JIB
GenHCZprXO/Zhce9LbgmhfVhOCngTjvyM0k79xIvAkca99gqimnxsnaoy808eLjf3MH/ILUSsywm
sA8MzCjSqtYxqXYPUy/jL/v0z8CNnEspnpGcspY1IAGw91Sd6FgqHMmG9PeZYFwqKCa4u/m6xzBi
R/wcAFZ9y0XiWEVtYMjPN2dZkLHAM0Jt2ZjlmKnsvAzxRgYKQ65g/sGre87+VUI6F2cAIH0J8Hpl
0yQer4dripx+G1cvjVRZDUG+knhcGZVp2OpGWQ/ohFXRjIiBfkr8Yb6f7NNG1UYPICvHGvjUKXSs
Yn+77v2d8tnfyYOSVK9R9alDaYjYIUVs2GGZKy8NL/NPIKbfY/OKryx7U5uyu5c7uHkk6m5NyPiT
1+pDSX8IH2iVRdr/faOn+GxJo5LNSvhuyI4uR1w7TDBrLvlm1MSWTLn6Ao/NboqCcmlR+3q1VHKz
lr6mTd9NhlkWgo/oy8JN8vuNGvF5eahB5buKjkUeOulUBq0OYhsnRcGYlsjYmI0vXxR7s8wYdvbs
2VG4qlSXfAW/HKzltMtM28YbGvjnk4AkZl64lc+DMPER9UZxwQ5N+uDTVzDybY26sF5ejrIfF9va
w65PDT2GIej5xlZUT/hfhD/LnqbtPiRGHqtdlPiJ5undJoeT8TbiS1TK+2O6HDbJQhC67uEUVeAr
eTXPafeHM9so6hHGSKoB56Y4NLM8ZYJmPXeK5tHyrW9ytnY84omch3ZKJUU0Y+gPFzEwHx94dTCi
FIqMSFz3yVsxhvheVEhYi5W4/FLGCqmknvhhn9/TcXNWOTslVTDEZOcWsExTbsrTb168EnwjIL3D
A7dM2YXfnb7Qui8u7jPUjKyEhKRdkowEH0RLVMsI5lVGrUXENBh44yuGKhczNUP9ldTRAEQUSjwe
4cvp5uv9N/m/e/yf5uQmsnh9tpahq2S04I0um06Q54rEvaczXx30/KGuJH+JRa1J25X9u/mYpQoq
hQw66gaUkcVnTDxoKkGKnSkueFIgmiqdLomwrr388MQb71iJ1UBGjzbCHC/zaHCJje4bMMdX7JyR
bH0RRp/hzSfRZYxx0xWNiVPLtIbIEqE678v+hmGOaIBN9YPSW+Yyjm9O5lJbTG4tOvQF8OJgfdVf
YMkqG7R9Q4HIoXp+2nkzJZ9EnaQbEiYQj5J4JesQiQzb1uGqzlz18wl0MINvPXADbD36gyQWdUGv
WfP8QaJyihIhsv+6zt8iI/I2CQlERN+LXgHZePp0uShab67bjdUHYpqGzXooU6p1SEqzMgtQYk+X
7v9HhViyhsC3G1rrqldXcv0jAI6aKNgSQaI4oeQjoBO/4IuoicBVnas01u7f6UvjFHG9qu469/RT
xjWjuUbpKfTJdKhE+jaM7seNlW9QaJ0dFk1ZRCfk2AQ/0fUgDON6h+NgAoc1SjVnBvIk2UsYlsGV
sQV/vSZvWZEscTsnMoxqNSxa6FLsSy8bFpyJVsZ9aUqr6hsTyKBxdqE60yZNPD+d56B0XFvV19cy
lxLV/GMpC+194awrzkESBH6X31+ORYij2yC2WmyJezrB7HXBCAczeDS96OoOlAVh66xRv3QpdlHZ
/6GQIazu3hjAeGKY03No7ZpLs4vvM9Be76kX1N+neqPVH3DmhlxFDtrdpPjL5JVlJRkbdQ5eIpgv
+iXN9J3FsDZV9gFX5+tbMFJXJEsdGWoyOfb6Vze9iPazk6OkAu/yEqFXVn6hLoK32W5tH5XyPDgo
50+btMDN3PQZgx5KXbbF2GPx3JJMVlpUa9ccNjlpyckjoyx/nG8E4fv1MTEuBK1chy8XHgN5RG+u
iFmB3PuyBXylxuCi3lMK/sDCLaUTkjkGz/z8oZJWnjvsLUWpkUzvpFWZ77Jke3CbiZoReRfXUP2x
Q5D5UozYRgduDydmyr5k+0b0BYgfZHcGty8cbG/Ef7YxWII6fHi0LcTxu4xDC6Hj9zS7jNczNvRM
0uRDU2r7wVIHAPcOahXB73WH0bRjznsxcJqq6iuRDghxPyHNuHHKZJ6+k6sCoRuFAhXZ/PrlBlqu
lnQwg5zlZ6/x+9qGF61VX8UA0QMTf8xsPPJtmn8mbXY823uNZcroDCLt5bd5iAEOXd7xCESRTsoq
/nnX0hbnzp9H+dUQhL0A5wjyP3Hj4v8SiX8XezBs5KpmmPU5PaQfVasJ2CXyVq7MzBUXQdPfzaoV
xKgTccthJTuT8wO00NGGl5Cz1/Nc4RY1kqnCHuRiRwOyoQH6v68P0UDl0f2jGaXJ+UXSalrCSOeu
qTJSm55xTfAb3vNzUggR1LBr1ukdT2UavKt8r1NqMe5Ph83F5vU1iQYnpF5ZGNXP18KWUp+15iIl
xg28WjgVMi4CrH5d4Iw+m66USLy5J1eOSmrYTPxwhd6cpEvMBuppAN0TK1ZthE03PTncjBt8H2xh
Rg7e+oMnL2DH7uIbZAIW8ECal5oanhsgpi9rb13n2wM0WLfYmEx5kAlxszMlRWqnWll6x201vXj4
E9c3HSeMjjTcVFWgrnAbfT8dq/5Osh4MLV7UgIXgTLeYJ9Pin732o5x7vULrV9kDUo2lfWLVvr+s
R/uA7AhQDx53RT8zUj6FA0NJDRDduy2dWYUE5l44sWs729BOoBQI9a43rTNUfJGyQyiS2t8Bgpma
8hFIzoqDlK3q8YEZL2hvjeVvOlAcr1wJwD+ZtU4wahNrVbsM8q9kzCuy4P6nAd7hQIA4O3UYE2BU
zr4vTGaFh49miUF8XJIbWUR89o2nKB2PmAVIL+xQh8JbBmnm/Av2gWMfOhuFjisn9ZACaUDZBcle
bbRuV9gUcmASEhfN37B/yxMUTYaDFKVcNmLDv5N5fXOvyWe+wGsVahQV/wxdej7LprNFLQQKBnWQ
9dCcYWXLWX2wMg8nWfYtGcqlrx/8i2e/iyBdoWIVx8GB75ri5WhnBGMWLcgt3Z8Um0NX5IQ6kgQC
JyVyWbTnmjTdx+GQLf6F3zHvEASLauIn0yyAJ6goeTrzFO4FTgZ/xAkfujU5M/CnZysHSRzGJNv3
VanQikKS2GSsG6DNNMOW0p7H3he+b1gsjm0rAVvRK6T5byXUncNcT2E1jlMD+XZC7Wn/9prhGXxZ
xZzPlhbb7kdsw3ZUCwBj1/9HBcwaPtwSoAzmkUP8lXuNnt2wzg3tSU5jgoFdccZee1k6tuof2Nid
idD4v0bY6fre7mjMRp+aHh+7t9WtxjBs0tmR19ho7xTjVbpD/TxKAMgEKIJnu+Uy2l5hGU4UjwBQ
QVjHV7Mmm0FKPK4m0TLKUo3SA6IA3uxOu9XZ7Gf/6yLWDGxPzJab0BirVmq0L4DpkhYjpWhZQu1A
CxboKwEeK5BGlPJe3bE0oob9TKl1aFbGokUfMe6HH5LJ5jvY7TTrOjm1u/MGXBuO5tOoYFfr7wXb
gD5swYypfVqaXMaifFTnOrOJhsAyU3+xN/T4yjPrxtbmn/szlsJaLvuQa3aQGHlWamLol6vlMUCX
os0/BquM1XK7RVXPcfIqHRa3iRae2lZvkKa1Z8IYg5euS0Y/uN9zC2zhjrGZU605OPM731WAB792
bJBL2KbvGrvUsfKhw74UVpmu/5oLSzINqdTNnQLQZGxrCdkhgE87rK9aCorahk7f7uTaYBBc+r23
YkUe+vV0Rimuf5NLEyPKyU0SCTBetQPsqH0WWoGdwAwgwsn6NV4rdz29WCAbyWbI2YgbPkXv+J4i
5XameTZ75MdK3olSM3wadGnPjz1xvpZo378OsugXxOD+2EDIG1ot/zXOnqu3Hy3wBJ/4ajjJ1r3J
A8QrJ3lk/NLfkXjNG5XZRov5GmXlBJRv9fdzX+LUQymVH4d/h5fWUyDnI7Y+3xIyHyZqkCbVNEoq
MN3poKSdY486uZUKLz2b3uwBj5aZdLnG+KtFibSRyEEdcetSd3rOIUUYdRafq1WkV2YlQpNRV11z
NUQk7VHv5SweQm4QJgyjGVczo5L5dX0fcernNzNVUnjuzBkD2hFO5ZGy0VkVAfPWnmdUu3PO1hd3
L8zpyjPI03ubrVYeMP2fZLAWFH77bSED0JMAasnKHlsXhAXxEhOeaJ7TcdsQ3BUalAiwxF1jMQp9
2byyzIH7rsoDgqyGhz3US53FF5KddSh5/pFBVI96BJ+/kT+i9XWdi240bsRqqNw+82PI0dZvdusk
JabOU6kTSOx7PIZZG4fQvRMSuIP5CaqfArFJ4x7rkJOv/tVKgz6+BwAgvfn2ct8v6er7zFSGGqBa
7akQ1yLuwWln4M1kewT+McX6f2f69uq9qimaaXaoNpo0GLZDElj8yLp+I+nBh3aE4IjLrNTSWf7G
PfLKrOZM4tsi3Qj3uDX2z75ePBFNE3xSI9Z6iaQorIdfZF9Uzg9bKxB9tjV3QS0ctY6xt31Xksgw
VeG0jn+8IbIaUAPhraB8sdKZ7yA6djLhyaX85F3iBY8X/0s3SOW39yzKKr3/4Z9VdMlT6S5NdZYm
mNlvieg2aM109hHA64x1pVsvIrzlEHae6qVHrvy2E+ndIEOXEp7HG6UB8EVAPCuB+XNKc+1XVoah
hCxI5EcAZjFCd1qB8m4yL5LdjNug3DxXkGOBVHrFE7o55NRS9WTLc5tS+ZycbSPsocF/y6xU3+US
4UYpHHZ/kAwv+HjPHmqWgxWwlKCDjpcPncfkv6CZrJofUHZ1sbp4sOs43jKFkM/s/hh418XCg3ci
iTSGFA1w95nbPirrhE+StTwLkSCyLiYxD3DrSXn3Oen0j8+9UPfYshie/nqIbirCmsgbaBn7bUpP
/WksqCh2USSvQYmkUriuZ6lH4iOI403Q+WV5tHBZ75icBIjGUiDrVPbWXK0qDX3o6j2weVmQ/9Xe
KK86CUsViBrgM/I8IQ3d2rgCgugR+IIhCCaHNTOI3Lrfpy/cln4V8mJd2yx9+23BvjGynCjrNWm7
2OLkxv4iwGhygnl/SEr/oQTMJ6VYYkiLnGeC/0qLvwQsvoN45Zf/aDg3R7P4C/PloqBW1jQ/a2Zn
miDspYBg+YQ5DOFKeZWMm9/GCfz/SvAicH+Mr+sCY2tmbFiUpS/dN7iiTfR6cq1ouPdn4dO5W5cZ
Htnhwln4c1DALgzwSQNVBhGRZ9vTHnNe3cMAgtnORSqdeuM45CMmkdfW0hwo6KNAhFLoZgNC6651
jHuqj4q5+wLVq5rxoc1kvaenqEPFqIhqQKpPJ7dTFM7GiZoJtO7Xs57WsNAoiLkezdYphDo07npI
KzmlfRxuLHSKQjG560FmJevSZnQdCcah1mh/uowNOsGinBMlOng5VqfXNO2JfrhxpMtxx1d8NIr9
gNv08sB64SAHzmMQ8Jea5HH+kfevRG8CuOd1LbE52QaJhxo67JXC+D4szhrtMHZBaMExbrXDgbEW
3mdF5gU8MRtgf4G4IWw46d7m2p6zcM4fEalCKPUOyxjJWsUiXAC+zHjKvrtRmS6raTncGg9dBKaB
pKZS3qdezp14Vv/cDwqgWJTD5fLeiO/2nxnMaRknzV4avVdimL6UZsiOxtycpbnA+kiXBeCr+VG4
euQqZIbumtfwja6LYGIITNVu4U4mlbtCWHUVf6TOWU9JUAeIXhJ/UqgkCoG+HVsBmLmQzWEGuEzG
bXtn7RfVn7k/o9oK1HpEAeLmZVCnJa3DJ2dFkLsRY69fqjr8ISLgfP3Ee1bVES18OrTSV4e7tC/7
heMvS+cYBRE/DEy+P4UJ2GvF5eGibJufH+KHdpF24KpDsg2MR3uQWx2Ud4wgIPvIYb+fLhwk3y+b
+52/pf841XIHxQYFrNq9S5fj4BfL+mFSNQhtKrT+qez+TghnOwUFebLSMRwiUghOl9V5b9PqRj88
eiYRbagCg/CmJhQAKUsIHyGc8oucZPDq3fb7KOCSj7P29m/NMfJL54/sRRYTIJvU4k7MyAMMNhD/
ZnoJsUsHpRMU/SS+NcITo6623/bXFlFQJZozI6dZ36jp9IjQBBZbvz2Q9qgO9bPO695HntcLe+WB
PoovJmiFNKWqbnjjUW9fgx0WRO+opCZSIgymRGvXrRmP7X1JoJ7eTN+0IyUa+wHzRoJ/0xLr5mzT
H08NtUIAqDRNyj5SYXu06kPLUIMBGyBBc76qMgQqXp9fEOF0Od5MKr1EIO/pP7QYesC5+1RHKUmB
6GkdJRcMJXj/VbB2IAieb6T7HMpiTnohDkKhMVTRN53ZS1ytjoRd9EKlkmK+xLynNHaYZLlY4xmc
ux5S4bkc25GcRBo+k3aXudHAarX/u/jxwOqyaLGx9Rkej+zrrl64sOTj7hApCGGcuK3D4aK71acl
wwtOaZwb+EZsRdWkK3aGCvIYnCoWMD4kqTray1F50io7hhlWyMW51ljAAJIRKKw2cWgJkF6AR6/N
w6EHMR+eSfL51HwLhwlyBzdG8N1T4t6Lo6nBw7TL7Y2WVKh9uhMa3AG5HFqj69EhYfzHDKiFpnHi
U3mtx43DgCvS7JhOTDnee/jzbhw2aSu1iH7GgOvmOY6cCmcBxyf5GnLqSoo64KJ/aNJa7HkLMYDI
r01PShxzPpvxyqvZV2guecXclqNCVHDa6kDoNsvK/Mouyujk6hvxOPMqW+DN2IXq1U7+emU0tFIT
y/iiZs3286moLPHqgnAkxjhAmqRdEvEQudKqrK2CjdXkZpYoUS7ESeCMQhMOUqes4u30e1v0NKOv
42LLRujR3EJdnEFPrdCC5ftM0vPidj5s3QvfmmUQHECQxV0O8Q4gvUUDGZoYDfH9zfmceVp4PKlb
oHs+ps+T2vLJOFlmiCaqT6rtgEFewVdl0uPLHRlOsK9xPIaXzYciHuojYLp/irXKbTKfZl12GjH/
WRfQ9VXCQjqDI9vv7+RGGu+wNaDgh9gh4nvgqHThWkLhIbN36gaBkRN0zDmHA4pUCoYnNw34xN34
YoW3x36RFWzd0cxXrm9t8NwZJ4mbntUUgEo7uMw1y8alvZ4vUbAyliQOFNE+yhv2EejbVuOH/I/t
nX6CIPuoVrTrzpyU2VXZYFLiMv2clR8XXd2h75AP1Ah42zLZTHgJBoYj+FMFFIInS4fmnbEmlTgh
2Ki6N/P47SIzj7tDiVHPcxKLS5RaxhsoA5gMpdtvuG+deXHJF9C7kqtt4L8MO6ZHokJhjU/V6g65
7KdB6K1ysKVxDGA5oXf4cGC3JnEzpqL7IOlJvjfV7uzuvp/6VG3A0Vuu5Z4NP5OlREtF7KplIP2n
IyFFdz0czB1CuyX2ybnIxrgZ6x0rGkeWMIRQ9jZSC7HvL7FKdJm7vYp8XM6V/6X7fFTIUfSoyHZO
wkWDyPYmIofAm5T8RL3aUQuic8R710dH68P8MWD5bAz0pB7LlwR4MgpRFTbz2i1FK1XqvaCuXtKc
GPbAmtpWaUQyh+sMqO28amAJdQjd2YDDxM15DZs0137psiY15AtEnZKCA7pwED9tMu9SR/m7zxN8
grdXbrymLzwSpAPOSO3BP7tnwk/APX2SQ85A5+axbm2j47v/39OAtXxCVU+IL0W8A3/U+wARVOAb
VIDosuwC/gdO+sRDnUrjFEEAge/2ZryI/yDZA+aYe0gWoGtqedkfgeo/iooB5DyUpcxGv5JDsRBS
j5hcnQ7A1pJPLmi5bXCQQ6uVO31089J/vhbuM2Kd+kZ9dZTlvw2OXhRyWxlL/Zq2yfn4f8iQvnBT
7cOgpZ/tboL2wbjUZ76nyizuPITzrIO6uPzFmrkzoj6vpgOGUDrBz2H8+wI2vqxfG1Ghl8tl+kaS
pzvVWHPg+ZxJP6O3ULQ5dktI/B+J//I8aQHcgowwiS7BdZZ8aVMT0OpqMpJw6j0N4JylFHGESJ2S
5OVFlB/W4imfn3Ddefj6Fb/4g8Zjo07EbeCWVpcKi26S7EaItKTs+uQvK2rld5ReIl1TKhoR89rb
+OWNQj0ABzHvZ+jfnGnu5X+4XxAPwpdamh2Tp52rXk8as98a0zWUkw7IitkcMwdg4Q6pMiFatC5X
mXTpfApvq0E/zQA9YUuKaIMdE7srhP8cKRK9GJK3dLG1d9t2XlBeG5JvywM0K6mgUcAByCfahldz
dWr7u5lx2CegNUBcXOzXt51tVGh2IzcLPKb/SQU9D/T7T/cecgOlgG8cnY8pGJj4ob49N6BdPJUD
bmWqp8ET1kDJ55qB+Ahzymh7sF9oab+FVqmS0UKn3tmOrcn+fIfpaF+YFx2P7lclOf/vaZB03KLe
c3NVIqDbsvMgLT38jUNhdtvUeECP86eNZGJVmX5aVQsggv8oU1v9loVKZQZOsvsshg1NFYXuli4W
TsdFjKo1qePWgV8X+ZqVqDp7DVh0YRVx35IdigoI9GuNz845DRoi5H1fW0zE6zbit/W47a6wIizp
1+yG+F2D1K1vJXOvezIj6uXA0d1iE9FZc+Dxh3lUsVpC/2Gnw9yW4EzQWngHYTur4P7gqwC3ifEx
SRocFjHUWhnIpf+9CCSZ0SugWeS4I5yvDevCEj4Z5WmnU0tRbA6wpXXPgu0/ozf7VDKzYMUHsf9z
eLbRJf1AuaNKrKTTCM14upjbV7mhDvTRVi4EbRMiG3tpS0T7+GhV3iuvMNY4UNS5xpZio86A356U
C4yq4GR3tNwJehvJ/PEdu7O4vRTQRbez4uDK41Ts4qdut0v/OrJs9c8+rO+MEHj8YHFIpkR27LKN
CSkVVPTmBfGIkZ6r6xzxThSvAd3PmykVfJm2jgiqobOUQy1DzwThngxjo4uU0CrMogu5wz6M1dwo
x2PyJWGYm+8kkqKpgrWp4ckr5Gy9+EFHPKKWIrpasIvXAWiEtJgbpqAorD6G5OzO/xK2zNg1xsVA
ClxYR5ba0+Rv9tSCOOMfI9Umi5Eu5ZfnlfGFSlYSoTcPL124h8MPoIfq00aXIjxVEM4fXbnkDPKW
mDj+kUwxmTA+ki6vK1EBU6IoQRrbcjF1DPELXZNP0G0ZOx2er3WLonOOT0QlYcsqHCdUzlx8/li3
SVya0Ywb93iRBD4Kp9ynzfY+8f+iQu2qJ7sLwaYRsC2dXlxkuyQVkuttiyq935npWhiLQDh1677P
u9KFO2kiZ9iC+e3a9UnM6LhfsL8gJjt8m+TBLrWbavcbQVd5vqkDy++Md+MkasbCwDvg+v9Zl84P
/uTKDg9ciZuRC85x73qAZEq7wEVVuJPp8behTo5nideRJtFAtt6/2gDPYHdI6YbMrTpdqWLLy3Mg
lIQt57fjw2w5t8zHgRD2RONs6rl2TfY46cLt/WFXREtSTo/VrA+6QvYXNaueI2Hw7UljJ4rg6xZS
WhvY7hXjSz+VWAUzeRp3qCKTksDy2HYpkXVmWCJ0AHUA1Q/7aMrGwUlE2M7wt6govTLoHjg0IDT/
a9ryKBUpAHtIvY7gXI2yTH0UMP9EwzOuScB3H0MhR4dtYilYe2kJK5FeZoqETaeF+cCqA4h4Z9Sr
ShHoHfBfCNybn1gEKkEOwOe5ntKKr5CAO784RabdYS7+jdE1qVKAq/a6YTeXBCup3Yb322Cssx58
Yx3jzwKGWKqcJILr/CLAmTCCkqwgPGKwptl0cS2Z3T8oN5QVO0zYjnCbWVQWjXehh5mZTBMQm8kz
YupeGWJ2MfcEgcF5HSlrtilkf2A1mjCJYsh2u7lYpiKfRb/nboRThTz0edS6ApFH6rzeeBz9lmq+
5jdKKGmNCTltxYyZSCw9NYPi5fH9EsWH+u1xb6r6esQZWiBDMnSWMzo6RRnsFixUzjU6PQxG7tWN
8JalOBUt+vVgMA1x73nc//MiqffPrM6xgkl2GzHKwqFNjZjayprb4ttqWCVgQj+niWsnFL9IDgP4
9fWeJHtyJmRZkkvlP762Wp+eG3RtcgSNMoH2E5zUR0AHtHFocvwz3q+onDtMI49WQzIzEWOIy0ps
MpvpS/qVXzPhNthqBuQsGIpn4a0nSAzRwFovjb47BoI5Tb/8W2gNu1hCcdagfstTI9RcDM4DBCB1
rQbKxNo3R8EjNHDXBLRlWuQSOGk/5e9gKuzpwY5PLqhqX+BSj5YACJAvGMDdZexKI0IrBemQJwc4
4XEGs1uuHISkhYzZwtb8LorFBgDhmEf8ONAPwPk2NiVwOPUQlUcMLkCwYFvmvyrx72HsNHt7gv+m
2M0DREPhYG8NPT4sUPvxF7Oa++szV7bzp98YWFq6xKlBmuYab0Ca0929Stm2lJUvCZERxM9OGZyH
+ITg8a8pG/mJsj/X/UIPQkJH91M9mF+cm5UC/PHt48yBh2M8ouyqVn9OcoHV7Fx1Xbh9luOmB4A/
ziyySUMlbfZggvxF11JXEvoxY1MxW/nAitM/Br1nUWfzbh3JgR6rwpyYm3O8urQYwk4IL5zz6mBV
lXMBukY5r5BBBYUEmwNzmj9tNCkcPoBm8BjdrpEIldsRPwK0yeDyoLySUUCiEUDvcylP9MS3Mw3G
0Kben9BLw9AxQVfRyT1yZnFvSkwy0Yvn6+lRLpF7xx3xzUdj9bs8VcbZx7Ei+Dc9/7sZq6rD+AfL
l4I/QmiFc7ma+NR194hse0oZSSKyXlA+oxrVNFIWvNU8WEyvWI++PZb68I0JyFNoK2ZmxhitcB7t
vBov09OfU80BVuTF51qyT0mHFvcMgJ2BjLKlBJDaXKKO08Z+OnRDIsKW7o3t7F0tJ/99DdDE+ngg
gf87Qj9w5IuqnWtxmwebYvctmUfDyoTCbcKPeXpjPN8kj2bfMtJsO0j4LOMP9xZV6SD5rlBx5XD+
oIE4Gv9d/GU+AQS5C3ZrakZQovUJhrrbd4H40IEWnq6xzKyDiBM2B0iyby6P1v0MIsYovanTeSZQ
RrllWFL4KN/0UXvHB2++NIw4NoAIFp4y3b/omHtfco738BEMObIE2BzWziqiVW8AoiF5ZmX8TS6R
ZDvK00AJnSLjVCy4BDR5VUo8CMt6Vl2KR04lGuDu+fIr7mS3fawmIIESKiaeTbs4WCkqKGA2Rm3K
W0LXgsW1QxRQdEL9TC8IOeOWcJNNg/kApBBQsPrLOSY4aVCsI1bmp2ZZxtPMKUf7ELAEPH5dpZAZ
qsJ/KsY0BML48OJUqg0IfRnL+ECdbX8SxQ7UciHt252xyk/exRMA0xjSNY2RL7eMIkfztKMkmSkH
/Grvv/cTeCKpwBvC+wRGqrTiQqkP/vQSa6d1B+VjMERIe+vLvviRMK9Mzhqzd3zFQLdugqNMim7e
mAW8tOnXUw2s2RVPtz+/Mf1n72/mJ0+xqv+2/BMJH67Sb4qF/A5TfHD/8BRp74UwyV9kPwiWn8nA
mMG4U6p1sDRDuz0ivcSPD0pgYL0cVOzWk6GcycHfzi4oQ1jJoXvX4b0hCFuvaHYxUGWrO+iY5hFw
0VzRuthhiBTh0sBA//RT5KNLDg8sfd6SAWf0saGfJr3m7W57Kcrf858nEB4b4gQe8oUU6dP9Mm3t
YLVfQkGAyJY4v6UJgzmj6FWxU/dRzc0CNg/S9+TmaeO85xbdJ7Oku4ygXoXrrgBb7Uu4hYCitQvP
fWnBe81rlKQjyprgCfE3a71YFsKFCgKBLoW+7Ucg/4I9qkgaM/u8B/hklwwfqtHVhgFnYuyzOYAH
asgadSBvPGMReaHm+JK3lEoXVWv9H1Dk25EATzR8jR72+rVZNs9JS1IsRoX3pfYeioAQY3Sn7BJL
3O3R/tcv9HjzvI7yfNu1cwcr0FnELAgHfM3Hfi7garDlpip7YgpzW3V3aJHNgcnKD6pDjD66LrFD
n+LrxT26BWKD0TvolsZbUxVacAlS4oAZWN7FD/AhO605euZ5soKnG9uWPm1y7MtDeIdfT51Yh9Ct
6jMSzXS26y8BUTDpdM9gJWx9Vc3mHL1LfxbFFzjQ2t/hClyKrf5IjN0avIYEdmnvqre3i/M+sXFH
O8p/q5QbiXhxYoGJ6WHfqqnD0YGgXVl8ZI0jkQtirLESsvGlH4cUUV93owOnEYEyqIqr7HUg6BMG
t+hgM67f5xGKuOJbKKJ7Qy2TypXPk7G1WmB322Cvh4QGEwAkB4UkMe8y5+uW4hqkSTRo7y4AsIWD
YNxG5dWRmTjHFI/KLCEUD41LcIre2DVcosEn/1iJCbnJvfjnV/HB8dBsZ6f6VKBlFkBCOc84NdS+
cbCX7FHcMfKRbG3s4GapBgR/2SthLHlhJsHfn8BOrOPuGnM0utWhCk127z9r23AXCxkkFKBjzEuR
J4IyHNdEkY9YNrC4N4TlEcuExOjAGw8TbTXe0wEayClGrRltsNyYOqd6eZyKs/DDyAaWd//ypz+3
dSlSKdti7xbxMYQA9hnEssoTY8pAxU2NSsC/krV6mZojHM3B4V3g1R/BOnjkuZ+IVNPrYjQr5c38
CHs0/Oun0AttVAc1dApspMJqwOgS9DThlsRsAcbMJvBD2+tka3B0DtXDl4USyWAWvI5rJgh2fHtr
6GP9rAun1rkJkN2MRTT1x9XmhFu1DABZWc0tSS+8/c3Tc+xJSyQ5thplvcs+I/CbOBaXZ7RfNQkQ
ZYcc84baUplSAS7VMjr33nVRrh4tDe7hez8T0yW17p4xQyqK6BBJyaWcxKkgcJ67sDekN+Eb8jBj
1hkAGxqCpWFmJ7HZPm6M3Bh2Z/G902c8wvcius2PHFtWYgCHbQvAGMVBSXi9TIuj1qnEbmZc2TL1
/uAZKuzQOWZz/XwrQjfxOYMS2p76z73Mc72Ge7aKubkdI9vuUuvg8YFgSJ3HZ7fVMUSMScfNGXuC
lWx+4kocQKZOKCaZ8KsbSvYdiVV6zTAHIgNWzevIN/0XXlsVhLzbG1d4T3+gntMxjFp38ZzTNEn3
ReAwSwJvJycq6jmnIrTv7L+AiK+vJd+2me8E5iV5oQU3qaSb8La0dghm6Q4qg0oz4yd0hLx10vpe
mSSogrxdqgJu3PxUeRYqaKtIgUNzE8v1RxChhhtx5EM9JtloE4+bGCRT5FE39tTe3FZZyqlcbUh1
kJ0+8kIeVNWpcT5yrfh/s4vAH/bqhV/E9FcLsbRvEtLbBIk9rJ5AHbKjmyiqThHF7ZPCqLBlBBVh
biJzRSRaJo4mTvmZTAuZhKlaDv2hdO1NXdQLJGTYYqh9mrYsSv3Jq4FldZrt22rumcToq/C/8Hqc
F74+R4vVmpPsPCVb+I8CzUuxQVqcAhXL66vV1rPrXsYzyZ9wSWsNESSwo7+EaSkTFl5HZnzcLUPK
XAnhdNCnaU6sPRoUDieNwH9gexdNatmmEU8NJFYO5EHNE8VpG8E1JbKBz7PTEvgtXDDpQPUc5Ufz
FTp2WUPWT2j3jo3UnUgDDQHlqvod8D29G8eIsR48uHZ7pDTkHO+fMEXQtYBtS0yQqKNo6u8VfJKf
0m7Gy70eMi28/xNz5/LqoT+iCoB5MFwBUCAQD5CdGMRWXtHldExJcxPOBxc9uJo5bqv7BFd9+Y86
x18yGL0F1yDZDRIJT/S3Wqo4gAS9TngX5qiETFxNS5a0mnLo3squQYsm5NfE96kTqGh/nTHaesNm
Ae+zMJ+SRGT6Vzs29uuZd7anvlkLLE+5uQviiF0b8YotSyoyPTZ8GWQ2mIyLolkpz4r9KOXP0wcC
SvwVsw1/Wul1QlXYl3Px7sYZfsLrY5Jc+WRhEDB7ARaKQ0C4OPIkLGkBLt8y3zBwLgrwzIQSGmKy
eQcWL7YrriN9I0wKRGpIPc37h1gOz89xANY8L8E6A27ec7EppROZUL2UZdmotR7hnQM/uhWhD/RG
wHeUJ938FnBLs6K5yCoFMQT185gt9enaGZiDBOcg4SwZpXbLBaI5CD1CoZK6u1rypMCZFAfxoifW
+niGb5q4ySlqtNI6X87Ky+gAmQJJo9LYI8iCK3x0qFXkD2qcqNtlMW1VDBRgyRR+Qp99Gag42fpa
psuF+O7okcN79I8yQ+j3t9qRt70HhSHwQMHp3hzRukCqE4h0MGRfHcXC7nBllq+1c/NTF6ikwfPI
//l76AXFTgFxV24JVf/GMsU5RFC07dyXRYFhzxx10SJeoeVKzwRma5N4MjdFWOW3jG1+pv4P1Xxp
v89oS1BDJdEB0se7yU1kCM45SUieeiayYF4VjPlztWrmMgrMI55Qi8T63aa6WUZCeiIh124Zj5aP
KfdEPatyCPwZlunufD7sF14f2h9f5FiWuCLEBqtgcrQTo77MXf9QffBr0oeqJdMrXBZA3gzL4QEs
ZtOov6QiFkI59xBOltxXMZFhIoBKDUsvb9uXvYayvFr1NWqym9RyFVldJdy1wcR7VarRrDtgoJg6
o/3t/LbVVSXGGz41UcIjOGhmxAX+2ZRQeURr5x47dc3o3M1Edsp1g8z6UavsmzThMB1EaNIBJQvU
y2Xm+xkt+tNcMqRX6+kIBcKWYTjD58zp2IqY65WY7Dj78g2lfjWagEF6IUcUduifoHrLVMon7G2W
DZtZ7Pmz0JHhmUG2U9Vhf6wsTvNi61P344YT+8iFpodULP0D4oXKmfcDGRCPVLttHNaC0V8fUy7e
Bc575zVOtxU5MfG7vzuHQ0ORHBgEHo2Ot4IY1p9B9VbvN2C5QJ871rc5InNB+oLi5VulvC6rEt5M
gcjOXxsTtMmxByejxyxEP4NtMr+1PtOffBKUfBDy7AKnUvcI88S6Ull+EVUNW5A6pi+78imAH1TX
UWOJug4luwo3EjqbkL9AhfIm+ezrQnZ11CxkdZjgFj6JLXOWsjj66O8iFAUTecy1lTccK8AUAYPl
zTtyfiMnIkMCY4QhnFGeQ47tWHUPc8wNcOQxlK8F//hcuIUWSwYm7G0yJzT/maOoh96S6a2gcKxF
4/iscGHzpbVszTXVZD6B+Gr2v79HQe8FAfZjvtSoWrseDXX4zEIK+21xxrePidTOYi3KVXWMrcSJ
8wJmSehrdPNhKznAqzUrn3xKdpm9nPuTnePs+isG2zH3wKyqB1mGuTmjrMQVg36FgvZ3SIHDrWUm
nYwVLxPE/H3HCllZK9u/S6HZ/69JJoL7qmMMle7etD+mVY657YTXJncp1tf3bm4eOBW3tKxI5g3D
l2toTpsTuXNeXoYqGzXx6yK0sIwdiAiHnpemfvQ7rT9KnTqCP8mfnvUwQMYGqq8N1kXywTyCCDrX
kaWUhxjadxGh0YTguB2w233OFC0dIR6YbC/UWjIHaAO1pqwb6LZb7Pg73MRQvoRzoRKeBpK+K472
ESMvMNWGDBQrRufnqA9txHecnYNohHHMvSRaHDmM+F1XC3ges2O4ULtgKcbIT4nFTCL+NapzgdOl
ik6sMEAlcyfnA/xAIempjVwqDdPbTtIKB2/yII/7s0dMj8r1oiANLlZlPe5lppxoHTLZlGpq162o
cwgZ+1SuYBQ3lO+xpAnW8Zn70MxY6tmOXa+HmRALDhuUwG1mWmB6U2gDa86kI6Z91n0ecvmPbud7
z6AOZw0wXtEntdd+Y+iJ+YohA41kOlEAH39NJldZdUawGMgURQiTmSaKZZ6fKC8MnHTvoGRiyYM5
5lkTsJvtwbEO8qgry+yWMDS8DYItTVFp/bHkxz7tVSLLeJSOk+ti60UUbSDRNo4ghqMJg+SHSZhY
+/dDkly6ZDxSUb8oxBDw0f2nWgHIFMyoUgAr8ioknnOjWWV32GOEa0RSha+S+K7J0fiTgf2vYN6J
h7klUf/emr3MV/NPRRSf7Q3uKFLcLJDoymqf8GcB2OICddOrQ0lnapK28kWlfllaenLnkpDmOE1T
hBAeUUsfxFn0BCoJ7/Za98mV8ThAagyjO9cUea0mPe3fthbnCajnQMPsjpq7gKsOdujwPNobWiBM
9QTAsNwQN8W8/6kyrpDiQGLBSYcNGKBWJ8/ZJ/mM0FsR35rVX+3woI67lzdm+Rq0/zX7RK+2kAup
k2GVimsfAUhaAg8JzkG7Pl+6IDE642v4GuFkVV6A2Vy1TJJNLxiUgM3n3zDF/lW8ZAnAqcP+rNRX
qDuKEB4XfK8Hnb2BSyccJHRxbyUtDYmJxaozk+tlPOliKBrqv34g0Wlk0xfVhZgBLQI1IeVpd2uF
8ehRwd4evt2fYHgzdILawVQGq4FhL/6awrqPkLC/NsWk4exaKlLH9a8xYRyt9wZJOwmxyW3OcBZI
F/H0vy9hB49CQe48t/L0YPeiooE43l+DS4/xcqR5oBtYPgwHFkeKo6JiJ5o4ZYsgBp5MyvNPTT23
YA+nwSbpbEFf2ZClZ7We8SWiGpussb1wV+UvQGcZlnhOaaVq/x3ejIku7VMU2mnllOsIqz6Uimj1
0v39MDvjtuKQm2mEYFih86FEpGMGE7Xb8Fmo/8jlH29oesF/sJSzmRBEb0f60G0omjx7AX6jbSbJ
EIJHZlp9h5v/wktul7wiwhm65KtY9gOpLGH3XRrwYmEVgmKyhBQU+maw/F4a/9q82W06cYAiB/SE
oTj4K9EEFQ6JQ48eAdQqp+gxy7rn0cMD9bF5avyI45dQqQ+waWZX56odhB9m8M7Uh8y/5es8pUhg
FDlu/wn4nC/XaR8JgqzL+xFteuB8HLv7mbB96Js68pO39LX+sXZKkI18yiGbQlPmoUE/LZ63sUd7
c/8pxJME3uHyvemrBb/UhGHCBAG22DjwWwS2zhBuYFgzLCvwVdkCAGZ95ivzSeKSv25mMnXjg+Fz
+lV82H++36JgnXtXRbPwK5CFX0uaMI/NIFyRE5oLzsygfMOwt0RDaUr5mgykhRlSfSYp69KPoPQq
R0eDtvVtOdp1N3UXgRzA05EEqA1iRrO/FFzZed4Gr/GiVCAnf4T2Y3Wn0/YFpovVx9ZWTETR4ok+
K7Wz1R46Ftqe4GS7krKIbqL/8MHptq7cB9KlbApX+zfJ+eGQesbMdQtqWGIgqFPER8w+26lI9xYL
KZcaW1yCF12maSeOTyeteqjV91PPT2NNz01ZW59gs9sRl/6JIRsQx4P9zxUFAQKWrKlNEK3W78We
49UOJ+T5PTQL/6RJzWX1fTa+0LqL1/BO440QMlcWwxieZ/aq6wyGNP8jQdSTEHKJVvJ+KvLdabiC
cqPM7PqStbb3AAoho9P1B5Zs3urnvJ8QIgZOFEbF9FEUoCCevgTCJD4siKL5c6jB+sn3Mb7OSrh8
26A/qsSmCmKmT5NWPcm2lv+uQRCG//xGiY8+zjxaWvkGk7oUiMj4hjK+F0cnxFJQXKhPjLvVASLu
b7xxdwvd2qJjiceHe+vfLTAgE+nPQF3RMpaMs9mwtETIJDk5pyX8p6sM/JcJBvvK1Ot/1/c1kiOP
HaYfPv7UAzOojD9+74CwWj4R1/YoRGbd6jB+2El17wLJ2Dj3A3AAj2HWo6S4hd5ifC2TQu3FXaZb
OyxfGkeeBJg3o61PKqKWugIkjgoF4POb+sR/DPHg8eb4z8kgs4npFEmJnlpe/igq+cM34gfeE4YI
4VH+mWZ676dIW1s+5ivaVGIzL/nJjkB4cP42NPzdKdgkr8RjcozKvRu+YOVLE516BNB87trlLrfY
y3gCLqk/FBtMmFnDzv8mK4pVnLitsVwtoLJeaEY+lX+gl0wy+VbGqZXFVPO/gmbPM/kK+i7tRFH8
tEPnP0srB+JZTfkrSs4G5ul0D7LsWM9t16ovXoOGYGVfKIU9bOzip7n5HqbnMuEFdFihKydLj+vb
KRFSvOktTTS/egy1lMfO+CvaE9xEf4Bl0l6cteJi+0hK4wdcHNdPEwUyDSizmtMrBwLgPxSIpOMt
9iRp1F1ZEbbmvR63evNNRX8iOqTLfPqo8K/HYtJ/kkGWil7pHKvnIze+kONhQSC8NaAzmmSeIpsU
Kf6pB3vgVnIF6eJyp8iv3HFF+whr/9qWK2ErQqXXbvRZsZX8X3V/bUE3F/BHFcgqW+uGxYDtXz9X
1lWu5dOdaIqq7+MLZv7pOzaIk8M3RJaUN8mtwy+Cn6w0b0fbolvMRG5BLpjFGhBpAFD1sdZ/8tsf
l5B7dzgoMjazYu/2TcvM3qRLU9qYr2SuHlkpztSRG4PaOhP1h9hdrYcHDBd3uHEPXDcYXSmpu1dP
HBo7n3jzzhrep4NS2OGXh2yln4LkjvOdZs7l2PzQeft3ry0b5SJT7a5uwIdx4nmTQrzkn0vFDrkn
zcG4LXJ0XIrRtpIurNRW708qmVi47qqHfSb7LNEe8TzU761oeGITT2SIzavdTsTXaOa/71KJ+eEb
db2bVbykpRIkwQ+gG5QGJ8pjR5zsLbI01o017BBBSl3A6OTVedDFAmFiRrOvo9tUYZOQAJ6zb6sF
DJr+H2l0inIV3ysf5jn6x4uVQE1xSDnIxR0+NM1f+WMo18IIzuTejTshkdk6qngvZCzsWLoLGcWi
AM6NxdpgvNi/NPdhRukv3bymHaDwL/8TkI5j5yhjAHeBAAmkBzA3oupJpvJEsgreaDtsT9OOaEXB
a9B+BDVxnLhKtpddeIm5qbNYsdCwtwlLHZf6RYJc6ZZZJErKh3TYGF7ZUkBzj1nTa94Ohp9pTjMZ
ieKj/l4pBnFn7uVde8oR3FfSG7QoyBtvWRhHDg/OSOBCuSgs4jeyPgsAdWf75Mr5HfUufUWMabiX
h78+Svy/buL4rP/1jJBd8+AB4tNwnzTkdInnUXFQpF3JV6qGY0FvaSWCyscMxjYCvbGmroihHw+A
s4HidNjFESJHRXf6lHvLNcCx4B6QmKPKbKfFPMOSO0NPxOYX3/aDyYz+3YXoiGJqE0cIZlSGzZkQ
g4f3e8sOGwcRGYOTGR13cqRraZhnDnqPXfOCMJWyGm+69SgaO6W7Yq8R4j3+KbKEW/wIyDjfRhWj
B2OvuTkkyACkNOiga7vczyDasDq9Fzz+aWwvodwbLfFiGyo+60G12CDNzok7TkgSdmOGOsy61Txu
txl2Amf79UJmo5OBIXHvP4mVC9HgVVVlkYBbmPio6m482kBFWXQZEDo6WX1Jbu88jHvGwlCtQoZz
gGybV67vA5i5GABNOeJq2ykWap/LCrX4seY8VNAAb/pQpHOLTiT+qzGBRE/iql5yGU3kNzyl9RFL
oFAl0kgW2nomKWbJtMau+uc11jb+lo06Ctj18djdO47B1ae81rLjAB8SloVlhdKSgFZ0WhJnctFF
TnmOhoCnkrcvinhC8nxoyBPsvicNw7zu1YEVgloqxXhADJ93vSGpEKG8hD1/JFfqSEfV88agpOLf
HEPLvCchfJhH13SeHztW9RwkJ36pVTvNnf1ZyyvIL9Uy6+/IZ9fK8WXC6mkplhXUp8TO8/XAGUOC
Gye9DAfCWV5nHULvv0fqbMsTWCAnyquHhZl8a8kNk1aD5LMbv87dQ7cB5s0XVLGscSdWWrIrLMGQ
5ohZtgRO1wW9dSxMzioYl+HLpOxQcx2J0N66k081ZUGMu5PloXeeMvZqWc721B5f4Yz49uY3FCj6
Z8nIVyWtqGFQ4JJFR2FBsbJNv/P1dXpDuxKFgeNW0tfR3Ihrqpl5TOm+TP2Bm5KmSAU4g+r8RX8g
zIM271oPQ3EhMDs5Vl7PA0tYvej71YZzKpcMYD98XPoRNTDHGMDuS9vBu8A8dX/XPNKZeA2kDmst
6i6hJ2J7mAhuqRBOs+XbCYng7diF8C5GwivOMRRG8E89UePHrKCoGhL4Fec4g3z7DqFgIQ2siwGG
S0nku6J9UgeYQ/b+tyRlB4X+X1Abv47nxN3xJMs6zQF+HT+S0yASHJH1r82qctdNvRYBgJX/uuPk
kPVyWC/D7hjykSgrT4LgLw3cvTW2HPm9o0FN+0wiaTH02oXtOWTuP9un0YQhCrTiOcqg2VQTRFHj
C3EdDudDswQSARYXQnF7Avbqa/FNS4n8LmMz1xwQepFAy+C1TQhOaU6JIlbir5gQ9J3jcFyXvVmR
BsqbjFP0wEELd2YhenHKLn6WJmAatDlOS0+SF286OJp6mBz68elj6qbCqO885+psj8hyQeZpuGlN
QNZYB0CeW7bnoi2MhF/zOYnVEwzUT4LPdK/wuFCGjQqesaDgjFRKBqWTVUBRDa4fY1EGWgOJCk8Q
QuZR0JfqnWcwtUc851rJYCaciAoGQEzSz5ul86H9wqBZ433WhawjaCHO5KrHP+d26tn6NBfEoU/U
DI35/hFMAL58ZBlBBvaG7TrwT8DWtiVNDOLpmEdUj1UATlfoX9zx5LHgwa8+Oujh0qAyyxK2j7hD
QDALrrQa6ic6F0evJX9fKDiMjAMOpwIQiG4ZJMHY33NYYWfMOTmJvOFONcPXk8tK4SqUD4C5DWea
6jc7ue6obWF04F7M33OzQWmQQdhu2CvNbB876Xsqhfe8eS7cAlS+1wz4wKGe+0ft/q1vH4U0Dd3B
9avXvrQBgLJKfhn7JnJPcGrnJroHndQJOZaUwZ02wqo6dW7LOmo/tz0vd5szevPMu6A0gDofyO+W
BlciV4mXfvyznjrpxrg61pm+bnW+9XrHJWNvieA0inC8fYuvedDZgrTdbqnkDqBT/mJwDB6hZcbr
JxhdbY2eoJ9/fiaNAWU/P+0gRAMeL6PaWsEoNz8JYA5Rp1xoLTJe+nXo+NGoCdAV5JF48tQ2PD+V
PRzvEGrSv8/ISoUU9OO9KUE74ges2yXz+DkzyRad/diAupR3SglvOeum7p91okQgiVY1dPTo6068
b8ejvnnl6Tqntx5UnDTuZF62YHTfYufCxLuSBJ0UoB1v9gSvVZjUsoBwfJOGvRQyBdgvsZZGZgVI
+8KwkC7plv9yGGAMzP45f6D5CuwtXv2PSiCAYluKs8o3/4DTNxW+3mX0zHqhOcg/hOQBOSPx7mKl
UQfff0Zm9rFVD8oqIwKtlbfMD5sYw5baR9f5O5Mzsj33R1pHmPyU1s8BZfb4rfwDTSDi9qYcgPo2
bByICA9djFwAcn99G0rnfwXauWqqiWKJNca3/YftF7T88cky9NRDQBdzzmBOT/a66dehMjMqOZQN
YK+NqWO10Ks/wlb5eJ11quwVGZ9SNsU6HdXavj+d21TqEFdaHnyPJq+C+ng1iKVEyPMVVx0S8Nkt
iwStIfyeuzGYkbWTQP7Uigmw7oy64Ly1232gsRnAxea4Yp+HP3nJERsWopj4o7MGMmr/0Sicby2K
Iswr4CnVpkis1DD3gGiTx4TXWpbgLA6HfYEj1MD0x7xpXcup7fY4rB6i9cdd+mXzTBJ+eqwx4/k8
+y4BNZwte7ehsreqpjoA6JC8cPcR1apuMlNnVdNwZK4NCNx8GBUo/lQqQy0DzQJeDzi5ud2KczVT
x7pot+wbD3bmZ2L/86+GoYkopU28s9Yhl3GwXsVkVK5oJTzDPkizO0ryMwDO5arKoJAJ/w67Rc7c
IWAx8O9HprAw3gcD9rLgQjjt3ffrYL02Pri66/Qy1FDFTKICjKcbhvrUGqOkIjeBAT1VH+X2nx2q
nHUCISRghid5aB/aRKgDwxQwG3juE+xqN1m5UsavqblRXhaerDMHlnJCU2oBV16x/kge3/0swzrh
yz5KQbRekiXxOWVV6TYgaewMCQ+QvJJXaexUEpj+cAd4gDaAqrtTX9rDdt9otWO+ThByeti/UGBC
7ipyMs3zBCbzuY12v6R0jXSyRcmdusDyh+rJuVMbuBuZPyo/KTr16Jcn19KcLYUp8kUVbHSf+Ysn
cPSGAoyUdH7R+9xy/b8tqMW3b2KYDpyS3mHi7LrfMwUa5dGbDbTwRLxH2WHLQbogf66oQYJZW8og
N/SmChG8SLRS9gwLppcimCttRxW65n78wiUk8NEUS3DKJW9zcvHM+I4YQ4NUCDuV1npT2dddcCFJ
vcz28KkFyG9OccUw1h1Z3VxTfY6WQhkBi8ctzaAl6pus9EskYqTSt1+tdP/ezO07uRF3JrpJXNO9
ZNqhCfyaq/NBe1RzTYCFDBEVsAffHKPYq1Fsxs5XeQFGRjuSdK3UibjhM8+JY3AjAyWONmYXRPc+
hYTOH7PGE52ZpUEuGWoA5y2cnwgylsvSySosQj3eKOV3IYCUi1Oo583siUgT6+emn4POwLLvOzZS
AkKePHsa8loK56pjk0XagQr4DX2+m2d/ah/ONCkBFoPK5M8K53BEugRGh4yrycOCz16aFBz+MHqu
vd9MG+C5QqbHVwHEqkfMis4bAZTaq0UKl9QRGU1JlbPexY0GH8qIaLPFSaIRPJYVeJKNed3cGrff
+aWAxsM9eho/OvMIOYR3wa9eKk9W31AtK6ZvypK76wqMdoTVfUIXJRGT7tvDaxTVziewGtlO8BEl
gZUhQ14wE6fwd5VwzvmSlFva6E79qc/EOQixwD/bxT8U6SqByW5o9Hore+O+ts+in4CmqONKrlZr
RJ15UvxJEtuSGG5RQ6VRz9CLg+xl7lL/xgia+8wPTEXCkvyrd7l3nSP45eWKAJ+x0K2qCfSkBsgG
yFEOeqXbXL7Yn3E7VsCGaqweup9Pdit1ihSeIXaKi37PuMvyD9vUzVIJafPzPjHixyJDOEdfZaIv
ApB1kxz0jn3eHIHd0tlWjBdGuYNycPzlrk6AJ8mqN813cJF4nc88bYRNIWC7tNcCR22xS7a9fYlo
mEF7mozmkZbOunptGYc3IxUM9idXjegfdretjRyv7p2TsKgHgDBXZjZBKAYl7drnfX6po9QQlCrh
5K6+YtuaCmTiO15GqC3TjExoV5qUXk1ap5f4jWicKfCW5Um3lEoa9qGX3WhAuz8Ddpg0RRe5E/xA
IT0S1ympIm8r7N+3vdQXXMK2HMhIhungZDBhSB8czVFv67sigUxceKhiJ0Lu47r80IPg7MZS2Hj2
UG8FA3EN/eWtai3otsNHN0gbS40pt61M/pdsjMichxjq86lxFLhT+/q4JDG6BQc1tYvmpV2WRcIg
k5x7ArwW5ku9GDjhKNVwxTCnGtYtSKK6XoQk0FM/4Fox7B5TwDCV6pVIi31awnaP2Tw7jtTEpg7f
nTpbECgkGxUyslBVcz9feJc4wDzvCCVjInxyMMTTs53q7GCU5li1VakAFoRIub/6aGL5YjXJTbMF
B/IQ/1koAzP1E7gOw0pYb2K2GTxVssrm9qoApobEzCtRt7GECbIR0hOHgMGXzLkttwOODVxZeXfS
JqSPEatFUpb4DDWO3Mro2zrRMz4FE/2l1W1nFIE8Kf92n018/XNWopkYRAIBbeUKYHHXT7IyJis+
K/xEe2HPcZV0+3B45kFZPEQtsauq8EmqUYmQJcBP+i6xt0PRpa4zvHoxnDuArjAwN8xDf3lKSA3v
1NnjkFZVDu1E0hFxjT+StbMcOWgiP2bDWADQWMdwUQqy3RwqvHSuk5KhyIHjh6zUjh7RZPp00uqL
pI5SMaI4o19TlHUeNKD/BsfZla9JSlleefbt+gLfq33W/qh7qYoANFUPALyqJkIaUKw0SrZouxXy
jpHEW27z2VNaluKr9mEUvrGtGiU0uFWimKltXbIKRT2WwrMDkudsZ61xgiytkODVAkpl2nda3xAc
WSVjdWptOFcUepwpZrVgYwMf/PJzxR3kt/GM+ZpJMLJg+L5if0tfAtqujvsT/jt06IBxU5slusM+
mihUGIxOiTtIZUhEqTxEaZ7fsfPkmfja6IIUsqJF6hHQK2vSISzo2sCZgZLKyiekCUzRgXEbdzwx
Ab1aysXYRO2S3RtUBXnho3naCjqeyXNDyB1U5fKoRR4hZOFDCq1Uu43DEJQf6wCQl5aLHBgSqx1d
Zg/7dzaWRtI+tyWZQGwwAD+JRHSND4S2p4eVKcqTavhgU7qKys5TCZgWqXT9L8a7/Bf21HxKqTIW
UEmZdqaq64Eden8n10YZvzs30vXP/D7RstzuuakiQtmXhGjsrx1xS616UcWEGiqj5pTLgRvAZoG6
oOzfL8UTl3wchbwNPKRvnpDyq7lyMb0ftpy05aw25ztLoWqUbHEmC/TnsLM56/YP8mkHtTgR0zbV
+LiT9a/R9XaAJqGNDT5ado8CxY8k5cEQ5M8gbe39WlUJ8Iqno/IASIFxhcSJ2Si6gcB6zS6OosOB
FPNY+XqDIn3nE5UTth789WtSje5mBmyQasKiUWpXuiRqQA5BvoVXdDO2tHpmOUdx4UekXlGnVpDr
DJ6ncOZn2eIjo/5/uRpmGImIdiySnhn/womAEUfVmddOfx/dHNZn+aDpdcUU+D6FnH0DWDmlWegu
CWQFFlrLZJAURdyCM/Ia4f/7t/a3g3BV3mC+dtySIjisJyuOPCeb8fapSvpVegIonKjEAX+LZh0q
pEn7S4XdKyyuxZBMzpz1YBx1ytNuTPN0bk1bsIZMPri8ok6FBG4wJd4zlZNAgC9b37PamXvlL+5M
cMKkrXU/A1sp/h8KbQ0nkijZeCHf+TQy4T4nh7HBwyIoLotDwYBMkXTfYWKE6nP/IijkctpvQre6
GJpiCZVP7pZIOXNmjtQQ0+9svFF3pge73UssJUk/7f6JzIjaVXXrYk6akVQILpgQswLfGASkUEw+
ZV6mUEEYzWPut4RhDAngI5Dgji2ghwJWyETDq6uLqAVzG0gZUXq0ABjI4gtPswxzbVOGdPjTOwxT
8QVKRwjcE5I5RmNHjlmbZXE6R+vrugvw1Sjl+Llml7pGdieKMStBnx8UVGgyIGTHcVtMpW8MvaSd
PFcpYQgZaUsMarczDrg8ss48C/owJI/niHbK92n54GWKGCReR3sVLnB4ItiYCARXAzrwnkEqpQIT
ivadmAoLFs+ZnGIKrzHTMdA5M2wOOPzYfCspyCN19gPc9C7qN7HCV8dy5/jRXjj8wJ2FxrtwloYO
X4nIt/LDPLxoocN5D7m0HdEwOc0V9FHc5V3QPQw0/mqBGE3jZq1diHO4945dRj3DJwlr835AgPOj
7J6UlCTB2mnuqPFfxEjN4h/5zocTH/dyAXsIdSb7iQGii1aGCg7H/Pg6PprJrvsI8AqNUL/wuuR1
HJXH1HkwlpusrHIG2Eg9m4iZ30hqWzPoKwPMPMMIvIZy5XrqC9U8TN7k/Ke2n8CyN4fQE5UDRqey
bPCWpAd8a9CVJBbMJ7DMKiWeMr16BHMOPanIxITOZqAgbx1zsTH6IqpLjt+Sq39EnZZ9DHPjNpKZ
JJXqR283iG6A4NnN9J5TTYPZXYmL/21EV81CCHzRLrOt5qBM3vLOtb8QQ6gW3uvye7ZgkxQGU5Dv
EkgVBEjO/IB+uuZ7/ktVGdvq05ZjlCA+TFQTYsqJh/YLdKYhewRESJKAeWl9L0cWLYK/erj7l+Cd
XEk1nmjDSIjgT7UwVyK+oA626HSgSfZlWLgpRHBj7JKmtiuFKR7wr4JpSBvaJGD5mQqpesNjsHvg
J3tywP0IE2+mcsRWN8aESck5AI3aTvT1tmozP9H09m3Q5SqU4iD1wItqwH/8cs9iDqQqsTPjQxZM
cNXK5s/fV1kQa9FvqvLipqmAbrrl+F5gxgZFITIjiw46l8Be3auybq12yCKqDdtj17XibbsTXBay
nH3+cHNzmmwRwjXEeREfmuRSgFsEdZjJtGHufnr5LCeqKFL7XbOWuV6tgfNk/wW1SmG1AzMb6kMr
rm+KOXewrH5Suxv9pVxFXz0rTSplsQN+P3kyewiHTqowl6S8uz7Sh6s4j8SYpRS/ps63p0ZxKndh
2q9yhqHwZQ1oWKsxsdC3JAZ9B9MUi+6mP7wIqBkKi1lwvUtqQeqFK3ZickqgOB0mucGv91bgor04
/37E553mzW11Tp9qr+GVN+ZEUIamvrITKE38n3Z+H+tuX39JCMO9j8kczyLcE+744HXPkdZ+Rok+
yHY2GdV0oYigI3gpUhfjJXwWTgMOezY6OwvBO2ZTDdAKMjqBA0/fH0qSk+7vb0f3/HoOjPtF5rM5
MDLXe3DMWRNDpkaZnfKnYHAQPjWrlEQONIMlYe8biwFRKQ4GjUK3yg6kSSfOoVEQpOuzOo5fJjiW
Pcnq3XbKj4nYvJve6DySP4XfaoiHCEnT8JCwScFebJU1CYt/wpTv5GNnVcePTeiC3hS97fpA1Y4A
yP1HX+zj71s0JMT/BT8x+GtwH1qptyFmbklhzi2pOy6BKplAxXmP9tKiQWRkRCcAPJhRg1RTAFvo
wkYgMVDzVyWehCZQaZOixdv8rfeU5pR8/5U6A1gauN4CK7pIbQlqYAHNpM/YXfSG2NeVLPK1SF2I
CpE4fxeXY0sNlejH9p1gphJPzUnfzfmGSUHbMPKKI2ZBCpmNsCgftoMiVH2pa2c9npY3Em08fefn
tcBPb1lu13AzSxAyVm48PtFeF7vc8rJ/jN1prlP7zePzdYuHU+8IrTpZrYXhw+4mcCGgEhSeyTLu
Va9ipa55FhGN3R9eU0wr1V9jqow+b9yu+rD4oo9UKXBktVZwhdvOUIPmNYgGQif1JM5ra/SN+nHF
qWuFnD585i4UROm6hYNJdFBS8QnUagh7YKS1XDTcOg3rIoXPHDBU5+uhklL48xgIaAfE7oOM/zQc
4d2wYI4UE1GcPVS33UxnPBwXPfqi1GHVI3PKnM1scIS8frzTROq3n4Ci0RVvPkIvy2dmdLO5x/kV
lDkcHRqjO73ExLUDW8gpcEWnaAKE32qu+oaoNYej9SiwQxgEiM2VulTTAfAEZ3LwMYfU4KQCWIx6
7TFEtT9mnqC69fe817a0dGxxlGlJm+kaXBi6d0ltzkUOzyDli58ULwJvg4SGJg3YXxSFUMW1x5CN
r85TYBMAOkrQZBCCTB55weOxACKg5lOCt5dBG5XVbs7QKTvuThMzWRhviEP0Z08CUkcIJqLQZSmC
9kXy/VbN40zPUmo5FC8F+6fzqOATN7PGszDf80EtHP9ciDeqh6ONwMOmqbuETkUn1W+ED+cxhsCK
/WW90gzadsOJ9RVHyjRkvMd6N1U6d+a6lBj4h4Yezf0IBCyRxLO8ejoSx7heCD0NbGAV7Xg6vxS8
4WTY4CVxolAOIGTK393XNwkyMZGHkfiEfyFLsIOemee1Qy6Ji55oDmu/XhNnrWBTxSF00wg1G9cS
d+7qe3+yu0d+gWcJX0WrCnyU0gte8TC0s7aADaCaWdv52SKTWp0DD/x//CZM6gAhvcX2KfpG8bDF
SGJOsAIyolhHw6eyfJi+6M4N2mwIJNk0vaJSlYsAGsmCP/xq16O4EVoF0xBDhkHr4A67TJ+g+xoO
3HVue8TUFtj9PMCXuhORMyOP2nZOnC120I4EX+S/z365ooDiMuwrl7B4kmnAjhgAEm6z+eAdZclq
kZpWjXh78XO/BdhAU84SoOrc5aOo83IOScV4wto4Ed5dVSGXLOiV0gw/KtDZMGecqAZ0v2yohgAG
aWjKHzbjeCUiwg2hsQBQhDUHFHYuIY0ND+lLITXc4Xz+FChpyqH9qmDsHcXWBzVYdddsr60EfiSX
CvR+CH/xbJJ7ruj26aiSTpbCRSa97JNbFIbth+r1OYkFgqcKhmJ3olaReiZDo+UYmy0U1RVrJMZE
x9cBunscO14oE5LdaPKVr0yNBRlvKJRTmPM+PE1iNCWUp2m11Wzh+f9n8wwhy4w69Uv39y9jkQcc
+SQAQzw/mV8MzoE1EXa0YmDxECDHjRmShKaUjY18dYJz0zXVJJfY1tfS6ZAdQiZJc7wLrVFJonq3
h8xAPcxRjflZi9U5CTiv+QXpKRLwinZOa/KRh2jN3E5DYYc10bjmGjC/ZSRJtpBLvToAq5zM49La
XfotzTsEsj0bTGfUI9q1nyRqnk4Z0Nx9Pfo0WiX3fmGV+1NZ9yryGAsESc72hap6q5XKyq+F6E1K
nUinIkPwir4D6d5696Cy8hN8cZaOonIV+OwkStZu83b/uOYP+hGCtLI0oKj1bBP18aEC6mbAb+1X
nMroVKJZF58mXn/hVR9DLmu/T86rU5kzlIQ2BMqB72jpjfPKEEngvgEPgYgB+Lg5ieTWhJduI44h
3+6+6THdcR3DmKTQT20YvEhPYy9zs6uZXq0V0w0+OkrM7H35R4CEP08MZVcD4nXSqcsp0SpYhI2i
uZjdST2vPyct507GNLbOViSQWVmAvPMELORXLbG9rbW+SQPsEE74WmDSXIuBbbadIFM3av3xxQnd
hUz3s6HMwG3mpt1/X4owDgVeXgTcXkPLJEHqDStG1B/vC1FLxAkVJi7I5fO3eV36/YtZ2dubHJP1
W05UGAzqy7eD5GJl+xyjZ5VTdAXeQkKhJB1JCIspSUrIKCp/HYmH445O7ChTJtQq/z/EEvi/7DeW
nAYjkVLdmIXE6p9LIc+7m1d7SjUMEnlgyw64psyxVZxtiOkimHqmwkwcYydtbDjEB1wdTTMaqSys
s/Bq92W/zV77sDfw/ua7P3wrWHCZK6Rtj3i/9HNuxK3naPNl4r7tUlCEMwFtl8a70ATngStTA/57
OuggQupbAdyOLChDM4+PV6/yvi4yxWepmJ8NMIwDdUGAPf6VTUWD1bdlvPo/X3IGjGSU1N9yFoiz
Vn5RtjzagOdvZ453I37skHXN3gnJEsMHXSuxRzfT7f5M1Uj05EnAQmQPpzlEA7nVFSTfJFyIP6yF
eCZDp0wWhZL7RZcRvGS+BoxakZBX0CmJSeJQ+cJ63Pg6I6Nsgd59CG/XbgxTtOYE/XPDV8jyBkjA
jH442xxnv8dZXBjTAoP6ofjqMqAtNcv9Ekw3AwOzGuMpaylSEWjTCdHgQkc89bvfHuNwZiCAQ5A/
oH0/CKBwy3BFDxSb/rm4zt9BrcLwK2RKcEU19ZZAElcAks3nMBVRQi5KWgmQRXtkEznFaAQ3UV7B
xpQNpyyVK9VYkUv3r6lhOnHYtGjAqHffYOceyKFCaAsZ8GA0I80EluxrN3DFm8mCS3hT9atHrm4v
nDGviTAZjFATWO7kpmtX6JL5d/soONAsRaO7unuBz+jbzhw9kwlhwoav6ZQ5mFKFfQPduVnW+cXP
nv8rzWv47hIEF0LVHF8xKvV5be56xHgFxpqyUHDpWjG32CS1/VVvlkBaEnI8S88aoOSC+T2ZIdSy
2I51eOQGX6VmJMd612fMyykxi7fiA29XWV2oZ4TgtqhVuyAZFPlC+vmcMpawFkBqymu2HETsNbHo
rbmg5UoD/b43obhRtul9yb6r9/Gqq3DO3YsLsLKzuT5X/4PsPgIIz/A8jrorYqcsH2dbVgPBhCkR
YpGUf5365pNcQtbwKmZ7lnITRvX0ObF/iyQ3MKfGlrl86cv1D2V5ZdXEFZhRA9sBPvxn34vCjRv3
GKJLxRDBiNgO6BOcb30r8dw0iyq/+hIZ9DU9roRmqocnAuAr2vb8tjsnW8nhCuoK6UpqnNeKG9bN
NvpTJoap+k7fHQ1R+yK0G4x6B+kfJdCWt+KYUvPW+6T1CmfN6QaN2CY1NGK7N2iGCAJ/QHztOqQS
YI5Y7jKuhk6T28DDo5Btny8aLaLQjRHKeOncJsvLmWBMVqqKFQvXNMf5CG9q47jcWjs2ZTxT5fGe
MFQZw82ax8pcugVaYntM3wsDkcXjtL97eRGtR0JWdzc8TSg0mO4xUW72cnDyyLp2xED+kF52Gy5n
UfCbQ/wlb/SUlrS8lk55MvTEhYjvysDtDhw/xivI7EvnqQ96rETJN3sv26Cz4xa3t22aVd8xrmhL
Vfm9J5dR9k2aPquUXlMoob6H089j63gBioJWXGBD7reXq4/cpIrD5qr4WFCoQCSbJIJFbt7u8ktE
sfb4LVTFzd8MBEuPDFHQtxIU1mm6JD/NvWEGPmcY9OOyzSGhbD5D4heiKisudg3f+tq/fItPKH3W
QDe51GKU3J599cobg3Q5M5SPPMtz2rTZS/6gNylp7U5/otsWSeReePO4KO0ByxrIJgMG6+xN02ch
sXNeTYgUtdZMg2XsCfJ03BJsKcjSZ3ZcrtxVnHkedoHIVOH/p0Brtd7lSxRcyYFvSoiKUYOAes5U
bspTZJpyp9PkEEQLyQxNLAGtvIRK7zLiMeRj+1dI28jv7rQOMSZ9A/BTS2MM1465nEPgfP2WvWEz
eXeDq3NB6JebnnkTSvOTvtF72DQpOB6lh0ARA0ilx8UH5BMZOTk+kULIfTZfN5ajkZwKIvo1Vy3u
TAjpBWI/uhcoLfkymjIB71kxbN5V+aOg6W/ShOjLG3QR51nKGDlPthdi9HuIyWjssPmBKbyx90z7
65BJ1leQ/ivaeWQCcQXlXzLCbQkdXkVE9icDGUHCqkOeohKsYe90uzWuVg/WwxBKNOP5UqD9py3/
8XnZRxWET77ODZ+RyBcCMMef58ls/HKPlvShZxGVszw1AsEoyXAzZy83aMlrk/YKz/YQT1VTkGO4
KJ0mh0yK46T4UMZEEiAIAFm++MkMWao1zA+kdOxCsvdbHm0GdoJZFvOLqvLDt91aE8MCzeQZinMb
cdb8PaZIm4/bD5dQFg1eI/krrwUj/TBnG/t2+mx46wXAtJbGc++INQYf8Y/zXECrCt9sWuoWwzoO
zXXjSLhwSOzTBx7SFsdFi1juRia5JNnz0mZyeEnJWssi/ataEHkhtyTiPK5mbcUNBv7VWPOuNvRz
S2EUT1vuzQdW5uvscA8Boypec6jwgpb8xO/Bp0pF351NpNfn9MwHQkggTM412oztY1ziRbX+0NcS
m6i6YpQyXGJGyC/M5i5xJAJb6zMf1fUYu6PYUU2LYLZgD4mSDoiN6EJkhA/P1ivGvwZZReyH25IC
GslQ4XzR39v9CpZ4tWChQzH0efE/agdixWg4M0T8QYh5AanEo+h7wiByieoNPjdsfsfkg1gn3iOo
Fu4H2ZeK37ieN60gwXZ+HDX8evQbtOuqKpAFP/DJcjMSakX9511L+/Wqp+4RWjHq0JEhIwXcg8tO
g+/ENgbjzyq4MvmP9kPDkOka3s3EHhSuySMFNBMt9UdO6vIynyWHJD3XlN2I3IJ86gsuzyUgTxgz
LLtdhJKPWvNhOk3k4YWlG3tjY6K/A4KwQbBBQ00qGejGVO6W0SWmo6Q68TkCO2GKbywuwm/LSsc7
KCGiw7TPshQJpvNXzVeCZbxUe1XFiPEsVIZm1CoZsmIjQAM61ZVQeo62N6VphnxsyeUYk1udwhRb
5DVpYnVGHkn5+UPIKvKX+50Tlw9XNs9vly8VdksYWDtnYbMoWCtpqFGxX/g3OpGCKyAX/YFOYgbD
KP1Fzgc+v46JgDEjOSpjVh5TQnd3wUgW6xJhPDdwk3swolOeOVeDws/HfaD+o4pq0fNJGARLbls3
rQta+/hIn4QwTkmLaMH7m/Wi7ssM0SjrISL6ENxwlDvTIJrG/fsG4gt6Ipfi9weQtnYhKOT3iXol
U5t6/2sGrB9PfY0+XmEziar4gC1Du8hLMI9PvX81G4NgguHy2HJmfV1G5XPg7fD2dPRIck9QXMmu
XcCFeA4sv7SQ+cGKo5oYJzYCC2ZieM32Y0TJAX38vmDMGukjmAsFvYjd6d+xLKTDuCxfxSQnuqlu
/kDOwj6LezV7FVlWk9e+9Lf3VqhMmm9SqDa2cedySEvf7136wQBQYGLhVV1TzgTrHScmrAPBOar7
yfVrwZqm6Bg4foBb/BvFWzWNh4pSCB6bKK6DvIfsCyqxsDSbt5vBc0r6kXBHHSdAO8hjesRDgbMh
qTgNN4TmIENwiiWQ4U8gRh4yYl+yjEr8NGdViyoPzTqLv/GrWsJDmImNc3INrglTHJezXDhwE2QP
4vOBbXLgSLqsXPn3fBtBHmm+ThDJp5ZzchbsrxHRbWiL8wOD3leLXsZ4p9YalnUYZR2ZM0FzLD9N
qZj5eZvjRlwy0oHlvIftFzLptNsPBAzeLHZYMlbhvtJNcshUsW78v+byBL9zAbGd2jM37ylJdRvv
aBoEK4YCVnNeX7CCpbj/DpZk1DUkvQM3i3RmSyN3ncg+LRfl3grvJpWWGt3in356nAr5Dsbb/0pT
UpzACpS8qMI1GElppGpW/+gX0zy4gM4n4O9UKda4nQoqXIsAH/GV9T/fqBVZkcH0V8wU9yZYTeVm
FClCy8lpNuz5HUD80Bhl2/RovP6nEfrFI+w3GRcdBolqct/b0Jd3Tf30MrvodlZKE7dTdNkGqhrF
vB4gHTbI9sVaEhzlGSbwYXfk47cuQ3X0SSLjDhBeSXW0Qe9FQN2+DhoiDZZrzfFwfr1vtqjkSFs5
GWUsMmuHSryELh+LGSzjE/8FdBTfrOBPChK0FOwB0rFVXajXJCKtq/ofaCxiXHec0TaBXibmtzFJ
ojWeW4feGhz4E5+5ZxIvXU0gqAJZmBgpww2w0u9hgm3qlCVKd7L9O7E4l3q5lDH+7Z38fAnXpGM/
1gV6w6acl68V1KWjnIdLggKyVf4TbBdHGFTsnR26rPiebDO+MojvepNQ5XXTfx/a/xoVRU5cvS5a
7gjham3p8TYixcbFi+GzEIvTu3GOJ5Fl4EGy4/iyRfNflwwUPuuMOi2VE++9YZEKeVHMe8Izw5/q
k68t0iNijk/3AttHent4uWaph+Z4asoJZj1yN2NczbSEBj1hq2Hnv9jIuV1wSbf6FVR+7jsYndh+
6V+TBl0Lt9Ypr1U0LHuQViKoErbf/phK27Efp8qVZzOmvr728BoZPmKX3+De8PXQ9i74wH03q63D
1m1slDEoX33BFipidx22pIKPhAoWCdfPCRd7322vFebKjmR3U0wibb7PDVWntfxJG/ztB5mQo29k
Lh5MPomLYgimLu1y0H3GsZgAy6MOHdl5CwBJBaB55SWmD9x/iqAmfJfddGHctlOGpuXxdh4D2bKN
paTTto6YNNMAdKjGNb/8PNbw0V+sOwYJusEFVayjcrtp+ltdbBK1cjGqun32Am8GIFEJvt/LDJun
Ki1otTm6ftHIHfjyIckcEcBtg2x+BCmXp6howGzYIH8BA420D3LTpisTmUuLpsGxYVB2JqhjyQjk
1RFdgWlkPywNDGOhC/GuxRbuqFDdykBLacppA/25Yks6Ecj7JoTFZo1aoU0VRZo93/HGQfkBh/6k
d8qtNbNZoZpjArcLGEs8TdDscQKsfEPDZdBPlUu2dptU2BQAffqddYU577H5dZv9o3DA/WNmKJDD
+g9Py3eRis0HAgQbUOwrQKFPbQt8T/6UUaFoUw4oCsWtMdN8bjpW9Ehh3LYig11vVdhIo4h2vKlH
93ut3ch/JDaqGyIfnVnDjftvfPc5fPSdm3iNQ7pWW4PA7otcql8sWJ3ctfUfdOLy/kPnUPAwtgTW
b6GLKmOqdN6B4K8iSCt3dfiqrors3V6gkTfFXoikJOIpnLomV3gLNOR656nZvVdoEnMafS4CWjNB
9dKV83WVySD/5JS3CHwFOH8Dn4jMTjDaX8f6DgdYOZkuDti1/bfIajLDFvTU3C8rRYBZs8bA4A59
rsq1MwllBizVZvep7xPiHPFUB12zziB1t9Zbhb5AROBB/gV0CUeequx5QHk2YYD15C5c0eOvsHmw
TBduYwbrQdBlOBFmYmAJ/dMZpveZw8Iv5PwVPxW8UFLbKuwR7YK8kCSNZxPgz80S2cQ00ZPPUtCM
5Sk00YFUi8gqLiHZiJ+bGMMyv2/Ua5zTo/l2zAlAngH5MwCxGfEwWpxUd/34HfBIFCtPZwTHeOts
XZd0oJd+mlAtMncRIWLkJsRJr2u3tQA364JoB8A1/GAidgA0kXCX2ulnItlTr09oX8booUndyYUr
KWvSF1UBBna0/LQObMc3kEI/KbkOHkgGZchukNlsR98ISH612S1Qe2WiR6pdzcm4yw4eO0CrmGdo
6D4bELkLuJMCkiMvMxE7L/x9z2FyAg8Vc1qFuUJLVNZpitn4sg5hmw616nba/U6j3IxLndsFE106
SOOc6F+IcoAyP1UziyUa79wU+8e7YPKkqv3pikPm/b2V+oejSrDJgpcDGIjuap5RPdCcD5BccYYf
tKnJxG+3K+C0/MkqjxjJFY1EE7SGgkoYeCDu8OU33LzCUS8Zzr0SkQTgcTIv01eiZZidBjZ6jDIj
pbWPPxZFbDb+Bt21R32KexELlkSZTD8J01rJX7qfZxO8P5LFa/yKicTfXh6X2eyvYahx+Ch9Jm+8
wXjmhQfKoF7AtaDGak+5kJaLfQ4NqOTsRTu5pkariXTGx5hZFqJjLlbH2q/4GlrD0w4lj86eaAnB
7rnIJ7WCgQPb8JcFwqo+kA3zq4+Wshzl6ixeuaoFxnae9nTbmRvTFn+smwvsEzlffgJJCzJhgoqS
r6CQFX7N7CYTpAQoPkcM7dr9wqwSO2MHoS4uuKZVV0PxHhtnRPCtMcoxDsKi2LojJM6HSt2LiUuI
CVJMKrFx4koXzx1wlS1MRA0xxO4LzASm3a9L9QjN1YVsQjDheNyZgB9ZAOzuUkEmNHLe8KpMF7W8
ow1jkd+FGm1JBZqO2mQxsaTdHjisXunuvTYyJX1VEX2eS60zvMjgrhqvpYFy+uoZ7FK0s5/TasFa
TQK4E4ylGDVvPQrFAtyjVXGsX3b1SsNKdhgymgFg2WLgu4YZNyX3nSCleQM2Vvr7o+kxfhMidqoL
0wwAOmHVTDvr7KRT1L/AX96CyT+RqYvCwVsowI/Q3dmu7YLX13JDrcjMM8ScJuddwmucbMtI3Yh0
JjBeLKloRt/h9ANVP8FJQxdVzyMitDIsqbnhTna3UjbwwPwsyrikdyhqo6QyCoLgl//GudxQyUMv
UZ5+JgIFwtp6sFFtsQQyGjCAJBlmJHecsQnjhUsPk0w2lPTmohf/sXp0eceB1GUiArtY6CtJ+XCc
YTnHZjpjY//ddlUIVU2ywPBwTA9dwNvI2gqxvv2G0MHD2FQ3uoKttrOOzSWbXCyl1EndAZj7+HC6
gNVt8WZAKxtigV+HtRvWfnH3QJmsWNWPadtb5CmGA+6zb9oaAXgc4Me3LH2fovnXf8hcaRLJUMen
QzIoDkvocsspY6EMfWl6VEDNOpkhZpqm52aFdW2L9Uum36fwtK5mySMm7H9pUCYY9fRMrGQG/Tcv
3Dh11dVXKW8nQHCUwvcKpdWsITHFDVLb6m5zt8q/0U7xYRwSElJqBq9UFO4eyMa1UxbR4Q+SKIFr
JdxhcFwB1+d1hoq9x7I6QudkIsmlk5mWOdKRuxL8Mu6bN2ZC9Ca3fK7txzpeklGmGBwpEP3fp7Xg
r8sI5HSCuXTnHraMh71RVPw09BXcypUVaiLr1qI9hIPnRuC7c1q43XMtG02lgO4bs51E4lek1AwQ
JYYHRv8E0AWBhVOZtHUiiEW60Z+DuD5Q1xiIB1M2cfuBscvNrJ6CwYrfIM9HUC1WQTdkXS+5hi96
1B/QiUihVj1JX++vYv7sq4P6T9RR9zXBdKvkH2CdlBtMaqJoeMBxlfnXZxQ/+d4l+XqJ01uO7Ryo
44a461HCa4Z/f4uSw4aS8j7uvZ1CEfO/vf/Lv8ZYH9VxuF8TGWtiiM2ez6emYSqWmNMQ6N2oZ9w7
KsR679lqkVg6Xspym120ewUAr0JN9NLT8p6YjHZWuvnVXBDn47Ng0C/fA8yRnfjK/sWELrAOY1LD
mjirxWw10TTU3VTNRxpSf1cxDX5yGeHXh75+/Yy8ACAvWnNxd7mfFwa623NTS6GD8cMeEcLE4fl6
1hY3U0kQe/y99rMSQwi/soWRbfRAk9qA0U7ymhxxnE6037e6pL6AidjomcikF/w4N+7dgqbwymV0
jGMNYD02+d4120+cdrMuyUB8tz2JVj/ss5sOZPyjf2eWsKIVJdXv+No9bjUnrhF9DjGy5eLl6JqM
XtJz1XeoZmca5PUVwpf0oeA2vP6s7U6ogiwTAZV/i+p5IurvsEKAg3yrow6UltLQEnAG7GLaMFxX
05lvtBJxHHDd9wKw5AzCNp+ayHNLcHTzP8pComrjYeCAW1pUfqesKrFdEZXavlFzKAIePg4oMQqB
g7RpoK88LPVt7bhWs+/3Q0MgbU3nachWoFT5t20zU6U4F9lcapQ7sHTFFgLk7p3ysL6rfqTzkqCH
ym2Zycrbdfvtf5Ppglz1bd+N70mGHViU16Axi0nAKmV6Hayk3pDy8CbpZHsVhbaMaZZfU5p72QAT
so5mOZN0SQNzyGCoG/eYroRwEEMmBz/MlDWvmv1RfalG3ulDKakBLo0Cqg0xYmb6YihNXSAq8SNt
sJCMhNU0UEOUdOtl/KOMTMpMNB5BVOCYmwOewE0B97q6CKVvo4k2B3DaFjeTiZysGKcyQQZG5LzC
DqtEM7BpwBhjphT+6q/AEssIDMt5CFBrckYdpXo5RogWgtneZUz8C+Peem2VWpWC1vXPNUXfRwnf
Zde8cPh+TtR63hD5JTJJdoVk7cDgE/go5xr1QQqidS4RKDp2yfCIeopOLSFXkuUJEfpbEaghIXO4
c4OJOaEawm5qvcT57Yt+P/miMmT26e5XFqOWp3C3PR8vbUiTY2qlH9cKF93zaX6LTL//TRmP4lSp
bjiJEI3q2VnZz7+umFbKhShrjojhig1TLyIpbMDvUBjQGCfnnxw/zTkieySZxc8k2ANzTxNhuUEF
Egujx+Y7knR1Xkj7Twi6zZd0w0Un48rItQdbgO4TSITvSH0iSwtfKsVd2x5UGZPn3GspJ1vsCsGv
Ztdwv+I7TPMkpjh4x344Vj5Gl4yzZy3FT+JQg6RzT79+Uc8lQklHlerqLnMScuAV3J8cUP56pfKD
gq4GP+ld7IHXvH+TmWM1SWqlkREoHIB8G3H70AxIRvhY50Y1+l3NjoHPewn6FQxzSeJ2U7gn52qT
NfgLfj5lTqevL0o3OWcEKyWDxxAgWge5m9uSR9pwsOd//2A9XZ7eFv6xQZB+lTBvBZbQZRqSdKJN
/DP0QaA8Yk1W9XJUwl5jbP35CMvQNoJV+ziNb12tTatRDvr9KnW36xc1pUjmzDAgouc2ZtiKBdnB
dNmAnDdOg/cMfQkOdbhQuZWMhxpYS0mzrc8OUEqOjQEzw/6vNIRGEa/V1TwpS44EIabftlvYLgQD
ULQPgnCPTiRso7vZYvfiKjP+in28gg2DbBODxf/2Bo+35yLJLxIeKMOv+BrghCr5yaxG8ur/puDu
LfwC9N5amKhXu1RaN5yWFy+nLiJNRV/USS8JnE1Q5u5JvpHkag2q1d6f2e3hpkh5erKk6IKEa/T/
0Y32M3Da0RRyULWvj9SU0ghdFjs4VLMWn16b7f4wok8irzToV8XEoF6KqpFyZ4nfRdQtbskD+nH0
6aaeoZq/NB6bTqsArTtEHNmc0zUF5OHJd0vHXiMpXG32t1nK47PMTQoyht8eXxATZdfSE7PRezVq
2bRsjQFvIkiJBqE/EBMsOYuk4IV6kDR/reehTNlhZKcJdLwOQwys3ybaqfyiM7g+sLrSnnPIwd8w
JVGZmA6iK2N3rbLQYsbYIp2r3LZkKrRjrzS3ro5xEXdiw2bx6tXuPuJq7UFbZeApqi2iaGphiPQc
UMOGAKyVP7tCANYj9ShD/3J9joUuf1QVq9HxhUFf+z4VKF9634unnNK3O/94KmHWHhce58k4tMU8
x97S19U8MrOSet20AMvkMjrLO0LeY4P+sz9JGIL6FVx2cvZ1EV5uzlkdgqUeamOG+Qa/yvHnZs/b
qqQ1clXbskcTEbWqlo9ROLvKiIm4TR6EEMQG98uTCZfe62M+dDu/o3CUIW1f1Trml6eZVTWezblX
ITNcbMs2yMBKE2I10foQhu6566yhGbDf6Te3EoI2KtN7z8JlBFRpjo4qxBNYYx8GFC8eCuWXcTOy
TWFwdHvWhhOX+4kGPcpsMjGEKXD4r7er3xGCfE3ncUrXkIYSg4IKbY5SdQ1eHJdJMn+i9DmclSan
6dh8WjyfFjCkLT/5S0NytYGPKd2ii3fbpP48R0D4qWXMGl78Uuc5qS3qKN5jzHS0wu9KCvU7Sm2V
bHDsSVvNI5biA/9mpUN1HTaIARwNVmU90Hv3CK90K9gvR52T41VydIE1kZEoYCsg//A57jFRF14m
i9AHrIQyvBT/w5Pm4dvOacmrxaLikNjMoNRV8y+kvEB5bdJuq87dVb8Kn5sJsAbgUh4UQB5kBghD
bQz2GgEOIWpi9jvS5wgfJCUin4DACUa5ObxOn9ynSuoy6FW7AhenpD1DZzmCOhJgMyWp0UfH6Ibo
IT3vETTF52ZkJ/7DMU+i9PgviI45k5IWTdHTwD1Svs42FdkptBs5+2n1QED18M0tlFJHNDrGI7j2
50RJ7g8KA9KE8sjMPea/xFPYLb0dRHYH0bHIeUL8eHsQx4LO5EhEidLQng7LzkNfwwibwRCPUCK7
j5VHx26N4G8BA6CJ/XFDIufJmQDIZjoazuClHAUer9xzQ+wt+3Do7tRtq6hf1K0EDgQ/VSglv16d
1ykg7oJc1PZrF9YSKQ7pr5ibqK6fnMpJocRdBugbvzAhvqfXSK04XfabZ+F25p57d9VyT4JD5MFT
h982G5ZNaH4dX5j3zUyxlq7erRhRHLmK/xar6cjfycEwyQ/CswN4jv4hV9q/BWSPALCBln4Dwf2V
NTd66TG9J7Ym4KTqaOmiLRTwRrYRQIY5F1jRINhptsUOXAeSAqqDpbFjxy4+8Yejt2pM+RdfeIZt
gWdvQT7wj/xgLoSdf3hMLCuqq3miO2pSEWEoAjVD+OEf2b1hAsY+evLclffMq4TvOKpj4wyXWuoe
7dEtV9gFxkTi5elVgZOEcCFvy4f8CIEzsD0jII7PznDGvsI5Ka2i+VqLCa4wq/MHrFXAp8kiIHt8
9GC99/0RjzE0sZ/ez55zGPHqX5GySc7HrziIKUT5U9UHtp/3GgsMo3FlFB5OujyPkVrGUIjk8K09
E98+0RgltMBGIPFGFc1qcGbo8rerflUNkhD7EH3aSJi5ilITNmmrTaQXScJaBLwBECyNtu+xOMUx
nE3baPuB7gpJb0vuC8cymEwGMTunrZ+/hyaIV8vUcvV7YDvXqF+eqWNhZHq6T8gRU5EDWPlpQ6i2
YUvCGmUa2GyqYxgXXDOFTlP/QbWtnLMalboiO6sp/UZkfmhsEh1zk+foTfI4AKz5Xeend1i2MrU6
l0YGV/aYW0lltI05ixCx7voBx9nY/Q6Wgjd2s2Z4A0uLjeOxs2Lk90y5J1BK/pMC8sot1bqixHNb
euhfwhyLN/ZAmIKIQzsZsvBMSJn+xOUM8Dxk1g2pbUJm+tF6280JL5w1pUlQP6FKqK4/rSAD7IO4
1Wo5QVWSFAoPLUIyeUDozHrTJ3qTR/CZ8HMeJdYiVY3R1D94cZSDLLuCDVh4xz0p3hv45T6SzSSU
jshSaGL6WDUBMLGYxDL742to9Caxj9QEV73Qul23tCr25uF8IQ7iOGzxb0QmKqFh5PEtwB7PIceu
4w7la61G2Evwko0rTh/Xt0LxdJC2br65XGaWQolCjIr0u6VrwSsYDnAuz5UXcEfmeztZTLvMEARJ
tcR/zOhQU6juHgq/RIg3PJairwPIOOZOrItptRf6h7Ag2Y4TGMEqCDvFjYNIYGvXpjijfndwI5jF
f6Ho6ePvHtamuyKIPrVPmS/3URCLDcznc6zvK9zxbyKemliFSWXss/DWUVx/ipJ0JqPE8WbSeAtV
Qq24jNJt6GRHvXwUv0eDKNpJcPBs3FRUOOYUeqJE+EZ1sY+ytTqlnZkv/U1jHoumIX2a/UIV98D1
2WDPIAhHDlLLp/3Ue6jPXidzXzq+yHF7UYuOPdTMoxXPrQbl2HHqN9ueg+xaWlkVkkHupVy506vj
sbMfUGVQUNZOqwsroQxqAoJSsPvzJPrhKL1Nm7kBhXStqQWv91A1oud1aWkzQgHOiNPzaJ/ZhB+w
szrZuK68P5RQZ3rjGHQXl/vhC9paogpEbaR9tdmlWqGcVo2fntrRk3Pab0EXh96EsXWC3WATa1tc
tFVKf+/+PjCccr1m/gHmEDLMm/XyfJi6IUXxiqidnWU99yl8bwgIR4Z8gx5xNrMZA9AnsOylLN95
V/YcfZlPchekaOln5b6MGx0O0vAjDT+wtxV47BBTw/ijSpDiBF5+59PpDfbk/UpE17c9LNx9wiYw
uffC2MbJqxCRHfgZj2DV2b0cbDD0dlwt5xAxMGc41FsngDkn2scqNAM6kus/bI1rkszxQFiJ3zZb
9gHR9tBRqPX36lTWwuuHzZr9Ke7UwGWUeoK+Ln3FbjxqCtmveYterwnoQbHRsRW97xKPDBjLL+/J
ppCz0XDwTwCIfwl9+ET88mAl4YaSsk4UIl8UsN8bwlGRSuYgUNASgYNLnjmr0ImnjqIOw+B+wqD0
jxeYEpgGo8QIBhmO4IJhlq01UAcqrukEC8hq+y+Nwy3tqdawP0m9uldaGIFcxVwHgibJeyLBk1QT
bJjEj4qVue5I5et4VbebEE5QLoJRQvzB/Wzfof5chc1PnMKcra0OoRApLIQVSF1lQ/bJLjGgjQ7X
x//5M/JvxtRmUjikkwKHGwRRjYRt8VqH4CZnB91k9GPCints5Y9p3DcufcqOLBWHdBMMnPel7I7X
9R+r00gzLxGnQlM7JUymIbUlbPZ8QalM9gSv+ro5ZUafloWmnt8ofj+FAGM8twzoe2PuqdEtEKKF
PraiWnSpkU2fQCu0v2xLW+Q4gtBmGKb5++/pmdcHGJQl1kQCB6h3JY+TUY/hI6rBPR++AbBzDA2P
DPY18xT8lruVqM/brrrJQXVuwUvJV15D+zZ18OKBRY5B/YymK8y6sgQHmNnAvQqz3eTG5DoD2mb0
cfmNzbNv5NMkmllhSRJcumArRsBau8JhV+dXDXSW7Raujli1vh+0nm6gq/lnIpT1DkZsNtF3nkee
H4Qny3DS/TxN+GTqizlQd0ocf1YqXKZpuAd8nMoR0XBO0JujuCDdf/DDW0gVdM7uraX+zSnmZahu
incgd1K+OeZT9P3zoGq/qaJCriVnSjCwdAGCq969wJ8PFFPEbda6irz5gvKYIEeIg6puf3q3yK5Z
9UgH6SlNhbATlDP4tmkAvRuwPYeNXFlgkGMUkRR7/OPeXeMDaL/46aUSDpT+ie1mdObjxAcfnl1p
xGpxceiRgQERxRFWn09RhRVqj4l/9fTXxXAzreQBYSYeRxqDXlnAvtOBM8cXyMmjLIXMhSIRj02T
dvUouccvqvH/DSg3HEs8ODHSGS1j6888uimvsI4/xRdwM8d92ZIDGJzWYg7/VNk6pIVWmpxFBnGp
ckFvU9GbrTUHgeCXAR0Eouj0sdEOpv3DN5q9QF8vQZLjWyY3qpWpEhms/97WXpH4QO4k9rBo3kzl
l6qfSjEEQRmxFksTQL1trDqbs5GuWT8JIDArVBwqg05mG+KylsGh45HV6OXNM74sN4QFOunjA78l
hwvs/OlxlRtSl7lCcB38LadcmMo2jEKvjGmL8ocj/Lm7Y2VNNxwbBKEmn/ealSghDqCPyuVaEOY3
W2IYpLDjZN8QHv4Ko+NBl5l6uYNQ2R6PrSpKhQ5qWS+5L+qRfvyrAIucfUPDFJ3mASaSFDFmrP7z
ZKyMTrRs1lq0TaKJN69Ltg7mq4K+me0bciBE26bx/N9iWCAwp4ucLeDD82wiA+K65ybX7WlW7E/q
LqyMEjw8eh6Ga+p/cWaE69+McFTOEtBzU/0KhMo9sBGS5uRFPyPioCQ2a8r15JYZNNEEF6/Q+qto
+AEUfZgZe6aseVFIChHgXy68hxSRWj0/1+RM9jXiRtSqYmhRKnIUVC7BkACtjcdponfhCfFuirUJ
T4kKPuWGllo5kYfDgWZ2CNIiYdPqWNT3IaeEJsicuNv159OfmEXUIw+HY1rsNvLnu5KHH0rz9Nyd
eNP7KJQO2Cn73UFD+snY1VjhIejQyDX9wtvoYEtNrfh8AkXjSqopmJtHYHnTOZrIX4606GGL6Eli
cfcHqWAs5mi+eJW4rOSfrjkTvv4SJ4chGl/QDZUyPCBzSbO4ZsG2qGcVsLXoqacOYb4M5qtpv5rM
jCX/cfGpOR6ctksQtq7w8Pho2/esiP/CAo/HzAOsFyCMLXjHK3p02aawl5K12w9xFRWf2kerlq2Y
l6ncG2Y9JGJV6/LpSTeKurIAIl9OMLhz2oKNtUHhJPjmSbbLdvLGjCI8oW9oVo1rd6b1qCaKG8pC
XkqmuGH4kEdH/HYRtoz8imFB5741dxit1oDduuTPxTBtSRGSJNzPltV6madhPel4wtU3sf9K/inu
50nJPZWZ+tx8d6Nx675YR3nd5Ned50xeAdjRA+KU515o+EB11eI7Jaft69kMv+HJbbvmbCH9a4Tg
eo+7pLsAWVfgftg510QlUN6LMVVs2/Ryoq8usbfucklUECRbUim7V0+ke2qTM2s+57HIENrJ6k7h
uEtkPtTwprxmAT+yITXAzy8YsmWc94YxiI134YitkBDKDm8/9mfLwbkAFsd9zR8mvs1WhbVLy5A5
XYOSIZaChu10ShlFOK+JBhzUyQLPkZpuBaMHg/aflNq7TDXDxJy4RvTNY9XkTxT5rcied48Q4A9E
rCDR/HQFAR8E+zwuyH2kX0QMiUT7+V3fJodZDG375zwaX+RKZev2HBqewmid5zxvc8eL/TuP4oqc
gksBu1ylzdf9EoQlbAOvH2n6NAmlR2TA2Z8qxRvj/9RjCLBodKlTvMK5i1+oYc7ODri2znAXwVAi
cdzHbWo5Kv6iH72au6HqUTOn2QbAdivKc3VRWiFq3czf068ZupFZ+B4MdF7OpkzDyxcf3jiyDsZQ
DB7XgD4G3XkR7EkybAWHDh/lgR4ingZBvAnaRh9+gTS7hTR47o2R/94yLmrSsM7d0l8H4nkvruWv
6tFaKdNc07ejkIH9kCEran/WB7giu4YFh0bv+OMN9hb1ke5aBl5HXyJ3jPGgVo1iwc6eds/B5P9c
mgNBsU5/3bGL5CV0OmQE1yRuHWqfDRo7tDMV83FgT1LlHzZn6yAyBO/yjQAXQiacOJYbdu2xVRw/
FMkzbNeHyQjerANsKJjEQNLCBLVuSdckWigGNlc2d7g3e63nzP/wbRRsZ9i5CNXiQ6seUdYheJEl
sFwoJw5vkz2KZQZz5YO5ILe722gVzE6BF1kLnkuGk6x3b/BpzhChjOhtFqgjRA6RYZglcE3N/cPO
MIGXBZ0M78zGdJsobLTCdEDeO6PR5tjC2tIOD9skIU/6UpSr07HknuYmNouWomaikxbiC/Rmc4gT
7DAPDhNk6Zprixe/3xnPIh+f8tHEp3a6iS7pupaKQNeMqr9A1vSjLS2btV4eX+IsIK0JG2x1KXLV
Kg8PHtrAiM+0E4C9hR7nfShav5UFWIIS7Ff4aguQlC53Ue2hL8JlLjfJfRJTvHYL8ei0X0Qe/zQM
1DJtNZGCfbgfMzd9TY7Mle5GntpbLwcrCr1BKdkpyQ63XfkaPrsZkEmSXE9KD8HPVPw2Bkc1xxS8
DwWrMApcXX6lZmf1ckZdrVDAplPrO9rRLaLson+ZnmqhKybkT5EANJFql/Z3nqwq8/c7a4koh/jU
hajrQdKEzprjIFAmK/BmnJXxKfUxmphJ7UvR8MQK1r7zt9tWIfUEJLLgorNvEvnNV/c0UOrrLxn3
g4DluQiKVzVSn6ZiPNSRPnhixdpr+5pBImB0ZPl4KrV1FS97FrI8nAsa4rN0Ar9gllOwVpp1oYSp
8xJZlxXln9bpspwwq/27mTsAUapQ0kAZw7wreSDU3lvt2yfqXbQFwqzWPapg9Tvq1fnN8MCMr/fW
3cuac2j5o5GyM/zUGaxW1UU0dl+jGvZ+LBxIPED97kGC8wef6rovJPXCkS6/vNuHNVBtoGRhtXaW
J/aH1QdDtdRn1CCPTp9S4q+WkIs4dIHYglJncnCSOWbKqzzbxHpYX8sNvipt2FJ7OZMH3gsQqO6m
iMIKYBryZgNkizN7Ge+oylvpEyas++KPMaGlTVBVqx8NJld7WDH47hTskrH3iOb+BAK0E2h2/SIa
Fk/IYB+nxbEJjvMP3SvphHrc3hZ4qRPrveNQrnU5iBJBBtGVRCsm01ZMc9qbJLagtTkq5/yc7yw2
rCf2RjjNSv/56WxMwNci/TDldxCuO9wF/r6qt6lPcvrOvpVJB9AgjkEO3ro28HdpUaP2E03NYVPO
MVS2VfGVpOeX3VgqW6SDijWdqmHBk6obQ8AaUcViaPQiEBfnum2t2MfdfDbLss0t/hhjtDg68RHU
aJUH01eb8Q6iNthtx/BxLynOYrPPUUznpKX8LMOPNH+jk/Xn6SaUtffxdSCUfr6P/UC18GRsWz9l
kzJlmel1cN9/iyoy8zrL2OYY/nGAAXtmA3lbfesp1t0VJvEpVnd6YCE+k1DN7kDU811wq8rfA92G
uMJVl0U68DsyvJfo4jvplmq7MqgpyZAjN9OLJlwe6f2iNiv/OkOsTRWqjkqmaXmYZoVDPvbyDSZS
JufoFNpz/QicISs6C57zTJoUn2yq9wLrq46PidN5bfKPtxo6ypQPY68UlpUvKKAGhZo9Fwiuq1ms
qVEPOKtW+0rSH1uOCYUEARGS7wG3S5zA79qhiAbMhkxXuO10wuJiqe3/D7GYRhfx71YyZLF38uGU
n2/kJ8C0nOK7RsvDuu8ElpN6vVlCa8Nth7OMupQbyVXIIk1+FoxlFH+WDj3ir8bNRNSvGEnRK4Tk
JQVC2P2CcKOZ64msG1lE8x+X7kJUQQ5m5p2fKIZz2h3EnJ+6OQKgqbX4Q+KLbdZuGlOuTqvtlXTj
89g/IRatPKj54JIh9YxQr6mdj9sqp9MxC0B7kEl93ynp/9djXuRXT1QQDvW2L0jxLR0Zo/YSUfkf
FCSy5gRrmgWn1qLR3XodHlJlhZQN/004q9ou8OqYr1ydhQw9WCsQTlC0hIkA9vUSwTE/0WyocZN5
iw8Eb5+9WYcr2IQHcFa/oRfboQ7n1a9jP3ryFzXpZM98cdcHH1bhvY89HdMvLKMdeB1brrp1a2JO
XixwkYABbJjVtpyLs4T8g161T6Pd9RFA14B4eTDrtjyT21z/s+Qln+LrXGDLtd/gQSqIockXDKdD
YpViuVyAjZVOcSleaW4kfzFCXiR1cKFeI5HjJY2H5tECQzXh/ioTWxQFlWtdpEzYqw0ovxCFnQ+A
n/jRFyBOI09HpCDdpL9m5nzExlBT2q33wInRqAQptT40TG797/Ngc/Io2C6mIeV13COcpG7ZCE2j
FkJzxvdNWkrDfDKCAxSit9WMZnWkgleg6A5zQ/13d7jB3Io/f57RSuqVqnZ3KikpGliNQ9QZNlql
9usyeevlUt+aTXxIGfHJpPYIwI9vBd/BqgmwqXiWrqDhOE0wpWKCFq/gWHLLHCow+FG4RvWYPKuC
dJ4FGjgK/NSN139uXegZKt7jENM4+GHYjrHO/aKD73et0+TJEAKGvmPeuIJrlhLEN8Z1DNJtfNYG
ZRCLv3Lhc4oWaDBK6jhTMlaLK9TBrX0H2fOkUVdgguTsLfe3DvQiuCjqvN0gtTnZuTU4uOnYFAeM
O4ymT2nEYgEB+VBQVdsNNzzV7wW60B0u91iXhuTxGUVNXA/Bw+sORExVMHivdXguh1/bSqPM7NKe
Yl27XkWRRgd+AnalMPqytk0DQnJor9k/K8BBSWiWY2T2eDx165AmyeWydI2c+C+8F3SLqGAPLjVe
q02sSEq9t+8v5InY8UossZskLXO09/W/uKtEXlic/L8zaxWbQroagxRptWtiAdzRQMan+Ob6zfVq
nVXuZKb2GOxlp7xtZtwpzC3eQ4tG8kpXeUvDw0uGria0C+g4xWXe2v/73Whh9+p80iLIfYB8fQjt
5BtqKyEyB7YciNy28Lzqq0eTOHCYV73PUpaOaz+DrcBw88pWV59PZjf+PEHFnWnkl7+kJy8eRmT5
bsNOMjBK6wgw2N06HRT94zvNQM0/KvQrcoUoz/SeIXpr7ZmOeOqcnJSonUOrKJvPIMQInq10s2uT
hIyP4gsOygn9HGWoB3YtKw1MeGYXYrVM5uftpBgQKHXCcV1Hk/nU8hdDrM4RucvXuiWdiFKcSW38
MUztQ1o+lFGPKxSdbhbDv4sKSSIKtdRnA2GMtJNZvF+abSzQSOCJpdZhLOh+rj0ZQJ8WYqLzvEGF
behNQrxftb4ffosWp4AvJQdXBH7PKhjNruPKKk4Mi/s063Z4zYoUA+AZAnObvVq2LZJsHEkHZqAs
DqkV6dUMNEd76Zf+JYIlhpgDnpMNe9jWWAAcnaELQNK+6Oe2tm6HigFBigVsj7G3CloZ2apdBfim
T4uXxv3oD4hap/CBOVVM1ym3NRPt3OVqRSIXk46J7kaVioMnVA19MFAHqjKeXceouMdJux4nh75g
WxAZfbzCoeuDYXCezp3pO0Je64csTAMzA+VIty/SZS32V+7HKWNrbc54LSG7ya+v6LsK5FIlNomD
r2TAPQp7hiI3vzffQA7kD2e1p8GfL0EB6C2KvdxJU4QY31KAY9KV/3HhzmmWHwbMkWNefL0QVbf4
Z42MLNFPxbIafEy+asHe2PMLeaSkepzCW5P/qDPCIv+WmQQy4rKK2HrnWShk6fpi3zNm7Djz1t8I
WZkyol6mDDcAK6cDdbK2i5X++rBx2dsTlqfei3p4v7/Dc21nKG+y50bcIClYs6D4E/PUynzjE+XT
VNnbqyRUrX6y4mB0DajxLk+DLjyEfKilW4A4dX+3xjPZ5vAKLkotfWcGYNB0uEqi7Vp+QGuBhaJD
rFM6HdxqpQqj/eBD2f3lLU9Uy7e80lT36+7rMKF0AJS3ouyLvNWOJILw4koy0JjueHKWmVlF/Fgq
pYjxVjVz6pc157/8tzyVYTvqDq5szrsAvqeTF610vy1fkw19bezekUouROw7JYYVDA9YJIANF8pf
n/SwwQyRavbU9jhtUoAdytQdSE0oiehFEqrOIJB1v89EfATZloTSXmGhuiPGMXkUGUO7BpaRZywd
d05B16wHm2wQAQtRh9Yk9FvH9DsZiS1MF+tg6rg3agqbptyf/oUEdJedM0kHxou1OoBLuQAcI9ov
BXDp7+t1MwtVpaS+3/0qHFax450Pn8yNUmUob76GmyPvu4bLFBqmw6PgREUfrDTPjC9pJqBSXltY
MKw6hNYE+I+klUUEsCsdN3q32lGENmAEei5K2W6nH2BxP4psT3vvaCSe7aJimBh/DD1DP0dQuVBK
aXjAueNtAILpjtOzEU0MhXcrCxpI8/g6dA9iYG8jiY38cw0VL28pHNMegc73l6xpKYGReZ8vV0QI
hhO/F5/m7QqD6NtymFfpkxtpb2TkAQguK8NmyuvdNEjeL4NspG/17JdODK79KXEBqJDDHNpWBlcr
LPcUiF03jgKkNxbqkjJESlWshbBwpUczSopmGBPVAnzwXmHSgtKgULbmAnRDuX6dC4IKiMmimCN2
5dBiP26KlABhSTzU0txs92wEQkw06wYbXvawwGqZ9WlJyAfDXbd/4blD3JvwFeVmGnHrDhAx0q78
3Nyp7xsy7z+LQ6PareQ4//ksYLZRbaceeY86fO/DGBsfv+73LuJkOxiVZA213gixz3pFT3M+gidF
WZGLSZYskgyXmWtjgyaa9yEeaT9fpipr/Atb6oeHFZUbe2aoSP47wL7Tmqc/64oB+KcduvRMpzU5
ukjtdyCnvxzqNeu7UycFU5pDnMrjWQgmhm/3uHOPqtK/iwE/xntkDEJNB9Elk6eNhbuRFg6NlKUl
JuRljvmhE+QywgHRjQJOWj8T+Vh/LWbg1ZO3cJ2ey5HMnxZZlUK75aJzNN61OQ4CLinfVFbLzdvF
KYUeaSOB95QPPwMeaXsgjFCiHFcS8Dh97s2oWGcXkYUzgWz9xsRGEDhRJFLkzd3f6NpCQmlhuRZd
8N2fuqtyKyNe6WXp2XfXA8JS2qA+ffhQUhF1D2ClJXxp5j/KlaQjxZqIlVb1NaiJL/IYnzz4AVpy
EvOG0lgZ3N+tRxmbnbvkOGFXT4WqH/AfXxrOsaxSTjabjhvmTB5qhEHREJCDbbigzQiC1gyRXTcN
jkXoNhcgdanmq4SYjtebBayu+qSS+/Zh7Pr7UHA0SIgFwF5wdz5o2HQgphE9xx1hBVs25ORFY1C+
GjEjsoa+2yT1huzvDAuBjXwLyvGCxcLMCnJFvRTrSdaUPCnX0Zx4zh6IReOTUsfg1/vLqNQ0Pk3S
GjyuU8hQ4mLaRsBqVaY21UES0tUafWh028A4Tre2EuTH1kMR1O8sWoQMf4bEPaUZgxb1+xlsD3Du
svidUt6oavoaDG0WwIlIG4yYxpEkuzk7wzmQmTZ/0BIIWuAk5uG4FZFBxzhXYgFgVqIcQ1kAnUPc
vl0ANEhR7Ie/mNAGbOw/WHspzi08iotMdPqVcQHebjBhgBfP6+M3+uuyKG4MONqPjFm9ypil0Qej
mF+LrGJ2WqQdagP05LCYugYSdMT/MyqT+xfLaNY1TF7iJPWU6+p2icKCiFCk+OKMEzGykGm2njQF
mhtHhNjxMTohbhsKE9Q0kSk+CsqZUIjnu8mhJOLWsEEvoPSGNraFQCYcVJOCFBfSI2T4R1xAmRkO
yzjRIY0Bq3U93aNFgedr2C6XLIPFXJJFnnMOd1CM9zgPeYghlDNuWStxNVn0msOybrMNhrvN24i9
bAK9npTryemCxRO4tqsUuIdESHF351oiChFBggXVFtKfFAu1akJmPZwZDF6ghFEsY7wN3hokxqY6
2wnWTYLKoOJo0zRPOVs/zB+JDGSFYSg2qoEGsAmv7ZHPm2bKrmK71Mr90voNEpg/MCgjDj7AN3es
4VH337hOEE0pGp1QVDFfOBZv0lzZ5ZOnyOIase1DK0t2lNTTOgGuIhffx3GrBqW3sxAr5yFW7HuJ
Llp+DAbMzLVwoKppvAzXC3CerJL4PQaC4ruEqQW52MwNAsubuLtWaOb92zTF2s62EYf1OVj+XFDl
ZBLCV19bX/agCr0JL4vvJRB8Pm3jxstzSXAOvQL4OhJJ+wUn2z+AE/AZBRsz9S8pJxmG4MdQN3Vk
o7qtgirOLlExMtMO7E5El30L3DL3uW1U8j999SgA8ruDMq9tDgLpUzWoL8pSFPo4lJmPQtscK+H1
NvlzNS+cnXiD+C1VB+/MRktHIkgzIoH3UnElMxIEfJrcs86oMO2WW7SpqwTmmytXK4/8OuZa0XKH
UyUhSPF7TO+GJneTM49q9vcydKdWqEcr4qOyQ3zgeZXuckfgbxEWzLdY1UgmXIvzuWqsqWh29Uio
72/T4rTQqpWqnCdGC8NNwM05+t8l66Nx2s1xBh0ob+ZjWzYCBr3StVtSMx9nO7lzaUPy6u2ro5M9
kKSYZJqxTLPPR/2L2PGMwDYB44+aky47wAywpg+RZWONLr2W8cOcEQPWepDuKktoSqdghYhehOVC
7TzmlcKax2njHui9BBb5swlGmp9RxDjhF/cCcdJqtJ4xMdGR2aK+hzuos5ofKfJ0IInDcLoT2OFy
dwH6CsdctH6ZqbYME3KPFVE3kYdtpuSfsNSd36UzasRDJCKhUEFkjnEdNzkSGsqtfQcZpbzCm2BD
44N+yy1Uwq1hkTycHrM0sOhrO9eyxP2zlNJDbenzswqTsW+dzm9aVvBW/oW8oB6hg+rnW2vboMhe
/Wene8muvzXxlJ8cMz9declOWPKC/fUsGjy4BYw9CfbM8xfvzxsN8ziIOBCbcgZmarqaIU64AEme
F2Edbaou6pzTk4KgzJ8xTLL9bbi+GzFpUxk0VgcsvGM2m5CPu3ZcTqHmgqCrxi1dWV38QFG8H8s8
5lpAN1eWYsOQ/yxVgFHsXwBJZbjIICCJYOLJNRGwo4l+fDs85C68maRHwwrV4AnybdQqbYDjsGKP
yn7SSEUOCdozUFxO2kbLPsZoYxsllc5mRXEkOf188w0/jNnN63EtAcDpzhG6DhPS26byUwW7rfRq
kjIPOAwAt41ewbvRfMogLBh0EPoKY+b8b9ujhZGOdTLFoB5tk2G/5NgYs9onbzhb/vSwMYqDInLI
Nu/i7hBvAOEo95pMvceCSHlVLfzLOYtncI3wI2uO138YPpF8i3dqNsjkpZVQop1WhUh+C5dpx6Pp
0ZL5T9wliIsmdz0cXIcumus5DJu4hXgPkYm0yUdm5ASM5ypZy+hEPd6g7cczyQmDxgFUthM1HdS5
4LiKRxaveZZQoCOf0tOFTTgswvQeZ/ShXPWruheRwkauftv3Qx+zqPNVkKPgO+fRY4F4fXodE7+g
1rg8nZuOqT47nAVHVTKqJFLxP9HwTB9xc+zfjUeNrQnSNTGN0h1D2CqIx82REGnpex18oN82yuGx
vFnvT5ppvhO1LB2grhzTfNAEFZvEyvyFqB1kp6T8sC1vENH9jowCtTk+ORkgkabCH2T0VOPmir/z
yn7OSFqh4zQlYjt8s9wh5KxPHw7t2UnwuoB0BoijSMJvceU8wpyEl3szTxRqnn+wenLoTWPs7nPj
2sFCiawQWm28nVuYZIBxMN6e/98h17+5nsxm+Y1FuJ/s5jrIjAMZHshGbbOpvtH8fVjwiChG77Hx
j/JAusgqwpCy7G4HOStNHPZGzAIIULcGGT+HzDyUOmtbN+xIXg08GrGsc+pvSDZBk7gtSiZK88uc
1m7YXBBZAPs+KaYa7dbWasSboGshe9YTgi3ZBulP+BBUZXEi10KY8+IhRVfXLWtTo7dRtd6CItJt
8RzLPEoeKh7VWjQvlk1qRTXX8ZCsTV4eCEDYJr8HLaLlpmiusP3lxcKv84zaPJUieLt4wVhSSMTQ
A83iGeeBbKF9dnuwWXzHMbw7HxWveKt63mYK/RBjnFRDnb65MeQjwzLPGIUIYH3V6uUPxmXGQyOX
71ZYWg8frPaIl0lVgSwncuz9rh2VaQiGQnh5K6CkVlEXPmD9BbFB/zY3B7tfmJavVHWAt3R2qV1N
y0iPOdlpGpbStWoKgtjLPFlB4wsCmyI48rOUxNAMKmkL/GEYbQ4OLHpA3K3HtQsuDfhSxcuKFg09
l8cliOMpJAcdn0uI5LnjqjAhZjPvkw8SzjiYdM6dbdoqHTfl3g/xLgBNmd/z4B3mP05fcJbctTAq
yG7YH2lOvhhKl6RPgqsN5skCukKtW6nS9yaXl1/jcH8hxAhL09xLGbvGd6GHb+dDhpxeCXvFQuS8
UJ/2lbRqYZD5HRc248GcionTzztkr3+VLzJa6fPQF7yUA20femZMieSfooxHd/5A/l8FxSDNj/3b
oLvZzGYcy/nV4zrRVFaDy3L4jhArY2Cxt0ht8I8SbaLaKICW+hXOCd6BRA/vp8m9s5lFbiTGmJYK
qc8sI0C4DYWOZikhWxMaPO6lGbSiAIcbp5hpkKurxAjLeQ1pu03lipKmkZAA5+yG4WFEFHANOw1B
6S8fbKVP7wdeBAo1xK9eTYBtgc0CmlPmUIb6MqUvKrDqjQ6hSsrC0yUDPbXe4+d+vk3Wh0cWmVYf
FmJQK0GpaZmBSYdz3puJFlNzvBlRYpVTwSy712HErklPXLE5VZeyjuGwNb00stjbehlbsGrwpO14
N4R3XS3BLAHehOHOxVhUQ0dKba5vz4oW/gnnhewuOyxL7EvXhSd07X7Yd8gLgqZrcPl1X/tFKpad
lgJf0ThYLLW1cA3K+hCcJvOmEJ/wjoHxV8mxESnuQ8F02xcoC3bzGGlLcW8gjxfvMYbzl9Dh/H43
8xs6sISMBu0LWPEahmKN7pa4XijL3FYv+u/e0If5rLcVaY+b9d8PdW/whxVznqlg2cIci+KL9gSe
4gdcnvel+bPGpuXTWBGBnUpL/pneIqDWu4paYKwkIsdLXh2m37C3REVU+ekw6mahkSmznx7Oc/f1
g17CKwAnjpjLb9t1lc47OevGKz1loUp7vkvWRoeqe5ohmY8+/WTvXCkZHWvnZ+b5gIgurX55Yybf
+G0yoLuU0WcXnenvgTonZGfyrjAoF90wuNDrIgGYTS0AunokDDktZG0g5pFjI7xxjMiM4CLpmmHo
to9QLY8S5cEM3gjsJgSGHf4J8ZjzUA97hroeOeIZOFiXJaIp1dUBiMu72+RxSqrXqF8OxlQ8UEtZ
cPTKawrFRiquRSJFt0YKxcZ+rLZNBjrs+Ub/74YB/XaP88qDAQ4w6RuclnKeJIwGoSofmRZQalR7
EmNefXve5Mq/nhb9TWcScYpF++mOIEfx0sOF8EYsZJQYqPTso9K42FzGCstqpmkvq7QuFfl0otDS
YTHF5rlSbUPgM2VIrSDez68P+6NZbwZRo7T1GGBqsB/siDC92zlWnm1jDw5UfHZFMvEn+i+C6aXR
V+IxmxODCcT8hWWBbDB+T4eBEBXENmyQ5X5KZa4sFs9dg+CJ4YrdbwmlgyHEs8eGryaDXmQZtBT1
Wzj9r6KDbuOI4i61TMKaj2xIwfW1Y95Fmf+RPw5uhgiphkRkv+DlIjrExgcwLXt4psB5oXaRZtas
XhgPlu2NKwG81E6+N0jzhv4DSnqaM9TrEmj0RdiyhRaxq/S5EuZazHgNB+KDXNvhDX4Kqs2v2VjV
x0jx9hJVQXkoQPXqAczXgwjyC8gbT7f7xq3HUlAtQ8GwDP+8ylj1SluOmSrzCJqqAEL526piowRa
yJ36sRpAOM1gxV9hhSHBNssiq0UUe3n1RY01W2i4h8tcxeXtFjj6p8m7Zgp+3U86MA9rn6NqTuwZ
Qi1PNibXvbt4qk1t4vsWyGitWbOyS0RLN82bAC2SjfJZ/d/4OB2xI235dEs0qBqjDYpb5Zrc642Y
c/toVZZQQzOaz91Ru5Gj+vyvKnS7+xmqpshI12m87VVyKk3NflnhNND/AKX2TQnSs15c3QwoJNVQ
Wj/v3AQpWPFPyBu8+P8TKyXxHeJwfpu7y8VRbJcdW9wLqNFBAaxqGOrG4i02kjI92+BC+eBxgXcO
xzrTDYzRVAo36u3uKdF661rofKEOBHgmImFNBi1/HGWYzGeTm630hedEupJlCccqZIp+mCcmMb71
Iyj/uXN2to7sk4o467bRxa+e8ALe35jVkRJCejXy1iOsNlA3K8PnftMIFK2VIhZpR2DmKNg+y9yo
3zvcgksxWBy38dkA235hHBLJnIN+UXdlz8MkxhVhLGGvCqugNLUM3kXgY0VBnH/p1e/DQjY5EF/P
wL89syvGUkzleRHRPhBEtEqACAz/kYbXitInZDcrcRukQAUoSOOlCWKSDCai+08HvrCGCJacQN52
yX9hO6Koim1Q6K2AExLAv/YnGwDi0OS2kgc478W8blDEtTDjHT0sb41vWvu7NkG/6IdKhlYxUBQz
b5AFtHNB18G4dkrUQdmjbB5AX5dYPybFseMO1GFudjM0SzaQhFNgejLUPHLboxyhtCX8KKyrMhy2
k57/yo5qmSqQ4XTDTzmf0rgM8lf6K+fxjwz5NeDWAa9sdw5Q70YDzmJPHJ0+C61RHsx8dbZxx38Q
grUMFZBkmTftDoif8+EHdpJZwH9ontKBlOXJ4zPVWmJYhntMP03S+y6BzX8nXSnFJ5Qe3GcG+ND9
Mr10llAD5Lq4OmI97i9G00+pvT7TVhE0WzTWMH2FMzxdlPbzOl2wQaVZ0IbzHOYzfIlrl4OgvqTd
ofTITO3KZ27y6oi8aJreUMc8H06V50KoTDW/BPFPvNhzE6byxOv6ftJt4jHPiS2xmElJUGVwl0XG
DdvuPRoTouKPpekpH7RP4zaQFQ4GaOgHrwr00PgJd+uEq0BGgOpewV32MmIK17tuiOvBsTJmXWuB
nH+0zkU/ld8BB7oDfE1KW9q6TjZvRstljUEI/ytNhXRlPSptheI83+HRr0dUk3buY2OiBVxp0Jud
ZT0e7osCMVWcepfgLmyQqCqCrF9uox6f8HSYrwqeiyzdyjgJDdLSfmiAu2WmoXW7WY+p8fihBOpx
7ObuWBG0o9uXAn+HSgKVAA739yhDdFPF9fGnO37aEuH3O2m3KHKZMVc2lqBOQ1LQkq/ODtJFVZn9
JhqKOVpt0GyHOj90bD6CXOVrOYUhqAXdHhT3laloXexGg8o+k0zTttRPgtcsnJGnRT77RaUcjSpv
nLliMqMrJglMxLqHHxImN/bdlbsqRsoJMjqmh1wSOOBwtRieU//p36hFBaS9KI4uxN4u/QB9g9z8
sRNGESooIB7Ioqx9SW0HhY8kQFP55edp9jqg6gEivwX1Nb2kBxeY7T55UX2LwFpplL9KqgQGcCBw
p1/8AjWIlXgVeBfMLr8zYs/iZUR+UhudhA/14J5bEs0Hpc7CGEb+/6mDypELqNicNOQKODiJvt+F
KdYqzVx6taY3URwSMatfgIg8vxWjoTYqfrn241kcpJ1tuUeUZtSpMRUTFIzOWrELQdcovzVAHMRH
t+F7a9e1lJTj/rGa0zBPEct+zz9iX9scI+0SZhgTwLc1TTuVIfj+rBNMBRPEjmtf/rQIhMfIviRt
+KyA4A1G2f10p7KsjD3pIiKRZauftXIU/alKlj7WfZ00lIK8Wh+EgyQn/alfTjiriD3DdtZLPSc2
c+EMBQ2qj+ftICpOOEsZS1vcFAEv/qqALxRL6cQc2Sw3zCKOLQpsOb6TDxK4NpdIA9/swYk8greE
Aap+/XKBBp4wgGXtlEpOpa8KAG3y3gBZPVMhGJIyVyJlakPIvV+HystxCyN9sF/uXRWAuLUJjeGa
jCdEJFKWLScFs29TuEs+jNKumk09OV70fxX2AJ2OuhqWcyn3iMcmyGzt4Sqb1pqKoPdsKCI6zIph
z9QHsh9433nXlYDDwplOCPdYF9njZCDVxYDperdwqgxsamdWidCp5W4eKFrY2RdEmUSKd+JetKt/
6KjY80qOoI2Lz1hLzppSNCy0ELHmDCSFz0wqqih1utl7HMNJMG5PY8f75kzZmIl9vbvEs8lw6ORX
34IL+aqmG15Ldk75KZYw0u+vAS2IM39hi2Mi59KLHyXpB6Qmbasrpivolj8/V19eC8OSgy9u7oAr
0iz//PT75Wt8Ymem9KjHSV7KEiw9I1mgKCLmPWPIta2xFqdqvTlJTH59EpVQJLlTRlyOKikocKpQ
hI8lGlemJeV9bikliZuzX46TqqIzcpkFVr0Y0CxJcWGmfobE3n1Zlfds0G72RcYIMNTIs9wK3RK/
HaZK8+3hWy6yZL1BksAu80SijiEJJE8skex3mTuVbCsnR3G/aeEHzHZlBKyMW4TYQIoRTxTc2bGO
YcY8aiSRAs4yDh7kERD9+VmOU/O/4HWGzHiTfWH6sLNbTBIJSlPaABCwYxOsjFLDtIlDtkKHJbi9
UPpMXwu9meCzjUNWJrnq3rX3qK2wBHZmd4BgA6HghrhVgmCnB4j5NgSHWT8TuGvon/s7nKrUeaNh
ng3Iv3AzIna1HMjc4fciBa2vuZx5qk+Jn5oxs/B7I/5vrJma6syp0ZRHv5XNHWUpJRjFiFEyG8h7
4as94cN8pr5ShAEvkUYM1u6njqCzJXXkA0RdPCyKc/qoXvw4F0vNmTfhfYmt5BaGGDmfBYszF6QJ
mRnoO8t5LAjyscU8uKPmhLgm9/+SCLowld2emdKmGPvTVuqAhGs64wzTQIMOQ6w2HfRyXh4DN2Qr
//KTJyBo1dWjgT2EDKxZzRQ+4AvRpRbCxh8yP3aXYIKrCZaVZj5IynSfJs8LwSYClbO8FLn6Zrrw
fzSNZG///uipy7AW8Hq3RZnnAfdbcllKXMQqw/tbykk9BdbuNlF6qWMnHoODSl4ifGgx4doD6oNK
y2YfgxogIsqdsq/ONGPpbj4QLde4rhEGYIhBK9NDd+wEjFspUxqNvkqIYPIuuG/1FVBa2csOuaqC
XtBT+hwaGAoyZc2tFC0SKcP018i3YPw7VunmmuSBlY+jskfnEk5C7lAQE7kdpXd0HcrHgiic7S4V
Gm/UWb3PAzKDnBm+6OCO48Z9gfGSIUldzPSG9s39PLfdqufN6O1MPzyslj0KgkFIQgGbz1NjSQdN
1OBafXM3WeMCYeTi2QTdK6jUhC2wPfLgdklCoIIhb/gHiD/lMOEkguYXtYjbEuSF3hVS9P/TocQQ
tO6tvoiKsRm5zwnas5+6GiN946NNkGIronceDCoNsyeOFOXX6nbmvD4LBRCQtc28xVUg7y44bwcb
FwZxR0LMn6mCz1kF5V6MIuRCqBUZ99B34NECzx/UWWXucREPesn/giIOl1Ed32vHVEXIaiS0W/zK
IUg1m0IF9tnjsGMEUALimdnXMHGcGQV66pecoeMrkoJ1rxJd78gIncCRrWHUEHa7H5nTYXc9xu31
UIp1PgVkP9RNsfUN1JSdgJ+VJZ0HcIq3Z4S1ZqX49aJC0zexpuO8Ka5f83SS7QhqUZmefA/xjbWW
1i6kBFZ0pBKUz3gmq8DeVTP6o9io8U++Js+UgQAMkIqLG8r3SXdQq4Bf3yFrL9qArVR3ncxt6/Z3
OQWTOzeXOG1pFgaKkM3wMVDxVQaJ02Hz/3xIUJ3CXH1JMcQUFRfejASdeEy0nnYluXpXrxn0urzf
V895b3sbOHnYTjS/sotvKWJeY8Y8axk9Y/S/IxHfpo7+Wiycb5M2hNVKE3LwY/1cA0Z3sP0ibRGP
wS8JytJd6YKn573BwLlEvRSRoj5SI5PtRoVRW568RuVyCP03hMELK1nljWR7hQYLiIAnxIXKvXXR
rRUku3zBDazcP4aEepUT12MznA2/2g4LGgvtI0OhsW2awEBDfRhyt9orjQ/u2u3HT2B9hc+pYhB8
F1K99EJ5VdCOoHow6ldRIPEjcIdEp4zzp/CgUbg4s0Hg13WW0AhIwWy3G4zLleNHaxQVqKa1IoCE
RH2f9xXkYNUJrQrLV8+s8d6lRLcmfCI7kPT1MXSRswg/oTcZ4iIRaTIsmFSFXojcsmXEelRZ4QYN
rjjr5P2I1u/rivCpHzG4pOAxFvEuq25FAec5O6VznpNfJ0vPWiApOtTfKflDLavaVLJsD712BNRN
WGVOFdppmPWjFcsR0NF2hjT+vKB/bXqhncPHi2kwjAceq7etFkT/nCM9QEEgVnRNJoSxUNPvVc/v
pSctcVWQK+scKsxIuBMVrpFwfrMiCm563n+aiphvHDb4lEgFC/3vFzMFh26fbikht5f6jVZbQAjg
c8XWdOyDGbv/9ylQRHPmEhqUokH+Gdv96ldcxHDCse/QMCd/Pq5R9aw7yk8YChzaEiIRdu+AjcpO
xJjEyQasVAreXP9pqQp6m3IyD6HwFGjUuDKRiA98x/q76/wt6zWTDlxe30Ynx9Ux6fkJJKgs6ULd
tRbTeOX6i1sAK9bOGaNMgmaGTutwIEyy6Hf/FKqUH4HyFrImAGvi0hoWUm2OlTXTUpqcv+ahaK1m
5Rolm7gHyHPTVDcnMjOWElKCcgfy0tKib78945gCPF4awQU9W7U5AHV0lmbWmX6dRIqIy6r0tTIl
6OV4LTf87ub2h30WOXGzDgGpMh4srIG2+06aKa0ofJV7E8vQl8WU1W6DLbvsgPKidJvkSuB/64+c
V1gpiTrjpL2hBuahjGz6PuksCE8qsh8reQPAecIeSe3DmTmFxEBKuXfe567b1LBIZ2l+BxogyFbf
1/nmXeX9P6VWCXrnGXVV6NrZGcCstL0De2BWA/87rTVJEN6HRqeYs5FRfqx9Cx2EqRPG5yJEDVec
NU2GXr3Q/EBZgE3olXRaMu9lkAS1a+ahxzpo9ojbG75IfvElFBt+QCjQIdOdqcTZ3F0WLlHJ+q4z
1MnGAnVCuXrUFwAS2Xy3ix4CNSZkJewt0w2aKzNcIITQi2GPliyS9IQB+0c/p8w50zbmEoF0k17v
68iFypi+yx+P72E91Og4OEu8CNpAgZVgv2fRT4DhMkHyjloZb044rAho7YOKCGmPB6PwVgD9eVgd
9wI8We5XbGUyjotzqHitwwnFMbgK8mnaj3u+d1EqGtb+Ivj3rFE1soL5NO47BmBrXGEPTMMpX4oA
nsPP1SpQgV3+N4y7inmq8VAMhAc3nSv+NnKrf5T4M6Ag9D4g4xUYvm3JI10ezN7vMEWU/2EHHs5l
GAg4/wECO5Ka7HObpwa2B+BDqwrzmB7/Jz85Pofyo+nYviVs4SSx4t2Sxs4TqStrttFdOCj6YYCe
X4x0Wtu2WXjUy/kTJ62POqId2PiDsAxC4rlrPNKcZ9gbW+44Bar+hqzsFRB7ewyQS+ve8fA84JEE
38/q77U88ZJ9z8kQAV3Skf7oBaowrxLqNkV+qt3EC0MqvRMv0yLp5l05dSWiiqvUHGFLfQPLum+Q
X6MVkHA+ai4DJrsciTB9ak3dvkU7R0iBFkbbEiURhNDx0yng0CbsEFdTS3vIbNBiOOn8gkMpjF3S
YFALhzNHXnzhJgcKiMuvb1M/N1b+adA7KnXaCitE4D9nEyJfFoXZ1LzIT/3Ane4b1MYvqyGb7m1U
cmvMUZi6RFLiiOS7XZ9u2raDOWqVST7sniL2qhHLFznjbb6HJk/UaZrOAN1y9VCRYaFs5c29G+JC
5kOYKFK/pRLHZJiySbCAdcX4KEqneWbd386ZLhJf75tw1Eg8TwabbHjtySOAzBGhpEUuA1gbwtYG
x5e2pOQo6+e9LvlEU8zlbkI3BJSl80Hr7IpzTGHMw+WDLtasGKxxh76Lrhbf2H13rp9fsr9Jr1nc
9JosC8veE5iA7vVUWIUALdtJUuBsL/0on0cFBSdM8q+NriPJQ6k6fNFGd5CZPGME2j13yg/dgKcE
n09T0f7lV9su76WVZ4+9AqZhnNz1o7qJ4+itKnFNrP3c7peTpjdAfln+1e5xdaRe4JwhLix4yt2D
NNiO7c8PvHbduzbCAXxJXujdK7Pq/G9UDgOXsZt+Juq8RwmLulVZ6/IqWmaUJn0rerDxvtNyOePI
2XlNl0fxGeG3kfcitU7YX5E2JL7WCft2J4PSQCyNujMynJlF8/22eMuIir3SkW+k2dGweIiHK3O8
BAda8GBBZcEuGQAug7o832sshZA96Yw8tsJPqJdMO1sfz/inpO8gkq8DUtKchfL5gywRk+zMSBvx
3oudMjybgX8mN85OA2ppIWdRCnFpIK6j+USoGumlsYfyF+R3sry1yUqZNGXasu1NZ3YupX4IA1GV
TBHE5aLcqsqeoMuAiuoO+b1NsVZTGQZO7bTbruHOsFZ9BQ2irMN+w33xxm9W7MW3CiMrRc2sY8gM
y00+f1UiCiT+M2i1cZq5UPrcIcwSENNHnvXxgZaZ8SZ9rZid6Z3wTTjypu3bHoDMqNYsrw/nP83z
oPnL0W9fx4pvOWayQ96KCa+MijZZ17HFqe1dUXkKzWaqGMmE0etXOY0JkN+YCu98jqr6uoLir1Td
j1Vs/PT3Zy7FmZEUzx2Spz3XS/+2eKpm6++EGhWr37pMduxIc/CP19jujHTRFu/ADBr0+M5Nt+Le
0rAjcfFb66a5RoQ/3fLfbqR+ybU3wNhGALqWL8IVX65a4T5HHRHvc6+nVzSLDKx29u8ObRN6K9Pj
PtyGk1PTt7hAE0n0D3E60BKh04UsWhIBYYpRNfkWxaCiKYk5VTLuKBJDUxpb24HZGqYlWzkftSXD
K5g9dg3tfEPkYMCPd3mto+nRQYgIC9/Ywqrw1zT/26YDXAcbI8TXLvrGkVjM9R0/p/QXJiel9uoU
7k8c0fBe27SYrHTq/9cGA3vEH26f4McmkovGlk67DHV0gejw42rQd9Nzehc9qDkq4+1AoheDawrL
YPYuv7DmAxQHkjDtO4qsmP85/wOwahF4XjoLlDQfZ7mk8oJEo3SzziRQKJDZWeOFbyluD2X/OXi4
68ys+Sbi0f56Oabl0JDqzddVUyomGBaWgGPiyGaqTln07rnfS2+Zlw5jXNgtpz0rJ73JtOy0ngcR
pnRPJ91bKbmDg7zolFB4D3sGIhbBn1pxiYe7vcs5WhyG+RAGb+7PlIuUqIyYTwQ6VGkDA68KTok+
Tvm9Rbh4+PQwZmRJ0KReNCUwIKJTkz2tnQUBzQ4WtdQUn6P5GNNc02ArgFk+Jl+v+W1wlIcMJF6F
s4/NGG+ACwKcw0opZ6J+KtGQLKRaWyRtKEH6soR/VqyVYkEB8qGrwJ+LSqotJaNoUdsbzZdmX4LG
Nk9EYRLvd4ejaDcyF0TxSZTa7kFRxAcs+D9QXzgzPjP0RoDdUDqN5Db9JpcEhg0GlSmKNbXi4oOT
QEd8eGeLWnOV9A6jVIT1CAdyVGCLNHHze2qv0sMLB8QoTYzlvJbFSY21H0uBfDrQYQ5G7N2QCjNa
NFauLKQxk8d5JNCoUlhiRNK+UEEgpAEyjBmIjFFi5pdb8ARv+HCit3epbij8+f28bM09yvrwE/Nh
A2g8uCoK3eT0IuTQRD7ImekYSGQICbEHzuaWiPRMvsyyPrhDRqx0eByeci1KY7HEVyCgXaG+0nI7
rE0FTz8d3Nt+8vprFf5vZmS2/r9ECLojREx0ksK13oyZkHTgqa5kVc6czwGHEwVml5t8H6HLtWV0
lEvzkwBsh8S7OqM4ERRuI23+CpDQ3XTn5Qmy8CGwDG+zukfr4TwqHEoLCvz379LBpbaA6iGwBDuG
3x4wCVcuVq9ymi7qoAeP/gHAfwzdGwBvJuXOQNLCEp98hOO4gPkrsCLrbrxvZAgzqZuc6q1nx60V
8XxAwPpB3dTxQzskK1LXFyxwE9Fe4t1nDpwI38Q4LRxVW4so+FTHg/yA58QuX/SA4GtaXigZlE/I
btrOBkjc7ahC3yWt5mXOpZ65r9i31jFSK2iPkNAUuUp+JgPKteNrFPwLbBLVVUnRqXbOBQPRR4q1
7Vc3t8kDLPwb0c6uabPWSdfXPfMVqwRqE9j2Qg7s634w7B1YLvTUPoZeDL13C1P94Gtp1Cp5Y6zd
VmbNytLDEEj2ux+NO51sEMcq1osZQkELoRzDjYyyvbCoTvSORJPhra5eTE24dmDyyGzNTCSM/Cml
r5dOqDP/mhv4rxayYaqIardzwNC2I59jZskXsARmSGzETWpU18UI6a9/nFpgqNYI+OVlrqm1gtbM
h5uG+S446ArNnZ/tl0vhgs/RjSdni5DnSeZLm8iESE2lAvNtUvEPlk4bdT3mPnevM7Yxqn/mHrVQ
1Gxw9FvISJCx3Ky1v1bfIom9EtwgZTbkIKdBSthC6+2u1H3gN2kxWm1boSPtzAFtUqGpYOGGlmX5
Jk8LZ0P0SnTub6GqKtIDMdtieitFOUpDXUqwJZShYARtqzuDP69IIkcTjb9uau3u3MSPralgJFNw
5eC/smJqgpB82QAOA8IVt7DN1GLVSCIBPkqXKVPnWobmtm49zGr7Qt4m8cUwFKJos+TNt1CxtAeA
qRpvpPH44KM6ypZL9Vpu6uRldxHmtTW5TKhBj7V7fPQc03xKtL1mL50mxgRQa/kD0H3gGRcxIASv
CY9GvMv5a4FUTSVcJh7XQ1LAXcYxzzkJ2IsjlgfEPIdX/okxYyX4qvI4yzBrvHOx4OiqwHKdvzrE
WEk0KLSieGQX/qhF4+aeY767Cx+Y62mS7VwO4u+1PWwEB0AG6oJv2ByL50Va6cKEfz/fxNuyKIiM
HRxcoZ45exokMKVI1Pjhp7J6hufL+C2oeE31vnxQvPkbU2CusLmSpMxMZFnAGECCRrPdjNcq3LYy
DGuFC5exv+XOjdSsyh0GptZ8Zc7u2fTtc+zQqmUng6VEAV0ngWu1mqjvOIxphcnkj+ssf+goYq3I
tx1M3WpYVMoyrq1YrKKy7CYpea6gObehXzMkCvbSlE75WYU5LgAyN2TI9m3hvbW4vm3hbqLHMiji
tb+emv2dkd2x4+pFEfigI+ATpBCS/00RTkSXwtIQu3nEjV7EdF4q213otBhwdVS0Ylt77nOfJ377
Dg28hMbw/nkUi1fTVEcOx44jdRkPxMtwuWlLdPTBMaIpW7mo5lJlGNBNPZMg8RXevFBNcIskBa8z
xYswu3RVt2CsU5+OLNSb43iuO253aTR2pqYh1FxF7k9/3JjLR71gtKB0me1xRS3lML/zHymUCEKK
aA1vJyrfPkmNrNG6DdrJ2HKdqebJjLuQvXOs9JL/LOpWQv+Sc3tsHJx3cTZ4j2+I1VrwCKc5yba5
/LbkMwrODKc3Y3aSjZXLitcY3YOjD15RDLt8c6+iFFjt3+GPsCJD6NAqt0nZg0OeeIhy/exBJRVI
dGdRtBHaal7GInKmoCbCXg0WojBZXv/m0PIpA4un1aDw0X+2BHE2Fdd9gAtiL4mQwo843W8AxxVz
cFvpbZBvtJAagVUCBWev77NvE/IyzW+V8M5I3DC5jbQmVNLOOo3602wtnyJXTPylRhFMBi1Q6h95
sHOQexaBEdzELSHuE4zXW6mYb3GyVKUYwGITsiBhlh+vrcCDaM7t8j8xpVGN2WyOFY2Y5MaDFFPH
ZfbaCu7Kt7L7nymWMvWN1s5RKC5qVeTIxJtVGQkXROHZYi2I9hqkNH/cZaGFN6MDndtXnlv/LM9d
kfS2F4rqQJ96gqnke+oZyO/RHHD1OzjA03pmvdRHU/75+rCJ97yqqsR3/Low/3BspK5rIwDl8SLt
CyyNmKhe6viAfNPZOOL8UNLbDoUb1+rp4Z2X/mJPh3aLcpmtPwAwswIIEKYHdZ/b9PX/vZZ8pA/h
GqP6Nnh8XeyvZ5vCwpXjfE0ofgN/1jkJbaSOt/H9790AVIEaPP8GxDd2hPjm3kP+Ngf6E/AIMHLU
WNBRuvFvsL58uhnqnYnU+QlGrkDV/dDaJpimu4t4NJAAKptEni3zR2GDDIe7vBGzUtR5f3B3dl4o
oqUMaiOTSxsYR1f9X4c72T0tJv7e1mmclGuRIp/QMoP+JeZbchIwAMARuFvmH8HUKHongg1J95mJ
FqJM9mU0B2bM6oOUNFm79qL738jt25tCLfbMNFjbB8KDOB/WX6wWx4+eLtwwN1ZyPvth4Sm4bOC1
yOwdltMZlS9cwFyDN+Pu8wm0etaNJaU5QVgBRyu6/dx7a55DgcEHSSTpc9rVSrus/pJqEPSL9Ybg
sXjoEpBbW23nvqwhIMZj6HfzmJmCZJ/YkeMiWQvl0QD6i8Q/dA5VVjbVZVyZCYPmE/s8C4dJ9J0H
Oia0UkpNW+NFoNCbcFlBrxIMwaoimgPpTuySjKaMORGAFyUBJWpkbMKpDMm6M1NnBLoXCt/8fYi3
KTcjoPpX/2zEqnsguCSqJhdulc5wayc35FgE2KkBZ7NdlAkhM41a68gRcYJNAt5YXojpiVo4oRCr
+CMuAbChxNdYql1eRbRNMr39D099f+C1Pg88l9MQqDyb0egA6kyH1DpmHQuEkeD0tyDPMgkmJ/cc
6+jryv1tvypHXD5o33iTMlFGiEZ9wGH6Mq3x6cvGSTZy1x0fsb64Pddo6N2aId2q062B0LswHTDD
5PnVxm7WSOk/y+iQajQAjwCAco3vi9TdgNx6w0+0XnBZ2d5+M82WIagIEE3i8GiEpe1nwhAQl8QL
yMeIpjNQZTn7WbYfNj0Mzrrart2OyDF1LeFMIH1DYOT8ArmqRFa8DdfclxvwhVnNZhAhJvgnO646
akl+XKibrlCe47DSsSYUCiGfO9z9gBDC5VqS4UGDalOGVy338/T9owaTqYLJMK9f2N2diafrYarQ
8wfmpfbtJkjXle69QwIOLBes7k2ot9nv1lEPRunwe7rhPeDHItCjManYEiXgBAFanFcLK+mfG49V
op3XaRD0FB7M4ikM8k5wJ4JtHjUJiamL5CSri3D2modh1zkxaQOK/1nYU+j3F2tLqQrkaGXXlLg2
KXqKh4Lh53iNtp6TD871s9ZZrKUPqT6FENuu8xfEiXdZ9sq4rG2Ncf0U8rRdfDl6toIu/QAwGN9a
LXd0T78qwelvYqntX0CQlN7nJ/YN9y1Gfz1KXcCglIeyPAltjY9EBrAR7ylcdJ3n341inWsXKXHX
GFnkHIJDtVA1zdb0v7coZgWqNKG3S/Q0lYzTLaZe9/CnZ6n/QB7AKaXsGFInzzNDq2lk5ImhFZIP
GcFLtpRNFgoSlhlQEQhgxFEkKLrkGbyGbgNVHTB5irwjf4yzOtI7pJOj3lT3Q1GB18u3HqbgE9SF
9ZdP2osiAUofnT5gvq3es+pT3cgoRiyCRsaTSdrlLrac5V3sgVnj3Kl9VDo2/JcKB+/kdUpI4FKF
m0M+i8Ba9fyxCEtG84cz7iWJ6hpf+7YTJZ2jQrn8buxSEzKl63sWpOCgOiiLy4lBAqrKEYPqU/sN
1a665p5msFDevsksZ93Pig5+sk2xw2Hd8qImZct5K0YPe5RMKdWNVJdskjLnqboF3WMmyoY+dKjA
gGLMOtvhFt4KHY5E2x+khpUfGjD8qZFdP/d9OPxxMuR8UmiDHPDn3EZUe8yYpSwsEMcZBntanV0x
IJ7ksLPSHaGvJ1kzHjQ1RIagaLG+bWcWCJWQ0qG0UqRj7dZrV7/TWk4DthqoBDPrvhOrWGzmp7mP
8Zg4ycDb1pMpXalG3F0V/LetMACiSbyRLZsuBBrvc4rh2feOq7UF5ede3VHOH5LsXZ6e5cO+r0qD
fhLYdezWXQ6hrz2L73vIV0wRgC4SCzDf5qxwMTwcfl2b2HNHIZcjLmiB9lkhHXPdAOe61hjn8yyI
T48YWoadLBuatBGMpS8S2565cUsGuV1+d9LcurkLeNiMV8HnBVJo0c4ZbKPziLH4/WiTKT2kKB8E
3KtE/YWUuEoC5SUArAGK17C4GlWG/A+0KUxNnnuhfRb4dF8KpGohESGVh4tixhrtPGcGUmulNdsL
reFUTc2czufSCfuuHahziG+9NVdzH1eFKl+vA3Hu049Hnw2Vca37ekyA+LEmxUzVZAou4xSM0dWg
JTAoctJhJA75dtVe+kCi/mqHVeNGQZvZty5SgSu3+KDjYEhRqTP2zEUxlE+Mv1dygrm63/ie8PRb
K1MCG3bGLdcY1E8ZdF+xDASZoL6q1/kmHKW/oqqI60Qg4dYa24hB35dSviRw5ullbYG5QYwiDzkt
UHZmf4hdLo+VXdDsneG4xmau8o2I/XXwjRbjPYU/4k1VSfFtaSXx7jHaQy6w1UzUE2yQVn4WaUF9
+ivtCDve4rV9bNexj8QZnIbJFMXm9V/UqSQpwPX/GDS0QPgUau33k5rliR6yh9yHkqcIIIKJxr3x
6nC0mq5HxeZs6HPPMmkpTdyAqCn96ffp8M8bgj2AH8Dwp98qtZqEImEkBAR0pM6Z23zTp8Ejzsxb
WMiaVlw6Q1WFEl+fJxxo79zmeOHCFR4jiDBXyL8vdjCDMlHeh5sw7OUKGd9ztaKJjAr2T68R88GU
w42y91TIEFCO5Wf1E1+ixqkancz5dm1q8eh5XEWHs8Rb+bFiu6HU/CT6x0Uxwn6x1/+nSC+d6vfM
Hg0njGClx7mn36s/PeIxn+Rk7ijlhEWRbNUELx76CrhZ/Kmcmu+ZMpXgTV+dluNAFONTfKvos0Ab
pr/9peotIXekYNXNd/7l08ubDCV7vprZ8bmJn5tANlcqDcXZp5zWopmrOVGcssjPAfcHdobvLUlV
l8hyvltK6xGtAc821dljqeZ9zWMIPLlME8d3KwaCrPDXQ+5LRAqDYSrgkzGbrNOsJpVm9NjFvHuJ
hsBS7BpVFsKU3wf54PqujdAnQVR1uwIC/PIc5WdC7lNMRvUoG1Jrcr0cuxjvadiknbqY/hcRaWvf
4/YAmycDHZNSEOCfzl96f1UfjtlLO2cPv4xHJTHsuFiN8Usu2tICfVdGfmoHkLJIHGg3fWhuCtdE
mX4dIIjCRPA7u+R1IiVbhxOQnMtwEuXqwWYs3jb9cmBoGm0+YRawY9vU32oGupYd6BOgUo6IUrQw
1StNdww7rsP/FXcQs0f9csbvGbDPMNhWFLg/12RJfoo+45SndYQOAg+T5aBgfm+fuHZ++RibrJz1
Vxi0wuShyXTOuc+xPdtlBGrQlUg0A6efGO7pPlZkJAEl//kauwnct4/EnAhnNxqSHSK5deH0itJG
mKon2tLK8NaQRvM+Dzk2AtD0M/YPWCBay8c1ePDhZ1qJ8vUatLZVncO1ubXch5AhDqYfX9Bvw3G+
8RaHpTUn+JSriSAaAaB83IPG84nvbMER4fTIE4wHuHNuEoNS74G8rAsZrOAVFOXm30AnnQGftSX2
ZNUl7OVb8iID+g5MG/4GUH8hiI6ABkerkcdZ/VaVjpJNzmmyrIOeccl1cMw96Ivi/o9HjqVMHeVP
W/Fi5XP2GIUabMp+KyBPJ2c8T6fYWOnOrO7pc9hzvfzIBzmK2MP+9tImjSePDZKPXN7I7NgIDi/B
gZ91bnMcerplQUSPNzno6Cke+BfYG/DOoLkK+ey1Pe6aKA1LHHRC/rcHmOsbkdKqxvTokaoiPQBf
oaIEgMcNRD8xcBp+C4yl1HHjtgJwUm32I6wxyCJo2BOAkoRxfdrEhpQ4Nyz5CLmulKiSGs81z7r7
5CvgJ4xMBk/4vafMkZAxnAa+UCM5Q0zTOKohqbyR81lxQqixp5ftJkdASIBiM6ZUA6Xvd4RZYOXs
OlVy8kwilDx7PWATucryN4oNVGIdZHoH5pMQ1EIJkW4lKrQYhlpOHEta2d7EfzMxgOuHK8ot7apS
e4k0u+Aa52ATgr3wv8AA0loywV0xFnhImiRahfOkljkvXGJG+c63kJORIUpB2HaZN9GrHZ6P6nVe
aM4GP6v7LTMMJvJSVruJbFZe997FhTMCy0oEzg1UobIAh4lXIdE/Jf4E5HOm8/STtkgrtIRCL/+h
WuRh1shvFf4UVyNWuYGq0guWETYUFs0lZSHLnVgdeM6Fjy9XGDWmR4d+5Ix2zpuet/B74JKyg5dE
nipAHBUstixgJblGPLqS38iHBefRJwgJa/a16RJscctRi9CADwQZmsPzOJSGuGXFKMSsZIsrX2pl
DgGxgf0QfNqqfB1XYDfh56PFCa98f1WzR9fKnukR59UoCZIF/7qx5G72pLrcyeiubvfTYRBV8sWe
05w6kUnlOj/7F4PPxY1h0uEkPK477ooyd+ypU/jz+OYD2OoY7DKTx/jCapOoSATxXpKt6Nwq3M6h
VKxp9VAI1kqUasGCx7owAMQt2Gk5JneR8Iq9YNMUn/WHuSwbe2ZT7DA62CSk1TjAEQB5H/6xfKoC
lAOY2Y9ZHv6HMuNCXK+PQ0O+5/vXg1GgcwitiOtohUvQdH3rz0NgRoFsC/hG2SDXqM817jt4LJMB
/LvKZPSr5oP0pZS79tuvptGy+yzk5M1spVCxwC7xC79T5JbILF3ZiVkGWnZpgot0AAsEddx/Nyee
t++DDATVa1DgOZnfNo7ujcxL80PxpQ/5Hd3ckeIHlwk53B4JKzl3pCct1XybP8qn4GtSPzhu5PU5
42uT82ofNV39p5XWO7LkpTP+z0L1UUdIQDomXnrjeWUQkiwWvrlu2sHi+h0gmY5qXkiQQ1VPnwEt
Xc/eQIhOdnYNPPYNZwnHWtfIz7T/l5uPGgT+JAvV5HGmNEpRwPhxBzcKJ3NjwlC2ATYRsggvVD3x
xiXXrBuacpJkoE5kTQdL5F5g233sIkef7d5unmgsSguiVbsfiUvnB27HU8ojZIhHbEfmWhL1IDL/
1nZ+uEt1M3ONUsNUL48Uo/B33lPjQmgl39+oOHtd8xQRm5vQuf/c+2ywcy7/RJ05Ki82dw9tSxNc
SgCznRA8h6MJVmE59kgxqqKKCqSOT4v8/FN0spAttiwDYV9fiPPsfFPt5TPsCJ1BzOEZFXZWrL6J
Cz+qnZR9SZS9s0XG3X+WWn4232URu9a5mzduLm5AAhmfWs4CfRWeLOrehhPITj5tWRtEHktmuG7G
syY4novOmoa3ZkTRzvIL4y/t3y6KDy8sBNZgFTIbmRtkZ7iCCX2+TTGO7rJo9BBlHzcjDYSJBy9G
E9SYxKDaL16qLo7i6mAQhbuU+JYSWA5I5VLgS/qBPbW/3CgDQtyYYL1WoVpQ/SlxKp5ITboFRJDN
dlESE8L8W67Hk2XBuz4jDEUCux/3LF5EuapkG9hhoMfNlphTcSpOpHmbx6yexGoKlibeKfr3ej02
T6ahBDbfj5cYVcCyz94xgi3ap+znO+4yDvjiiq/f7fviXGdqplZ3PAbtUW8n3Hw142+xFrkorkEG
6HAr8AJcqPdEMCK2uDNjYrMqPXN0gEmGizVqwa0vyFZukQP6RAZCN2BrAidCV8DIE/QxIFtkvr2h
2WGLv4ppUhCuHtB27tOQMbGLnjL/Wk9ApXpMrIv0+zveI+LUda9/ukhYw6JOOQrl43NSMbefTKnx
pu90m6wOuYrnI+gL+1s70Kjw42V5eqSIGIyUKBReYmVm+6GsXRCX6CY7D02oSPQbvE/1+u4dzV4q
IIiDgkdeE/29xpstDJLuQxByTi95NulDk0v99svQhwvmy6WckCecRpIz1bn2p4i6YPHDjJUPcQTy
AYDVPYi/X42I1VYtwgQDcMHlDTPuQLUDdiBVseBo/oAO4I0NLQ7VMdSvLB3HwZgzCkDLQqgAFRVp
Ti2yTlcQejpT1zIRboov5INYB6WEX2kfcOx4Q3CPKxT/q9G7sUpvY1qcXeF5PeOh3S5LJEBRLLC/
pVb4AVICysJDw7hMgWByQVzN1LUk8crJf4yBWsNTAJbM+mDDDlksXar1TJiZ8MiFzse9HkQos53q
QQ4Zw7aL2BI56s2zyT4Qyjq2CT7AlyJ6DM89NKjjAp/4N5tr93CLL72bris8inxHk33KPVeBXa+Y
OWEJxvCMtZ03CDT7tu4AiojIq8dueruQWfERC5tS2U1rR0F0EERRGaoueuzY2XRKf48uDG2FmnKP
utRLX1w9NZ6JcHnq5kpKJGtVj1nJKRbwL0FL5Hw5ElmaJoqEQEuOFrwZASgfK//0fmyq7eEIshrw
jbl3OFJ4c0huQ2RnUXG+wNP/RrQOPaLKDkrO4AIC+07StuquNHxncZjo8bdD1khzswCQRM/YAHbc
iuh6Co/WBCFAEXUVV/adsQelo9PLyuMploTulYKOvr7vlMumvroabjRju8gakHZgCdpqvfr++vFS
SI0rizNHTMZY3Nj0vui/nxnRxyA6HqYnvpAbCiWWp4XxVZf4atZfssS1TIwN2SDebLojfoUzhGia
8zYJafxoe1T6OCbl4mnfwsf/UWQhDMTyZ+iEeJTYOynf0K0WOK0yL63vwqmZdkVxPLdP9zx3CT/F
C//hxiU0+HA99MneThjp8YZehuInROhVWQcFOyZu4PJYaSGxrhrSzIp75bct/4a0+KzS1UNeAYXZ
H2kipmtE4PzZIJt66kqAv6z3R6q82Gt9Swsr1+6Tyr2ube1sFqZydTkKoC94WZVBsC+iMNbDPI3O
yY2hdx6VdUvY7rOyFK6p64Ava0MKDlcIvrC5LNSX9bdWpUh53P3jm0J/R4E/t3pwWSHbfR8Hphah
U2Ncl74B901mtrWW4IywEn52phCGq59c5eq+i1qGppDTfCDCyJIHrsGqF5J1+uUedBV7/WxoEmTT
W+VPmZVT6kfvl6NMGIGpn3U6CsXNcUHxOV7QsbOUMlKOrR4ASUGWltMqELoBy//wWQSwPcIN5k/2
3I0RH4NJdNScDLJ/7MwXagVa5hHcM+44GzJOIXCNpCDAyAEztVeT5qfgyR4Q04Uq9D7zKNTrEJ9f
+diN8PHRkq/hnUN/shwqvdezzsBuXrB848pR5RPbUV+cZXxyoJr3h/vcuxexx66WhE7tuXk9WeoV
O3fyH3CBLYh8ddl3JyAKiPrgB/9a0gbUJYqKPS9sTYH5nnftyALJj+WuVpCyo0XN+EBsHdH18Iu1
DI7fRfVQXUcQq6ZJc1zPHwjKvv/kCKYTbPH+2zP1XW0i9NFGENTIIqfPQ740MjlO0Q2wE6xdd/lB
RMbd3VSQFhDuA13X4xhxsGOajzVmwAdNltwFjhET0pYSoKh1ztA8S4lvxfOgJoDCxx4Lt0PfCjVG
WvWgfBqnfxZwjKsWzUYSqGRLnYNwvq6Egq0ewzLjiB9P0101c+nO2yPRJD58XJ/2mHlR7YhyLIG4
ZlaQcUBNGQ+aLeKtXBKYS8k6x4cT3i70waqNLPkxnfFF39z+o4MICrsP4wAGnldUKlhT0yCkvofi
Udf6aP/wBbbdYNXtXPvzMBIpRxFAS9DiaNwwUTABl1j5j0aRxk5A0u1hsqWA1pjKg9IeRGcS/3fC
U8PU9vIImhpRXhli+83rFg2AySdZV0NofkZ+VwIMy3Ghv+6zVcBdwRsmpK8kF3su0j8TeeATr1/1
d+GmonOoBQj2VL7vh3Oi18ZQ6wW6NagtRvi5BJzHNpkNOCMiOOgXstY1r1Zby7b5LXaV1kcYh+qX
/lCxnL7Qcrev51eDX04aAimKC7in1LATnb0DcfWOQjhRKYyBazY77dG9XOnknvsqC6FGc7jH5ejf
yDW85EM5hWIVrnHkrAzCu/aulqN9ZETCBOiJPhnACeH0zRtl5V3245YaUHbhefwVKDqRqXF8ojcr
UYznQwTyzcNbOatTpfb8hYjlgZ394y/B9EBxp2YqfjPh7rRaYQbv5YgxkUByVzikQ/pKB6lTLKDn
tJwWaowmYr3XT22J5t24hFIh8coBwWXbgMJmwrdNl80JY05fjJ7RR4FGfRR08AX9xWn+sNKBRiFC
4CVcOlJ7Cp8ZTzpvNTAsGbMZDlYZHSP983Ni7RCFMd2rBP5XjZifEf/AyRICe2oBHwYKVMoXTLKb
Wu4am+F/mDRKVl9d6OVB2OtpTPRieNmgp+fxCMb4wl4dWvFgUrVTQRTUQP4s2wdj5w6v3SbA0Tzy
D2z7cv26ZEviQoUntW+nN1PfjQkxtz5OEXwKTlavfQaT0V5A6WP+6nxRtmgTZ42th821OwoQgFH4
bwh3nDYv3JO8tkEnle5Q5jH80I2W384gN63mF5t32p+TtF4W5WyopXkcX/INRopDhO2EzZHkGCVz
tP3+fU+a62jiWm3jNzjgJP/nogi2l8ih1P/MjKtH6PfuoY2+HqFw3AJVqiW8LRfjwR84xBUz43ww
l6kTKbBl0eTqrp2dVM4PaT4FaXnFkV5xOzmQJhLZmYkG0is/sAkeYd7irbgMyvltggBiGZpQY+jI
KtglT1jKUSIxdAkmwl92V31Xzh/K2coyu9YtzVNpZisMiKs98yL6bPAfMk3q83vHorlL4ZLpQTcj
BEk/P0RDC2MHLXG2OMjxhjKX8tiOzp37cMXKnY97Xl/e1uLJbV9KbJe8QlevhTkDfUiK0+6LxCTc
U2eaoykjVFv5fyAFe/4jYgGukFWJkheRyJJ8Jh/K6mB9w6TmC07rDu/4Ixl82kBZ5WuRRb6P2eIB
6f9oJ7r/qr/nnDOSnonZhGx2OivRrGbJiLE52KJXn31EWgYq3E1qduzQnLCAl+dc+fTY6Pa9+mSr
NVn9/LM6KLqBI8ihZW3PBY/KotXb0nf2ozNxWqysnnlA1pWFihWMprDg4aFoFQs4urAApEleHDBd
j4vnEQ7yzBSbgaHn0S+aEnymAT5SmqQKnJFHm1USfnhjET53aqpB86k5XPtTxkvlIaRdHa0+mHVo
L4S0cMWHIVkAFqh6KnluxST34yCXZPutGBuxT9usYUkJ+FCFI/HL/eVlFfIT1xYeoDZi7DHCasUM
vRdZIGxk/+JSo1/qohFlaCoUJ351MEp1DDbvsQsIX7A3fuSdJTs7x7lt9jvmFEP7Sq2IaRwcNhbT
x8i6qOV7GjIHOC/SnPp/w1ZW5U6oV3bg2jSDeKGBJSd1I9j8DjhdBURpV+r+6MjMof65sOjigldp
ASfjWb74FX/cjPyC9LGxwhbS5EVjEluwLkmkHJNPc6UNPIadm7cuMaGN2A5QpgksYp/PeUNPBtZy
qeNOYzoT93DkRBrRocEgzZtkL88mwfdlf/+LSL+t/HbIkf2sCmV/bqdb/1iYZ5Stn+yjVue56p3B
hoplDaNSIJknh6rS7tpBWk/90+5ReASx/W9+Ew0Ta8/FaFppGxWZBZ5LgJ75rF0sz0MxxSr0ChNT
I140qHkIHqlgSk1OhUxD2qmP8H1C3rFIz+O4k1XBNkst/x744ot/BScJy+C5L3iyuJ71JEgpvqnw
lHT117iQC0LDiEfBiANKvK+SGEpggczcSTceoKOHNnLMTeT1uPNrI0TYK61QfanZW7j+4/HMr+O3
9FuIMCN37KRSpab0aEAEjVorfFgTE+MUQ7boNFzsRa/PAumZE0lhTtAlGDERsdKJwblCVpzJTf7e
Yp659yd8pik7SDdnwS0oczLmH9rDVjBefMg2+ewgi7NPZxx/khcV6kqBp67+KuNhQ8qbdy8BNUnn
KWlpn7sX6lIuMmgu/B9v++FVlKTJR4qaCh7wA3Q1Hpxlj5U64AWIRvHvGVnf5F+yYy4KpwMC+e3k
AKbjMhGK7hY8QibaNyvLJcKBi2ER6ilCUcg5hEETAP9NQtjVbTEJjy5RYuTTI1avT5AeWjDmdM3j
Fqxu5o+crEMpDXkU8hIh7Kl/Jx+/ZHYFo0SmZh0TIJFgNQ+cKBV+nn2PYnPc1v8i0dStpfvRgvqJ
bI6CvSJ80gFb7dRqfy1PV2tpS+o2dlO6TW/QDnPDxJygmZx87YPAG2tljYIZDKTbGiaqeuhjpNw9
yKCRLPtNtY5BxAwoN0Qm7g2kKadJjU4lO71KVt+zU0ZDRPF2WHL5ZQ27TpHZ8sKQJeYJuTqTtJWP
AiLaGWlT1oGyRWXaKKzCTgzH2tJYPQ24dPFYsH6Oxm1buSzF9v0spQe5YTI6vTDZxztaQS+ZHStQ
vx4NMkhmCKqFqZ5lY2MY288SRYTZC+4jwS6HrhAfgJIeg5Yn7vnelhdBO0u/7BzlqGKo+W0Im1dM
+e/f9g5/fNOp7bcDhKeV0muT9f3o+TnYUIHJ5N2ScB7Ugl2heG7xtkIG9uQ7ES+QbZ5uBzEzcNdl
6HcNkfAgpOMt+DBFCLeMbOZJ1GbbYZjSYdcSI7hyfrzvw0bGkEy5b30L3zUVwbuVz+/xmoMoeLu7
3WwwDIofiFJfiJiEcb5l4bgKjoVloSEtPF5w/AusMCmID8Nnm89QclnzKy2n8xYvWGmzSNMMajlA
DUnh8qT18C1DRFcj+doh/lU5T69ju9tkWgkJXq0Lv5CQQ5fvnBFP+mU5MkhE0EgdWy3oGaXtinLR
ZwdK6WKtwblwJx6dnKnmMnvYZG++RFHgORmikk268bLjYx9ka+ObM/8gIuDvRKt9MR5REP50MNXY
EA9xVUQfNsZk22YgfTDEXkGFkJ0PXP5RFUYBUtqAcHpOzDeub3dGYN9q++zbEyj5iIpBRshnJabR
X4agOwdld5cAWlPrsZZX2nI/BwFNIlY+kkX2DLKfRMZMw+MxbNe57djsmMyYPFlI3ePrd/dduXtl
d/wHVzHoCVO7Vc3UOoJvDMvdwVxouTsEzgqzz6PKW/xqCGB55yykxZAocP41YIt89CxVDG2xSVzR
dcyRtWnWDARztqQg4H0zXa1mXyBliY2yE15bEqDg4ety6QYV24/v8XFeRUSmUqYuTOsr3Zo+wNub
bHWoPGifqI6jN0VXviWxQi6dgCApmirakoqY1uCzJWQDC5zT7DhxUxQSSPDptgeP+xTP71uw1PQ3
sqEiYqOROq4baUM2ayUgAUkQ0Y4Dc5e1oDWBKgLcvVf3poAkjBqoNe/OolMVDKZ5uynBwUkGJj/Q
6se82AIg0IO1I40zk5kaCSW/TgfHBnoikN8ndViYAoDC6C9Gsj+REyjXN3U4XZIIl0hmZHnrMgl9
Z5NO4gl+muepcnf1eFdjZYZYpk5Yy9S3W0a6h9vg25zgB6GLCctBLi2MqpIx1ENYsNE9p8MYT42B
Ch2SgEPbzsNy8dnk3s19GPtdXerNfqA2PTr2nWQMyVPWYe91dkNn0D1bjbfAvjE/vxAsMcY1LbHK
03cCGruMg6b3F+wraFkaoiORU4KOECJF1aC9rwrm86KZaFB7Uj++KMrwWius1f/shPbfDDwS6VbK
9g9YM+r3K/vw+vl4G2FaEOvqMvbFBtfaXBWnkRpdzV7J0e/mJ9W1+aXfsaxw5DfLFCgrS4JEZKPG
ATcZa6PBdtjcbn3by66+daQcBTbpsPov/1V/JvZnwRHfIl1wYc5kp6AG7fxnJbjZ9dsTxA3K2QEX
OsMCHHQjsOzOeX54t8KXz4IFMGEBd1jsJjetiF/DRX67Y3yHzpRlz3fisZxRqqJInmmUZpi77a0e
jQdHYd/2+M1urTw9pjKxlWtwJmQOa/3wYQXegYZWV7pdPSM8evjrZ6oYmfwWQ6sw3GqiHP5MkJjl
/FYiaIdPwk4HKIXmxVyUAB6St4rrFhYxeeaJMxhXGRj3Me2oe45pXlTIHdt+WqNF+MojR4LfOriA
6URpGLzfUR0UBV76Lw7ZuxwajLtdul/vUBFPJF1sLAf/RDn8gE3utSAgZFTqXIEQV3tOQ5aFhFBk
Lg9XR/NfLQEDIo2s9iEIQwQkcHZNIztxnBI2fvMm/T/kLNUYa6oGqE4YrSezxFBqS9BB7W4gN+39
dCU1Bpp8knobF/cM/wLAdrdZ8o4UL72pD63VNoy0kniiUsM3twumNs1Wo3GBUG4WERV2Gfom35pk
y+CrVwhsWKz75C9Ygzpm88qIck4b0QC78s3hrxyfqt+Vh6NqfzfgG1a5GKaqA3RpRTEhdh5KyHPO
1tFWOz5sDjDMtaY7QFnuqvElpYQxvzXUXO3lTQgSZQ9p2pW47QeP5NYHxFyN8histlXoz2lLLjUL
WJ8Vce0Oq5aR7jsnYtJPztf15SGkF2wdgPaRsb+Q86a6zcWi0ah7dFQELrpI4xZL4z9a1Purwdlf
IqEMd6sPg2lixbmBjIrqtvweqtye0zvvQH99FC8dpzKD7RTyXg0NdOh5KkwLUs0eMh9tMisJp9sg
ZFnIMoFIi3IaYst/fwugb1R7y8U1CC83kaB1MUqX8OLmAmcf6RXCbbwmc9JVl/dEw7y/XaSih3Dv
0WD8hRQq4CwmRY7dE1x3LP8RBZIkuPDCJfsBgIZXyilKjcHzHDDbitTtpTV5FO0MGMaxuNFEi7CP
1iM2zHFJdmHQD6/c9joOSMOyABJmF5Rz+igbr+2vilYVv/JUvbcdTUDLEUbshO9AKi84PULxrs4Z
rL81uBUGHpZFgP1IghLS5qflA+22dzakl5zDhPvtLD04EMU2toCwzt0cOaiVXzbug1wTPJvozoI5
R7mFZ6x+KM/6GUOwf+jjRB3Ak9mfdt/hCgXWVn481VptRiV1YYFL8vzO/p2KSvkSwTgP/yNGnom2
HnRgmd1wvYWbUnQurFSMwEfBNsNpf4AUuVkv/fRpVza8gX1BR3od8SGtUGuk+mkznDwxnh5Le+/B
ogpRu8GCn4JAkb0n5QcthqohWJoAun/RbX2EQOyoZbn0l0A4/tzJlxL1R03gF8aIZmbMTuWIbF5F
02p7wxQcD7a5AdInnrvCxaLG/SVY+rtEcL6dAe88dsZJfmqpnWvOcmou6MVH7gRYRL5a6Hdzh/rL
No2rc24rlA+FGc7CRmOMLKDE2CVMvY1XcwXNqanRPIUXIe16D9SKjGgI7WzXjJH8UYiqr5EfEhxb
Oc12zXnnjsridsiqJVdlaYBHvJTbsT+pMwCa056JGlR6NZWYcVXYZRwnD6cz6z3Kvhx2zow43+aI
4dx4JylzAJF+s5WL3OcfSPw0nHCczY7zDF0MBIAN/v7iIn+KNm6es8Kp4G1Mz6AcvKUX4c8kBy9h
W3PQNDOUpVmWcqQvmslec7DZJSUjLoSaagnVokVJo56Ig2hqXWeLH6ryg3p7muF83Om34l5T65B9
o0XVPlrHppfTeNq/urgc2wdvgEJxvLLJMr2cv7SBDPsZ2sZ+VgosxGrXvYkExFCvDBTf9qqVAq7x
SbYJE2y3PWQ8cv6hLCW/xpBCyk68QydHdlXF4bqmkyHZmHd3YRzlceMkTaF/8uvfOpPFFFFt8Ixk
juU8ozfQ9evTo7r4yrcvkXj3wJxoggF+0f7ycoeDwsWpZWoReqO45cxhkmyTTcPymc87PwZG7Q3W
01ay7dqnb9G8BWUBHIZy6qZ3UhpAvtuJDXIZyErEY4z+asLgzGMSWbiErmHqTrrKn3lZX5//5JX5
UZ+FfaNYQaTkA0tlu3QTSux3bilyCaBgb3cdqV+aDQfLASiQyhA2xXB4YS6A+YaOWWzEJvkTNqgJ
9wQUb3aC1KnDckAOsO3+V3taE07CyTX4Vr0jdYDcacKXk1WidIRj/8Y/sKMBzv2sB9FM6gL9O/Wt
aRKihOhBxY/A1XqOH/JkioqHM8NdiJ2Cv4foselID2x6uHM75Y4GV+CIHM3ea4Uip3U7D/3CsI4S
hyDKkIE0Xy4aBMoAI+B5GZFuRYAWpLzHcGNZKjVzUJ69c9YIdlkQoohs4R4SFvkND2SpzH9x/twF
ZJ7ay7XcXXcceQGxSDcYQxDgLfYv2nutI6T6PeVgGjallJX0+8ELhyMfPoAUCQRY70aChv6up41U
I9ZCI0gVxOl+ECxKfRUd3kzxSExV2WEkSHU63G3BRnnxh9T9E7uKxOFAibH8RaDX7e1uNapBFDDs
xXsAW4hXHltBbqTTMzgQotcKAklbyzTJcP14W29OoLoBpWUuWRLffoufbDuX+yjbnaUVHbljO1Qs
jGMo9ci151rlDJU4tJ531TErR8YpIhq2+EAipdNj7fhjx4Olyy74RuB3lRNVu8w4GWPkDvj9+Gwh
fa8G8Trh1ev2chuxnAyk7nkrkUiEIlhLVBu10P3LogH8T2ymm3HDtg4DBOoL13jJlnL/5JUWqolM
AICN6e+D8ttkc6UOo4CMWwVdguYSwMGPSKCGIja9PBMj+z6yN/8BEDIOAUA41FgwdstD98kqzjFh
mMLwn0/OBWpvbdtoYTwnmrzh/ZOAicodT6Nei/uYS1L3Bj1nT4GRk8ghGiZ8lIxwPwInIhvyfarh
B/zTzQle0g52jW23IUFkBmwfafKWFRSIkdK72dBaGuhJwZPavMqESVLegEdmrgF3dDlsPSEc+zNn
Ukx9oqAMpH1RE7EKHNlYSyPcoo2scSjT31W+zZ5dMQsC53W1NqQqA5iP0TlnCJcVUvvLkaJg7LEi
7iyoE/VJdtsH11zVQVumLwXG620+mchVzmXBGRFfvFMjTgnrpOoc6gibsPHhcXUE+0UGT6hxcITa
dsEtixM0efFwO3V+LAdOBbtJd80uieBATvkRmNpxsVbg85mm6rZGQlFJXPTLaSrC1S0EQ47LK1J+
97zY8E8TcrhoTzUPy/ixeHPAv7mqUwmvfIvQwSalRUsJ/SHEaorDKoz8NBM9d4RfZEvUwe6NjBxR
qCvKcRsyPD3YdJvKU2R1C8o2emj/honBi/6Jj5v4uZ8BeAkmqg99C2b+M+ohu+VW/htm2uHJekeL
ZLkjp8NcyyPAuh28APBxdZ6xP8VKf5ZrXB/AWSNcSbGTuPeQX8kwHC3zg5omr7JHnWFZejvxy7OH
66xmJQVMo4esQxIMl0XHtrjmeqTBWXU6FbDgxGzMQ2PDabfyPRNv1QET2wcvUGFWhbS0HOXtcprz
wf0fRMLxBrkJVYKty/jHDe1mTSaPAD0hEs5+a9yRvrJcgWgiTkn0VLxWXQxAIdw5AM8MESmVqTbW
LXCP8U/loiICviEMf9ncVrHYRKVaf6CxoFYxTpdQPvk4MliYxszFCmObDQLD/1WzamdZmCZk+2R/
PIEX937o7Wg8MUrtoAYUrqGJvLI0Uwt2ra0L7JKcZtlutb+oNn1RstyYYcd/cnnkiq5cxx//rLIu
FzED0Y+xUtbbCS8/Mloo7XVjUiiLgUsbwDoU+omUtsaBJuZTs6SyHKzXfMeCCRvsnnrnLjeXQUbN
aZiFvb+we1uw4SF5PcprEUd8qGFG5uWqUuWLWrZhfgpLB2m964H/nplYCsEz5JGEM+xtdD6rip6a
52eWAl7MYVOiWvmIogDB9IhEZSLp/o3cUsu5nICpJ+lSbkfwEO3QeLGjuMOr+47bg8ZunKZp67kx
e1mK2dL3LBO0ULLdQ2Kk28rJiPXDjqvuLqfxByNbHtWenuzJTf4ZPAmMDvVIYkSXX/bXvQHLUCtt
Er66S/htf2vFRPQWs2M0Y2A4czzg9s1/LTGYTRuldmgO33S1WbMY500yaKeAa4cJYPeM+j39CK+k
WtJXKQszAhBGStrdIryi1Vgo3SDbv9xS25CG0mjF1V5GGkJEKX15q9slHPLqX98DMKXzA/7nBlSq
2c//lDDW6DnYsnoAjnsrji8VbNdVfLJBp9TWTduaTYXryZd0QwmHl+zSAqevgi/QOHyT1t0kmlXK
oF0MLng1S8LOR/u9xW1sITn0TIigsfNOybB5yoyiNJ4FYLEz4uGYjlPjelYuzmojAz6FXNS5hjPi
nTqjdQA+keIvxdMvt7vVH/PPrRXnznHPRvYiEZGPhwFPEvFQ6A4Q80n/QfD6AUXl+3E+8L/9L2iM
9/HOzAEAgIHHv2Sh7K9ppjKueIJ1ji6SkJBelwjsC1e6bFxw3p66vagLqvNzBQbH7ltnoJEbyRTA
sV+fFpCaSXcs2QC4BtPpKIZL58lp9UP/EIXQZA9pDErfFR4dApumvYdgGqe2oUHvQ2rrc1qhmunU
U19RSmlCaNCb5WjQjN8kzyuwsC74THfsaXACJbf0FzYC3HLs7LAWDeqiK3+Ig3g9J2UAa72ffl2/
jHh1zxF0FWizhy2nc8TM7rjKEFrXa41eS5dNpUJhMlK2Kq7qPrb4SMmdew3AwSfFnaCsaorETQ9y
xUqZf7zZ9at9TuDF2oOyIDN1zlIM/OjapXcg9/Itzbk6zR0PYDcVZJyKXf/kLusF8U2fK56KByFI
e85zLZX1NKD8aleEKbPIExTzIFTXhX8PcAc8P7qfyeJOc8Fnp7shri9zDRWHUjTgQRF/RUm39859
FCCNvA+Cj+FBaBHXtP1pjd2uubuyUN0hvcErHPTjkb/uR/ik5+MeisRkmlKAUAv271QyX01xKaVY
AD9Ck+KqENoajBLeg3aGQ2Fcgz8wjYSJyMWQ4MKCoYnAdlTBQ79yEe47Uk9sO81u8EgIzuVPklic
AMmbCL6BuXPEv0KRln16MwGzcnk+spbmzQeeQjlJkgc7yi2RWBNnwpD2UoOKZQQPN0Oam9IWxaLb
6oI5mCbnZlTHGxU4v9VoqdNq82azWYriuQwKspo8rQBUUX1F6ShBvkoQrpL2zg00kF5qVe/9+JIU
djR4jjZdIl2RXdkAGcdsDZ8rJGneLzKDUU5uTTXlPMi4CCXroJpME0+sb+MyporUoXqh8z0yxcuR
a9wLLkL+oSTzhwt5fSrLFUq9Sfwrd9RIpeU1TdgDTl1xhMVxvD41FcdN61izOL367/raI1C2lygY
6ia61+7Adv1j7pvLKYLHJuju/hvOLnkRMgTiwZ3AI9Z5/MUUZZWg7thV6Jn1qdY05xf4e0VEa8DR
AdMamG2RqRsFSOlEN6DWaTPmodbUayQPZdpAhfWqdW/FeDl8BZtftSXzHWqEY/COGhFInIVk34R6
qUlblnMbYfGXfBsAXhzpLCld1DM0xuiqosHZcs6gLlBVsd+LjGsMvD/0KBrVuXQa1Jv5WMcFchCH
WAMvn79Ix1MfKfDcL4nIVugNWholTN1oAhXdJhnWEUU2Ul3z3kQ0N1RV25c6NcaAbHQcC9GPgv3u
1ve3CE/1773hBLxuMxto6zPP+ZgWcG0pZzuO9wnf3mUQaotEm11oB0T29ntTQtdBVM4e4l2Z5GnT
wdmDGOE4n3UYzEVQrZMweq8k7xwz8frqTHaOCXcYVDk+cxoaCV5gJLi/WjTZK6yP7l7QeD4UjA0E
kjCABLvpgclpo0MLhys8PQ5nnXfJdJQlWtjYAUtcwG62q6RUL8E6BPaDT2VkaLKdyJVNdnUbq8JJ
d6JAmeLhMvKmsKz9iU4jVjWvhKE2yjCgJBpsNL9JXm9W7fYwb/5CJN8ArT98mDk8bzUYlhw1hpBB
KL9oPNk2xxz7jW3SLSECno7chbMolZiq1OOuim2oBwm+HnjegwOT5sT2sHcxUbBdm8LegjhjI7O0
Tzv3lFKb6w2t2tt11wR6l42DMP46rCHewc8FXeZkE22J1UMqflfSG5HZXfXdEJHackqPR1hLruhm
piDdsuKQBH2y6RQSlRlLsF2KyjHwlOJ4WvqA+wkyqsxH1jQeXNJNUjbu5AbeKzcQEc9cwU9obusP
QCzevgaMjhq80JAfGRVte67lPCt5bbkJxz2WAFHY407mBe+tzcvXacyi/mLFzbnSD7q+oQ2HboQV
Us06UPu88u6/3gRUFJ1XmoOi8oncm19/7B1bJQ5N52ZEa+Kv03AYEELkV8h7oIk6WKvDHlKsqzey
eyULYLTp/OVhBoUlxqru43YQLjntBZ2JCPLUlbfmK+7ZklSZ+hOYJzwq9GLJnVV+B7BDaKmolK7/
AX+EYJtph9kVHxRJN0QCKZS2OwK1S8Hb6znf3dyHrRrNZI0YydHzB5ES/ROEs8FTZog80dd/26qC
5vf6ZVsV8XcE95rN4iY6brpI5WD4OrwQeaE/I2a+HRVM6sUzqk0obVRtQgGhJaM9pTlcIQTkH0LS
GNO+PZ9aau39g+byBTQsiZbJHgxvSsMH89G7vh8sU99pV6XSa+6LOdt7BY4VTqbV9z5dv8Bl4YE7
mbCzV6s6GvTCMNpSJey8vMov5nkRaRu7JIkEOAjXZSw9XM1WdyJpX4ewpWL2rK0rsMwnD5+bJ/ah
Rj9D5dOf61i88lhirzod2V4ij3o/5H4t/02mWDCPtexF0oe46CM000yX24pj/NfrBA/d52gRaPcL
RE8mKavadkX3uvAYzbhhO1I53QnZYD41XuZl6BWeIVEyt63EdDJtwjqkrRU8gzaMuJbyXLJBZxyz
o5dQD6S4miuvCU2v5D8ykJ2uUeelVRsHWCJ5KIHbKRnAVlPhXKHzfTvdBNJBEV8ptrxUsHjQ03b7
zvfDoLXKdZO1PegR6h9PbWOTD22TGvBiSzrvLnNQizYdCkZY/lMBTZ8xfACE5kc+OvCEBnkRU2ff
VFjqCV1RY5WWVL4RHVUgVCSIuPyVcttOFGciRNUjF6S/oJXaPfJiQfzDnVwY7frNE2OKtTN5GC2D
hqSEpPdjpZ6jmrgwlNdDw9E+gpitYip1t+Opco87pdf85Dhs7LnKx8NKv77RRMPieZ2LgAX6vMy1
drujk2cNhiAkZ/6snXZf7bpdjGe1CNItBtjcMSkhm1+0mcknlRjfLq0ktq+yU94smUvjYWnRfADI
r3efawnpRra5NjJFpExSjNt96jfyeve1v6n0OCkvvyUAx9/PBp8qkXlci8+dHksypYt3Un306UAl
FvUwApzUu1jRKIARXAJ5uMR1XLWrF5/Oh/bxKF9aMPw3tmVnoWAHGa4UklGGlmE4sPXA7Pg1QIIt
bPAP6zRcMiWyrsY9WO0V+KUc/3UV8akMIkLHViDa2fKDA8niQzQEOc8SAggEViDnGD9z77cMW8T+
bWDt/nebpgsD2pgX1uwqTQK6huzojaExdrgSgPinMtB8DnCHNOALI1BJNmu7LEkRbUqAQFrVppuf
Qux4WbW8LxZgRVQ3M4XmDr7c3gTo5f8H/ukYhD4K8aGDzpAU86sTo+57U3/xx6k/bHW5v8QgnGhz
9hlMYB3gVkJCDkStBpAIzZkGZ6frqNHymVjnJjVxWPMN+0EXjgf56sdgBMAyp4SdeksrRJCBSnER
OOdCRnQ16Bst8G5woJRKXbeyHwhzkpg/EMpfnayRA78fJJ65EbuRf/X/nBmAWv2atnQNRIfWWA8Y
LGzvOqResJzcYHeC6FgoZAYewqE3a8Yp+pGc/pBAjIhzvH+MC849kefyiemqJEh08+Ez8EFfHxsa
QrGCgRPdkD3YuVc7JzfKkFJRVD9TvW1Wv6VhT3eTYggXy+K6BYIwkTuO9CrhvyPH/r3SRRMUcKzf
/GaQ3iTXoFIWQR6w1SBZg5Os7mxzdEM8KnZLT65SwUO9yx8HFg5ikJh/ltFmF6djXFv4UXvxWtTO
HlvDCtWFHwJERhbZG0P4cby+DuiWqJ2G2KL1WAY/NfOrfVUAr+zq+BxkklJY2biwkYAEBvPMPlnU
6YpU/HMKHJb3H6Pm3a8dgSHC5+l1H9P3VP8G6rOdYzgeE1Hkrj74CzQAf9TnEbgJ7Ak1XsZqzxRm
KS9DxNItbn4d3pjofPgriSLkeZEwVCooNDAeLkm4DfV+XqQqjhsLxaMlxNpuaRMdhZsHiDLy1oRy
Q87nOlX8rPelr7gi6nYDGiwEisf0/3D8kNt/mq495MxnvW2AcWT1v6N3bwyZhOIpyb4E8fOQe/fu
KgvavKW8JatBc3Q9zWm4+TcTQBu14cWY/BB86s4Z7BPwpW1mrDQw078X7sWW74fL4VEh9lXfH0ZL
IHcIcTPljzI9s5+USbZ+nOpYevt25VmKhFWSQ83fHQeLxP/xxH8NrHIaTnZT2C2J7XBXNA3EhniJ
ZAhxfb8qaF35VnfGlxPnPUobmDAYichmTzZ2EiGLC4thoBXQFkuxMB6vWTxKwh+MYWHhxzXr7Qfx
WOvDViDiTFYwIG04IZAjhZsmuXQBZK3YFN7m/E2UgWAwaQWpxthZBwo142HK6dWSFGTAHwCmrQig
P6qsh58HYtYHRtNCCJBjs2v7qISPq6z0N2TxnjtcE6G8j1dVVTwvl4vk3DTPk0f4T9opaDGJrXUp
kk23t/upue580i97/BcLKGvZNbk/M86kZiL/uy2BeJuRmSW2qCcfctv9PL16Uxa0y4Goo+kBREi4
h3ro9uKHNJyZi35c96IJPUUD4Gol+A89aaTVHZGeftIqCOOZxVa/8qWv1obD61SuRS1r2gTanR2Y
fgeRY00piNUA39tnlVgEfblJl0DETKprQkcIyjjchcheBQ4YsG/1Gyxjon+T4zurCHAZMUpGogPy
IjF8xBcrtBJDE9DG/p0eDCqASt7VfcJI8l58rOAi9WQtgC/L9JCxDtBnO5wyjASJO5NcZ/BBarow
VCfiQcC7EU0SqaljdqbCVbyo9zbj66pC41Fx2XB7aalcDxVo7Lc08JkbZuixfwggoUJ4hFacaPJL
bo7hpEM7YA34P11TJyWtX416SptvPdTyoS8rMWJf/syesu5ZCb0WVAtr0mbpqMfdE/BNag3LS5qV
0Tlg1b9NPDwiwDTm1lQnOK6DlpZbuTxpmH3aHxV4+GbsUnbQLecpkXfjQunaMv28NwZPILrDhQ3h
Wajdj0blM0zWLcVM8wl7TXcN3KqYq3DNLZ82YbXiVxtf3ZeaM2kFJZPjChIV2obTcgUGh7NvtJuM
MvoO0Swk9leBrve+MsrvSik1BnR24p4f0n1/syjzyJ7F2w1fdh801b0AkJ+Kp5Wowtl/jzwN47C6
Zc1uRQGSrWo15Dblb7Iup0yw9fF9wf3MoNzK+0xGxi+POu1EknRtvX8xVzX6B+L4ZknsiicIh+0F
XzEHY6Zzg6eFyUJB5sOGRT+TUbvntkD6VccmWmE/spbDgY/UsoOpnSq7ywz+nKKnkUAgMR5LBm6I
wn3LwSQ7pPCDtlW1TrQIxJzKVdwHGXvKcmrNsJUI76jGQ2jIhG/VQdJV0Aqe58fBkUcTCL/+NlWa
zNbIyr7CMs+URfuTM+JY+vh3q1+rJvC2Kbq5ymHUAbhB/3iUQhU3pfqh/+XG5xU/DmD1ewpdWKJn
hbIGunbOIJNFXGxr3cpiBFHWA25OoHQo6qt0a+yd8S5KLLxmQ7nhYuK6QF8D6LM7qR7LJXg1Hb63
WkbnKRMVvVc8zZGmg3fYUmXEP3Nwh4Q7Bin971FhkcMJA9fM3CvNyFOw2fWQ/6GvRjlFtIxMDEiS
Qql0oLJei+7riabSrQ9mZgYXvHnUUOgMciXVVGsQmNYzVv9M7BZN/IfLwWtd5KtmR4/sbS/SoG+v
AWnagEMlxbFw555+ZE1R5g4TbE0y7x982o8iaN0FuSlIiw5TkT/puEeY/hLdxgBadHZXEeOIzYQm
pkXRNJ9CWMj2njVVbDRItd4SaSLID0XJYxOjKZ8lcL6a0RoelqNaoN3CYNUd6iUF3NvBG0tYGASZ
R4vRKztYzvWNOjnYVFDLtgPTrkYlXuVoMxZv3FMbZL2fdWDZk8yIgCM89FNxtdTbirC4JLB63jqI
yvfoyQawEN7udh/HzBUTCAjBX1siD511cwy+MW+TN4FDIrkvzg3xxBO3LLsgBbZsSyRTk5Fk/Dy9
42EBiuNg6x2FYMKEKwMpVLlRxI/NZ4w9W7apgCuTE1qyVbRaANXjB1NuAZUPGSMhsAArVgKDM3XP
5xKJXQyus8PAZYY8MwP0Gcsnow8FktlxA/ccO+9xS9Kz5aIBJnGx8jP63ecPaXsDnWWfgszLNUPu
sMq+f6ITV3t7GmjeigAJZo1Ka0akQoSm2yw39jiMSjq7EQmmlRey0rsDtsV1vJ7nMi14EfPnurFJ
P9k7qcnbm3GmIL2XnkzSNipGQU/T84JQzPFv179alJoz+/97bNZ6DxwpRgBmlmfLga2ah+Z8J6j7
V89RxDo2Jz3k+UJli1B385pPUpzoY4gbv1Iz/EO7uEF32xQ6XNeIk0GNHwCLbFdq3PHdD8ECMs9j
2eEpVosRETNlrVEjIB8jYh0b4n8ehbcT4IcyvLvFpiboRM6iNw8Aohl0z04pOHo7lbbVxIfs1udE
6KK8iAXTmzsAuHDAbmZAku0HBxnktJZkLdQMvPATovQCKBId/1Ox5WGTIbDlcU87RGkeVLtAF5JO
2Quz4IsG57Dl03VEQ+TnFovjPrQIUd9UaoESmtuuz3iEg/JiLfkgb8rU+1IT2mvdm6u8O0kigRYh
vBeejnTnmFRMqq62MX+Sy5iUtpBsclJvalwhM0jsw/4tvg2hPrnYSu/czvwbp8WaPLk4UL6w1FNJ
vQga7t9ehrmYu8EQMk3MOeyY5PxbI/ZDBBTNc9cfInHTtKxFnC6WiQ+Cz1vLGB49XIVojCUCZjZV
HREreFeyycfGOW3bT17phCm8jd0hEndp1gNTmqexSsKfalxQcnp86XLm3rOyXu4XF2xEk7LO3Ys6
YfhB3rSzXf3T9gpVyEipilWLoOVDZaQQOienKXG1x7QIqmerquipc+YFM8dNKwmlHlSvMqjrDotc
/e9WsaIiCsJu4fnRhGQGuwk678cWVOn/zxbr+9dPDyr5GaopQl7gH2B5yQ7WplbFsH6Mun2o+M8h
w5SM3gfpLBhOTR5Jw5DTsBrSXRgQVUSxkwuO6dkQv6EF7VHnkL1NGFORU0Z+D90CgTNXiahPRAVo
LYxBCDL/RGwbybs8YWr+/wL2vmV270ewZs4CqM/G/0152jG1Wi+rPoJ91os66PqRe7nQAjdX8ynO
0k4eBnx49klcB/SbQceqokuIm8z4jPrIks0N69ZBT/ZZ/R2N4kvdPlcDYC32fdwHSzq9bnvTiVnz
T9e4hm34TvrpWDWkhASnAd08uVWMehc3w/VE2MIzDssJNioPO1hLbo3lLvCX3YrBsRN3DnkNL5bp
MRoOcMBhyPjliveKV8yTQMLtlu26R8n13mVrJHsG2M4BSd94BnG15ZRA8huvpoj2jncbXpOmHRB6
EmRBo2P6+fPRKuL3qhALBIvk4cCMRNOafpBt3aCPxAXynE4kFUG7ExVPuFynBRQLx2R/G9fSy85f
RRbLJJbAYne64sU0lSlDOIHPAiXAmeDBQqnf3NRuSIG5yIxw+IgDGZkc6JAtduwuEp6hFjt2YWE3
5ey7CabCyfaqKbksaVL/KPBdyzV/psuYM2SQOZchL2W9HRhe6fklsD5eE6TTkbEY6VUgE8YFQp/z
m7o3rzEYNcjdSigPLYyYXkxYvMmVnSLobLppSEnCU8/iC1nHiRWMVDYW3UN/pRqxXdv2PfmQNhBW
T4v/xuW0ipT9Mo+ZJNnkh6oZSHwc9cl5COj20yzPpmAOYf+nBsJWXVtzngBle3/ItVcdFhfr8eRW
zti3CUOwXvjPAQcgOfs8OqybYc2c6k1Vd9zTIo36EHvGcVLRzGzQMHa5fyTH16/FzPxRiwPI2+Vg
qf4FzbQVcrmnb6A01RkIy37agSpn9Nr3F0G9b8v5ykuFpnYJ5FcWbJynQxhFYQ10zaj6yEL9joEu
sKZomkr5JnfPrA0BMi/8EErwLCmF71HO9I6eOHD0QrMYvEq55LPOxgw3U6e1ETf7GaXdiHmkd5gf
35dN3yzqefP1N9QEx1y99/AvVr9WSCaNBgGRB1O9LvAp/xN5bYV1ZPpLXxGEQcucwi94EwG8UE6b
YXS4VK+I7OoB8oHljB74ckngCqreqS3jNz1OsY2F61uCi3vBwVokuhN8dqso5ivOXkW7mQVVkVU5
HTokE2Eiqymfb75gGslbssifWNPWSAxC8TDIf6mzufb2AEsA2tfqlAlni1H6j7yYl5J0Wb1Fuebh
WhwMyCDImhfuJwdq4QlvGLWtQEO9vT74Hkpi4MRulrhTolY68425hI4yNL1cs9aYsriEw5NJ/mni
RAHgk6pJVpMKVuIyF2QrxO+cHyqWo2AqwEstCqhQcqM7GHMHStYZtqGSu5BL92kFkArtv8Y/SRoU
Lc3iAVVjVHn/oSUdOscilwC88l9SbJKEW1YU5OfeSyBEsQZyBrAQd9r9EUKx/YYmSXxIXsKdoL48
jLyhLH1EpyYhWmfTqpLGjvCJx6SmtjJMtc8olIivK4ZDl/jgAcXfXevWIAu81XHwNBUpvAU0zCdR
AXHiQG+w6sr9hNuGbsX+y5zFRl/5RZrw7c31gwcmtVNkgB2bpr5VaXHWMqZKRALz6XUdnt4+txuZ
pZKT76iUzsanvuISk4h+fGOcIDRibum6B3oNWGIFN/6F1dqfFWvQ5mNkA6UgwuO3muN3RHI1WdMG
5FUsHtx8tZdBbptYBfEBCSwmKIh4VCofs9lSotrvsCJhxoBqeNZBUhLBBEby5REgeGHIvlgZJucK
C8ccSSYtbI/BtW/x6CtpbXKPwxL5BBNoEnWApAul/dMYdk/Zwmrkr4P2U5KjHdXYFjPd95kNMOj+
pZYgkI0nhH/uMvZ8ocTGoWptznUgHxE/CLtYTcre+AE4To8ZOEDyk/+kIpKbxyElD93NGDK23J5I
VoEC80MhPrxq2LJFhRZIcn/RmJ2/nG/CPnDiuiZcNvzLzjcJIYM0PfUgdgzv23Oe5K5blPdM7IGa
VSdt+yTaWfWK61i0pMOiNyZHPdpDnyEotNipUvZE/J500S5oc2ZzF8ch1Q43CTYeDM06l1j9Z0FD
1nIaT5AzAtDMB4rcfm+eR6AQtOKKwzeBr28F70dmc99ffIAB4RHl+DbbK/L1Q6vQ4h7zSt1qXg+B
SEbTbvbC/XRsga28jmlrssaP026HihM6YtyuuqnKoNMqdtDRfDSEYw23CZfNAuCB2d3593v/bFyo
rPiyIqNFKIL58OcqvDks0xHnRtLZ99528djft1ZZUcyw67C14Oa9hGqU33dpSv035ZTWkRaePVOa
luYurduBXz/2aJQgXvJC4MeKvZ9j1PGO9KfFrJTIw4V6PQ4UX+daD3Zt1NU3mNH2N6vSdLJweuFN
V4c8/xTu5Yv7uNknWeqwOGIlhBujKXf1O9zPnnWZGhwi6hzwN8ZyUwpG0kClz36rHBWfMDAeFQbH
/pVtMyoc5dlaXL9EiKaA5NS70IinPIa4s61obZ9UExFO36pb9oVsSCRoZAS9/JHDyuJ5th0cTyDH
eROH6KZCVb/tzeaaj2RNrRHJquD7YOzY9Ow/omdwEYv5P4V/h65P8uOvw558a/URPKWnScdevbJm
V9oTuOd418QD0U8Ee/BZaXaRNSYV0fzGZ7j1iSeR1XcGc7+vn5+b+D79vP+n3kmdDPsAi12mHRj8
Rn4m/KvT7AE24lm6FFqi8yhw4Vdl4ZhYh7qz723OFt2hTimHuT0Cj6vIkDzQ+8IZP6ZxywNnLcJv
ScnhKeY4LSlISjmb4NcUoWSJ5Ja6agaAZB0vSntQKZ75X6GDTvEexN8wKzGzGkL7hI5IlJBqXZnI
7CY5Yg47WSHJGj+e3Dwb7hGrIcAkSRjLIhA3rxhEopwLQLfWRmWb188oxflFrBzjFoA9iuT7uBTh
UCTbZQhnDmwh1kDFp+vsLfbPJ+aHAhoO5UQHBdj24wy03Ta3bTYzFlfRKmLbulhWFOQghnSfKEVb
EDHEv3MGkM5XwPf+oG0tCs9rbQPpicbtgZ24neIGCI2EhWeMkQlJkgjPAgN64uKgRY2zsiWIifrm
9g00FOM0dnUfYM+kIGKUMC00PTlkLnZr+i+Sm97/PGvTV4z11kfZUd3nXpsmdb4XX6pkjYhGICQ0
ukcTN3A7RCNFG2jIDRLsg2xrnFFnNA2V1i1RlWsQMAQhYb/DMDQRj+syYwPgLwGGEn3QGqinRWxc
l3WImPc57FGHYOTHOVT/TTyM8zUH9O7UtTfKUOi2HcZvvRr1pF1EC2p9bfokqDz2zama3ayeAP53
wpd6K+yzr9yeS07j3ea9rdzudkEE6K7Kyubi/4vN0JGmJcb7uUY/i0UOKxwzaKVBn34wxRVLNqii
SkTfZzLfFEjaOprhtCbkDf1sCuAIzoCWiyvKPD2D1rZ680dfekfC0sUK9rad083Nhd5Xk0/2fdj8
0aCg090auvEWihJecEigID+g604EcMNaX3+tXBWmOXZVoe9s68Z/nX3XKF+uhtoWLSSbdXr9wdKX
G2kUTwHm1ZB0U9NNvUit6HRleU6JcWfh7qlSjSASII2iWTLH76tt41dNh8RxwMSn+gVNsDON98pd
qgoOyNXj2boWg6o4A7FlqR4WcXi8fdoO1N6v8UPYq3xnpO7r6wSCuV55UYzuatskPtBnCPqBuN88
S0yKec5cYX4tcHTVfhqLZ4h+tiF+qSG8mPV0bTxyDuf6EBMRdyYSnZCkQSSJHtSZQVy7Iw4aF1Js
GYB9q87x6W8qumuLlxuw6fO87i41wQeOuemrDW8UXrEE6OWxXqsGbjZaejA0PH6x8b86KoqAcr9c
0N2K3SEaP6flR3/0pl2gCY4+sC8aJ/7GE3aJQKm0jm4Olm1JxDgFcWj2ZAO1RVe+NRbRbSwFKuXr
hlY8gLFmbFl8BHowr6PWLrEOD6699580tBhjWZGR7FvasDszhg2iBnZOmGMaKucJaCzqcIewrBJA
oVCt1XAk4TD39WXteZOB6MEMoYW3xJKMRpWsuCMH9eHD5CFz1fbHJ5hjcixmPQtqoSuJNT9AB0eN
usqhGhhbkZI1QCXxOShxJJFNzkClmRSQaAYf5sBGzRWdEALaZIaPP1ASx3Tc7YhnjGkM5F2sUHTB
c1CekQ+oUb41aeiCQgqlyfDNNVdXu4xDXvvpEjOOcFBiQgoGo19wTWrILLyHjkKyMuX42LXiNPZ8
ydPa//+JopuAK91jNdrdDMTVA+DV0rjQfWOEadrgxVj1SbOhQr5z/NWhLrxegGyD27mxbHugGHrz
MxFVdMWQ5yY9NQ6RP9KSpivz0WePn/DO+criE58J9DpDrwg/K6fDF61xBjocS1/3Bo0ZVh6vrD6C
LK9Z9yxF54P7OTmDRhjxVdzc0xUl/82Z439EV9Sez2W+EMmHWADF6Uc0d20OPzbUuuhscrNduI43
YWNNqkvxzmUszI76aR02Tfuda8S8Bzaky/wc2KN73tYC7GS21IDwhf6+PJrw/XjarxEp0egieuyF
Tmv7F0BWvyzqaFyPkxgUaoC6pQSqbe/F/7VZiytfetreH7pZdhWO8W3+7Fa+JKzCxU3RzKtkl/pU
cKcp0g0HzBQlIE7KSV54BNo+Y5Qzb2ApQAKSPoJUnf0IWIoPC6B1NS1NxS+szYHdNlzyzc/Z3UKk
FGuwIyM18brwI/OSVWOarULcW2aYVjxdKXBKyA6HTlpRAXWD90DfD9dSZ7PvlcDxdiyb7+SZBlZy
8LcLU3/m27BQ7SKV16RxXi5r5jZvgHK6coUbCx2rEMb+aL+2yzOw6o7zAlUx67uaSrnjDmfZQyWi
+gUoVRExRqG6Wa5RGXgMQJJVeK7F2AWbkfUC90HE6cnzN+Nz83IpVmV+j5JYi5KWEAJRp64nNmz4
DQhwjMRrT+OeL4QIAwtnNcVmQt54RI9Kb2STUvI7/gwjXq4qNms0POqsUb1smzNoXKyy8F8Gl16L
8r7tHW3uWqgb+9pcLJpvfbxyHwgnRjODWQSbsCH4VQcasJffl4/7aWcPowpB+WHpIx2uzERynOD5
eJ/FxskSCcIXKx+RiNIxypAz2caMFkekd1ZwlGrYvVnwwTNPFfQOY3dRQ8GWhHLO/EmhKjVahr91
cSfX8rk8uEjOQGPVJjS93BD6pN4s6M5fP5oIOzbsYVNhj0fV2PxeTpXwAgGhzWFPSDh7gVgPEbX8
ZmJD/8uaCzOLeqHf7G5IKdu0yNeZNL7w+TQi+CDYaoZWwxokkwVrkvI58qenV+D4nD8XzQkfptUm
Gnn2qF/JVsV56ZMNXBJHBrqN5zstPTp1yXojSm4IrmU2cctmEW8lBIo5NYIelSavl37V7cqVmRRf
W7NhwCE4NWIuDCP8DUi8iNzGSSRTBGlYoK575NDbPgS6Up76JJhjQfPumxxz5xOi7mIUKcM++0aW
FWvYZ7p+9N2NBe543UWC+/eaMG0PmrzNcBxb2v7eV9x/LeybszxlWSy7p7s9CgR7bcp4+JBIZsTu
n97McfrqWWh5CjEtDNyVPk8XpdTgIWu7t4/1mG2agR8ScDeDJJX3YWnYt8Y4hlUv4RZhS2N/uAxw
IGcB0faPxnc2MOECLUIpNx3wTPIboBGJWVIZ1Lk55zhnNe9xumthD/sHW7s/6rUDQt0Oij3HreaA
1Sa2wlIMc4rmKoIisdhfFpIWcmDgOnCn3q2HfQIqn/iRgTv+rqVvt+joFN4UEGJZWYeyTjvO5jN1
U3JJg4GYqO/2hPcm6KridX2JhAkF7kXg2Vvn7fiszLjbT+JHom5iEXihIyPz2KOOUDLY3esO4WZJ
PEH7qzlaidJoFclKqIazNyyfeHWU2xzEnB1emitdh9HebNXxpNds/+MO6l7sq3Jl66TKIpH0wSOS
ZsZgU95LH2nVYU9pf5oGeu6QGE5Kj3Qsvt0AfKv3GAuPBe/fc8APyPNc2gsrH0qM6St7PgTCNwDy
eT2Gvn03tWNgtt37wq4K/JOdlU9lMpLfo4cY82zNF4MvM22sOqVp+IvmqvjboBH5+EkE4fzhJFti
DIkCNY0OtTBQZdFZA9EaXXl1Ygsgc0rC0+h2fjgHMsVLZMQb4BiQCdpSLHYDSOTs2kIcUHANWT6/
au/MhPgppDHWzYlTq+SY/343DMKkAQQK2EO7V/XStEYp9//L9PFKxeZenv+EZqmwM7+SEGgiEX38
9hbCr5yMW+MkVESPDt5eV1XTQoXPbD7teKJhMCZqWF3+N9dQzv10vxubMgSRIV4jKpSqZYINGHZv
GpCsMz8Wdbd+jzMan6MaSgDlxUDAAML0ufFngZWb6EpWNiq9rKUGPJmsIrdHqVqdjyvz9GWSLVyP
MIEioW03Gtfx8FP8xPWCzVHZVQx9ZKzNocpV+qWI2pieQ73d5jFefHqwkLLlIv6JkpADt9EN/aBy
La9XR0d7IMM0U+vw1afZKnsAISV1+E5RpLxE+Lf4sG986IOQ4lDn0OVuGlwkn0r3+MAWMBKvKcYy
WCflUQ673Si0gWWzMe/LT7ui6rJmp/aPVDq4t4CZpQMTtMJ7cQwM+ITkwZ+SFXB7KDD7HTydmbss
FX3wN7IYTjEIHXOA/G/DmvhH0dpVci+6C5J4lKx+1JM7yriL7iIKgrRgzoc/kYEArgmQKLk9NyAG
JvkvD6aOjz3zPDVoktyFzBRispedffH60aLrb3m0xWWZutoqhndhN4L4wawnrTaWhLLQl77xBX3+
CBag51IPpaR/UsFFdOUR8+J2bQ6AyT28f6UxJCX5bTP5zDRRn319ta8Rv/Cto2n4SEMw8I0PwWV5
l/D2V4rvu+bgWKdbW4gBI/ez0yTi9a5sqO7n3mpy0Qz1sId1TgR/vi46GfstWJ+A+Kf94pnphimI
vzcjIFx8/BOqIW8hAj5szWwPccHRZW6CZbMHqXin32/uxaQeEFJIJjHnv3yriP124rUFnl446p9S
dMatSETXA408YEIzWSFEEVrUKhs06rC0rBnf4mCZerzG2NdRYIH0OJfmp1wfiuXX79kA1bxYgB+0
mN43ObTKyy7w/v5BoEV4GMinwMpnEhwkbu8UtOxTTckU4eFQy/TOm3SLyHpWYMbtrnxpCHRM3ceJ
2/Lm6EBDTPKwU0u1Yo3AlYfh2WCjxtemDoBGxI2uxBQiOKvT+lw8UR2xU6TBK1THqtBxJrPLFePI
JvIkOcRhjSCPIQmqpGwZjN+OvgJh1O7t7r4KPAXYklRxy0YsiyfkFj/lrsirDNMUI33lgm8Te/h9
YSFkhPgSPLsvA3inRYgvQFdSMMxtMFqEtPbP2SSVUwbBVrkclABSTLImgCpcGtaX/TVB8A8pIw3j
LJE0uwF0xhViuZORI4jjNFqeh4+iiyO0KqEJgbu0/F4xCBdSktGW0hLA55ut7xJBo3sEIJ5TizU2
qm5TQjdXqpCP0nJfjMIWKHMpFWUM8jojLHIXy79J1arpNfeaHHc4rO7Aiikr9oNfe05GNAxjAoZ2
hPJ/swGIEkIJYRwf8BI87vKi8FF1j64064Qal5y3DSfi2ykezI8Cp+kZGXHSJ6jsWd+4X8E6yHCd
EN1371JCGh6ehu3EeCbaXKPsvDYV6v5J67ZxBQExEq2ZB74DeLsywOLqJ6FMOnk93C/6PwsBb/x1
qdcYUJYKRdAhBaN/hbB2oS9Q/nMrGaYAWX3py77tSZ75MmVThZ/4+6ZDvI778fMyvxhuoKTqH0we
GUZljfQSPTwHBcfyDO/V5Dv5adSaf1GGex1SgIMy+jF0ePDY9EPfHl5qTKX/A4XxKuAiVadoUVIr
o7RKRrKRrLo7oaRkPD+Non8+eewPbwiGrlfTkUPbrtOjMiurFJY0xVdWsckuQmnhaEvlaftvU2DP
MO9EO5ohyKgWbUX7YeDb1x81aVdrDwIvrfiV9b+XaT78CWViZ+G5cuDa63opOcOCdpOJUHj6SNaw
aY3vdaceaeJm9n+8A3hrIcSljWdG0Hl7l/c1dSpLZ8oszx7DWcyJT8cvnuIpHcf1SRoUH01eowQv
cCh8+OqoqjVyQ5Q4U2mHzXqdbdExKI/joG7HylNq7nEdY32saVBZ4QOCzNUT3awugRl4nYOK+p7X
svaPYGeKTu0q6ZdUzu25Z5gc2MXQp141cdMQL0rc6bizWWXzH1/zKYHoVrbT2fw/pYOcl/lb3+0O
Ue4b4OrWHQa3aCqr2SFeprpcm8hbS9YcS1hX5w+9tsjT3bHmctbzOnTeCToFqg7WVduQ3k5Gpa8m
LLTtBJNUjuuxmylAyYCE8TQALTcN6HMeu/hzez55Z3pRHj+FC/qOyWBAHTC/sVB4yIlFWxN9qEmV
SfTWHscOMioh7O8OvaxLnSpxYIBHdD/I23vdox/f3ouyGmZS2NA+grklV7R3T5E8LnWYnG9jzwIv
MU0r1p7HFK39g5i9fg02F1JHJ77cDx6IRbzPnlBTLI7fDNVMmqv4hDr3XifY87RZYGamn3higds1
zn5CnvsebxDwl0OaYcAB9p3p5QwrvwIkALHSopom0f8wcTC2B2UMNnNv1tqVcrKgHgEKoOvDVgDD
0OcsjIG5tpB9AcSS3RJPIpLkajHsH7RCsuQESBBtVw/YXljDzH0BcBGun3o0EIfAaOZe69OO+rBm
vR3HSIGfDRYrZo2FSzzB9NEGQfTka7MmU9I4vwMYiXOC80R/D1u1V7mTXNIOuaUL0OzAYJgok72g
8qCzgy66j5tXgb7GkH38tvox7kMGkFrsGVmq3HI+dkhkMH2EVtXRIJtmhSEGnMP0y7dN/Qub2sKz
llbXiR0o0LsvIxeBVok1gPyovzNbgu41nn2ca7jh4N55s9XH7vbLVHJ6zxTrNG71aGklN//3AcYX
2TvCxZKxUTHPNIzGWQyOwW+7Ytq24Kz2GA08OlSUMy1DXDTj61QJ3dkbP8IfT9F6RRlvRIaPT5VH
GPmjYtubLlQf1ToQ1Grxe7LhVMgVaENr/Rwop7wK7mqSioGkl5q91U8Qde5sSZZY/87x/MZQr5Gz
GVyV0Cpj8ybbAr2Z7eGSzye/FWoV8l0oDZKFhImc505ZuLoR0pBBn3O4Fly5nWh5Efq/gnDjl4k2
iEp6FJ45n/QRBHR739LHxTjdDKvJQuZx1YyUcEtJwY86jMaRBwbnpw/EvIdTQ9kYhgb2HJIGINDM
jjjzQvuLb+i4EOZBvmC6YfQQJ7nez49tLJx9v7AuRQK34ZvQSNm3KlyknedFpNnWs93XvRcxQAix
sjKcedcm+NMstI7eVrwHG9VTQJsCXQXiGbf/9lDdjSZJ5u0aS8tGSLFfgePmmvIHqF9rn2AZRSPG
yQJ0RqSerIdtUB9NDyU0lPK1tbVQkAhkQ9/LCVtix6YEdMmhnQtqSsTm3Hxq79XoS7qdWzb2XdtW
354K5xyan3++zZmqxIv7qiw/xKJ/fw5sT64/NjSxP87oWWin+q12/umzukLg1RC5sgmnWr4bmHNr
9SuHVQkVnGCuRf+8NheIRVTzWXa/MhMOiJgBHJHJYu66aw9QTVBvExxOk30pJbcLuuZN7etNmzok
TXyhphanWtNAYetvl1RJGfKV/vSrqjYTSO/8ZNVaJp4460hBAZOt2DAO9dMAidbzFSZc6cWi2VUf
pMjv8+m2dSIVtBcvhEMcUK8gdWRZvETtlMzwajgAwNLJY3Q9F+dYVkSTArIzz7Y38YWlGSZETcG3
L8Jyq6MmvMtQeA6LhSJ18iY7c2M8EneUGbgNYMg55XSPGtNl+vTgg/bf6Y3wbjxH1IwbQ7c1Zsxh
2CJ3kJcFtyGTKMadNBQR7d9KPI1qGOxuoWyjXEy6IvlV7kvnddEA0zzHB1eltSdjNDjKP71/9qV/
AEb9IbRDUJzasGxLodLoBU9jf9/0zn5yE1eoUCU36a+qnBrdZRB6qNe67WSSLyrJdAS2ZJh41bs5
vsivNlJX+7lie9NDQiQdIhTD3msCLFrmfxDO0/bcUykpbByepTUdWOMmySdmfENGB7BaC2wIe0lZ
wq0uGy5Q0shRcM7C8it7jojczAKnbtdXwgCC1s8ShLMSTtaACjrTqJ5PKOOYNiJW6iXOfitWAYhS
f1RdBNSWShZBewyikFX5BnerVvSWLY6kxgkC5y5ZQbxcwa/e2ZFgaP7jInZDxCGSEn7WFPHxBUmU
l6k6yY2cXdEIsVdqCyNSF/ouxR4vc5vb0Q0DPRTl/fCoJxypwd50Fk4y1qPck03dhuEF6MtnNU0u
TZP3yQOsSdM6yOz7R4c5w4gSRePout+pVpauBonFIAQoZSST2ZZQ8NcuHJA1UMZgIvzUWlkK4PzJ
KHu8H58seFrn3RUrNRMApEB32wkhgRDpoqj/KgQhSQ8MfhEbK833+b+t8HVo5axLw7I5hhWb9BFa
ADybljuaFy/S/bHQrSJBB497oalDanyu9x2rUaJf71OTbGCaejRZMSN8+ByPUwK8NGGLTpeJylt5
GTIfkIFC1srjS2lovodtLaUXoZA8RdHzciIAZQqUuzrxPa9GkIydxAb1DPZsFmKKiJ8xAr6tj9Lm
LXk0bQMkZRcTb38XEeeNnGot5iW4MSRO+vXTaouQYlv78vUxr67rb1XgYShpQOCrm0fzzu3tuUwj
XtimzaMzxssiOyQsHjMv1mxLms/n6G01DqGD4mo7DMcyiXQCZxlrbhZWeFBTg1EmzEmCY/UAtaay
Kx/rPEq7GfEopCHuK+VfQJA3Wgc0BeT0PGlsdXHMBNt3BpoO1YNYVPknABTkC420qCptYcSAVKAH
K9pcTl6WHwG1SZbkO5IEe8VZoNsW9rcxQHJ8Gh2NrFynLD0/Vuf1Vxvo9Do0TyQMqBjTooHLkKCE
guEbtXe2uDp4xBD6rzvutN46SjusW28PxwnH9EkAZ0hZxDPCedxr4lEem45YmXeToWsnvnRSpKgP
ynLAGWhwgPAG8MtTMCn6O6nJVLwCnMCrlvLWr9wNVImkwTjgBFx3/O5Eagi/KbY5CRNmgGZgOks3
9/fqOWMQclmknkXwdhduFkhlsk+GAoJ9vXhMexV3o/QziaQKrYLdxv3qDUW15uGEMetlTV5rC2Mm
LcKywDXdQMG4XrQ5I2TFxxNEhgf4xzB+8RiRaTcDW6QG4aqh2duMkWO3ISDURFhiAWhH6ZqhRoX7
TgQVANLbcplc78ZeVGnBQGhWVW5rHe5+zbaLBVX0ywYD6iSW4om4p50EXaC91WaMu8Rv2E2+50UO
XeeglW7zyzY7ETa+sMziapePbg95haATVQmdtFRi93wqwXN6P+EocZT09VBnQzjA/QXXPJpFjica
Yu6WKRKE+UrGkxuBkvRa/7EQ9LfEyhs2GACFnqRqkgFBBzGW+rDMT7EqwJmPIM6UuqkSJyW9Tkch
Xr76rKtiUOkM1+URGWOJeGJaVNM/TuhK9SeeXdbiyBh1fW93OalHMkLmBZXqegbtJTHmqISnClZx
+414+TY7LPiBSegvbGQZeEcqwFa/Fg/LUjupnNtfWi8FCFUSMjjibYkpdV41qAV6IIUtbATo4hVb
2e3tSi3T2wrc12iVtD701CE8r+LfuHLzMZ7X+fCOWyRs+mqa8YFZrPihR7jDaDsRe9zWrkPW+f/u
h2C2vISIsYw0K9zfIYPy4Bmi9xjf+AdswVQkEOvMKnFERRVe9EtYeRkAPnx6bjHMf3eRgTvc5Qks
Smxf/Lkx6ttAdxE4TVpi5IE1vuiO3ndpBYwAHU7EWYML8sGpdiIQ4INjuaob6tNtNyWaTB1CHnK2
S7FAUIhQIzTZ/Xag5+ZFJWfmffQalo8koXnSDPfLFsuq7x34n4UX8l0/t+0pw0E81MtJAJloKBm3
3rQw1SPW/ByPcjc2b94JpL8UGRs08KxbuAvgJ8W8un0dxjWObxnaCGCHk8VpD2lW+2wusGvvtRN0
lXq1xHRCoAYDqQMKNuLvFdx+7x3Uz38n5ge9F2regYunIbNRfQwTLJNMNRwOrs0R5lQG8T+7inav
FAKcm4hO119K6qw7hJZekWni379vCXoYydqdesD3IalF4yezUUbUYqOPir5lEGBha+Gr3LlFTOLP
audm0pi3Md3FualsA+kTtqcyFTrO2sFSQJBfjMuAiPj5++iRvuAHP4G9VbwUG4Ds80N9ZdQsH6Uh
Jy2P5Sf1BrEaCwmiL8wwALmkNCaYQqskH5lwZTDelVdaInw8rnnIoxs7Tb2Gf38IK3/LHiReeUR5
X78v79Uueqqz93Eu02oseaenZeZO4Pi/39rRNAHWQ2ASs3dCwe2QF/XRc3iKHWq4/ZsaRFZIRrr+
IcVLma/J3LMs7AviUD6Gr3dY0C8qDK1psYofhEFhYS32owCiiB1drlLHKoj3JobYoi0L+IX9KxLA
uVEqD1QffOr9/iqtUYyx5ri4fQ39TZcStSNhsNnv4PQVikZUYCqdoHdn/5cGDoP+39wKUWWhKQFu
YE9WoQRdpcl2ytfvu54kUiryG+hd7GbBtQkEoc4rSetcXeTgUXIqENpnET9UFGmOD0amayukVoAK
hxq6Bcs8Kx+QBa6Amx7yiMzsoR2FM+5x3W2wRf7zZVE1rDSP7Ss6zTwZpZ09XAblGDrm/gjv8icp
xm2uYc8KRXnvwvIB3ydsJTw3i4noEKVjew76GTJfbl5u5dWfo2NBISgYw8ESJRUJpku2LChTuIbm
zwaaBGHbmJfImPLnU7d+GotTDm596/Z6oxymy8yqqZkfKcJe8rgOkmt0VjMS020JZON19KvfbCkN
mFYBOHMBeB09E2RYGEdb3ZWBsCDJhBL9xfVx1M3NGYBrpcXwmwc/hoB8EiqiF5LFBQojsxWAOYxU
d2JvlzBR2YSNil39P1VIoVkDLYGCcWyV83ZSNVs5PDsPP8Qd59ZoXn1kxzf8qXXkEy9A2b9NWjum
TLTuGLaqLJod/lH3WiYqPFkg9UW2Bsz88s7bHOsOtbIgJI2IOwMw8Tr4zb3eodUKCSZakMvZL2q7
+DrwIPVOMbEjXT6Lj6t6wPetJ/em6RwmfxIqxtQlcQPF4PgeAX8eEW9vFy5dwe/NQHTxbTboMNIg
gPHU9hPRr1GwAEVPQdQ1TT9K7/Cnd//3Nu/fDS8sOdUs8XPjeYF/Yo3++Teat+SBNfnpOpJcv3xp
ZXIkJqXUsTZzp8/is9ciNuKva9+QbRkxP5MUnnYyCcdeMPInnUWdcl96bQIgTF3Kw27tG4VyhGpN
6okPm3XTSAftijXMSekHiCzTeMJdHDf9FZAtuUXGmreAh5w7ogM/F3HwDMMilvrtk0pfguutyJMO
bZHNg6JYHiaBxW6Q9z5A8KVc3J78PAtOjEA1OuL/44SH0SaL6yrf7AnKvrHSvN3rrZx1IJT0Uy8l
WFgfuOAWqMZwL1NPLeiq14R7JINy/JAfapdLMFaMRFIp487+ryeDvn9owurnZHFuRtoBPq9SDBtk
x/YkxUqKqlZAmvqjFIrjMAN25+lHGnaGIdjDSFLMejIriJEOUX2xpUzo0FQaRiMXG1KuKm0MKAmx
TixNQvOEfJBnGHvM38hc4mQKc3eDiDNMkGlVom4IrVvgp1X13HaUhskieT2iecyTWoEIH3WO/Ct5
39nau2LjgkB3EIU9tONIOw11Z8UMRUMlvSOW2LE9NYMJA5WjGliI7UgDxIHDkLn1iISkwDAZ/PBt
28sZFSDvjc9KAvaBihU3fvxZgZ51CPEsHhbxPexQ4oe56ekyLwNAVWFBzsE9nlRskZYtPpskeCpe
jtkuaj+1mTrfkt7+MvCcZj2XqU9FRvBIX4U9LSAY6n6kRJUEQ2jSkCKn4dgv040NfXHIFBLygYkJ
wCE0s2zamFByubGZcJLBmwxYg5Y2uWW/4z3DAPTvbtkdxFS6wiGaBVR4FqB7vgmLifTeI/BX81xm
ykj0kJ46AmR0gN1cXLxZfRKyOo2QUlbu1zVAcDN+LxJhU7rAV+sSI5jyvrFUKyqEnZrz9vwFy1F/
1kapKtsw4cVNUmS9q21O6Iu0OD+RaGePMnGQNBliSaUMXZR1hm8mhVd/8EfoVkF992mxUXh6p0nC
u+0Xb4PEMBLY6X/Jup3yAkvi4OanqrLRbK6vhRaCIbzcDr5jYbvoeCFL2oOb9zYo9kC/4cLS75RO
cfMZ+9TYfrWcGY5e1yWpUkdM2KEFnNXR1wF2tQy9Tic4B9eRB2J6ryFl3oD+NxhcT/C52FyMWtme
ybgG6JARK5zYzihNDxy4ALDy6F9ihs4KE52KKWKG3+IgC/XmqrN1YrchZ3bHP46E3GWGWFXix9in
vZqvi+Z5QFm7Le0NT6iU4irTd11ibiNDaZlvgiF0aCThuOF+hkXqLmsNMM85RpaZt0EV8I7ogfm1
qPga9YEWu03/vDIvJ9eHDVz5VSEKlcT0sufPeRnt0zRspFppZo4SYFjWMLAbea+Yw7V3g8riW8rE
LPaoi1Sh6eI+QKHezRJIKPlO3Xl865iEWb211hOX6taF39kcf4muWieev/jdyoHhGW1flN/bWLif
illmDt9btdpuzkZwG3BLd6vapOl9PWsf8nBUhFsvuIX1trkkvB9MdjmBCp4v1wnD0FcZUPkFNVnN
33q3QnQ8dsiAoby8VMFQeUMfpk9UkqcT+2naBZpvrJ09+oR2m42zN4mRleCAhJ9Aa2NKuDkMYgHk
1dROmKm5J/ktWuZwPLItfWFEQGqYv8eTTQQPPqdRd7RupBzVQea+ctEJlKidjLI422HhagHjH162
jefmNby4N33Rpxp7HV1cNn2nR6dnMjHTO77KNbE9BNJn/yK6xbe7uwxd2PKQNsZ8foOBK2KGajdP
NDJFWDrlMtQtZraGtNHoxfDB2JUDOEQgjLiPoP2Q2t7+vDFRn5HxhA+4VDL8fR2UNj1niZLnb0MW
WqR6p4K75bIJvQKc9xt2wG31L91uGk0R8BXsOy2RJJjxyA4UE0bUWoLrGY7IkzOJmVkw5Sw1a235
2cQYDQ9XnHOjpTrjWGyEbEy9nWfbgLt0Rbm7Vbdg/DfSBBCcO3hC8ZaaJ5xmztQjGOauHZuVwW05
YQEw3U8x5NE673LO8aYc62ELQLBKT6qdv4LnqaJnYE1h1DT8NTBWawBPI96ssKYoWRASAqgTyI0C
t0LPXjaKwo9nyT3b42waHsueW5FnSAYFJfneH+5Oke/+TnwwjCSm6oYQKdrZs0KeDYwX1r4mseSV
x1h6LGdJTD9QgimriPuBWvGH1m8jq5h4F5eAzNpJinoElZP7rslZ+knAPvBkSoe/a7HXWLH/72UB
HmnMBMMz9wNxDe40+j+kqsJ5yQKGrPZB1CePvtCHNa60I56STlGzAZvK+ZxC4KudEFAns+uJgzN/
foUhTRNoB90U+AQfknB/Uhk9H7v0u+NtgpjYpBEuXWgsyURHz71+eOQwSaL13MFhHjB7oM4jS53J
dKJCFY/AH/eP8GWGA1pe81Z6D3tpbRIl7pVC1K6P2LbYIPbkZ0qo2htJrHBB5pQd3YeSHUd2NPGA
dGdIoBCK+DQSeSlI+PLYTrGQP/5U/qcjKXcJJcDA+ARRWcqUHBg4qMznu5wH0eMXm8mHoO7TsrcO
k13aXkn24k1Xqm8gGIBGYMbs2vJ7pOWEQUq8LyVEvwuIllYCoxe3jvOQz1adZzB7JMJx0ckpJXbn
JdlZLSTMeciAE1bGxGXdlgaQbGR7z/kjr0BQmBEGYefeYHC9S7hZ7zMjoPEB+BWpzWkc4PAlFw5F
RTMbD5oJSggg96LUA2Uc73q0fmSJjgph33eeLT9fqjrjD3cMlIgeHwwmy2u33zDm9YRQjSVJndmR
n8G2Az5IgCAa+hg6pdVfymrz8t4xDVo+yWWM3XiOUHqziPLYhzYfJZbSqr7u7IBBoVeqxoEhNP1c
O3CVg7oYVvo+JjJiI/gZXNeEPRCuXRfjn6vhtz18a0JLptfcDddFAvIFTQ4E5VukDew6GVNfG/Ty
qIsOzWDi99LC+QPI+s1hD3rW1WmNyNwS7qUlLWixCiRPkorN/4UDbBTPNmvSSGfiBWdZJqXqTOlY
fAYx649s08ImxbAV31ucuEotCFY2lysBP5zyJhKuZkLKZ/7j0mJEXOpIq790r8A1n0KTi6c4/eGr
+MOdonBd3agk+DwUA/z83jBJFp5DJwF0LybElWP5fLFOaRmYqXYrHZMc99z/9XhGW9s9Q6UUU+eb
zmyfMn4WRarMlxK70Sf/apXq84fecHYOOK+rChkXgx/eeGAsaw6NLAY3bQ0Yufe91XgfLxqaOaSA
ViYyTP5hpk8WTDtCP3ONrFntrhsNeXxOGIv2GAoN8p5o5V1fmnb3TUfV3fEvtq7MOHma5Y9qiwfX
atxDUD85qXCdIkus53gIGYMdeCzuMjYSoixwjThN4mztID5iLLiELW4EU7hKz59b5o1IRRpDsdpW
d9NJ27vnhm2gIezl3Z8qLslwLEbxEpEeD8ijnRDbyVYECcgbG7RCFYahiEmV3mxO0+WBTX/X5m72
gw6QobAEkkQz0QM8VPF897VixYlt7F+hO9SOEXu2H+SwQfJILtP8MWv3AU12yA8Rd08ZfdEVqeBU
B2Cpxu0OXzHjZsKBEZ/BbqbGGCCPYRRVIl4tfkRrsoVV4zBHEt6oSbCwxUiak1nI5oPI6tyoabdx
i2ynsNw4m9rvYxrDCTb0I1pZpD1BRKoZKYsUoYlf03czb+vWz+OvzNJEpQi4Chs0husyrboSURbC
7DkE6KmgSBR5yypjOwmY5mqv6bWQl5hRRQhR+4FaRVsQ9WBvVSsqjytkvqboKSfN9NE8U+Y+XH/s
qlS0PG1TRyc+QoUO0Lvi7J06y72jyhbiICZ+Uh/ifo5qzWJgrlU2H7rsGH8Jo6VEAy90yQ+QSqmA
V4tIx4VBjvhC21QTPhU8Fb3xIYj0+tUFhBghB8Ts2TnqQ8rlX7A7bS7FUQLribni6j3LZ90iu0Y+
kd37JCvpzmMU5VUMtR9U4QbOJlGx6prf+GJoWKADbWJejymgZFEWqiieKKdM81LuQ2hBGBdPvkwO
SXcQn1zgTxdPE354qvIz2z0AZJ90SgIHKuDIs+JyxQlABx3jEj2UizFWpsdEYuIfcP2id7QKHDbO
NLSkJAIiAbrrojC7GQ4azODxEkxA4S9cFpukolxvk7gxrXSYD8yQEfktlYs86k1Ozm5RTsQlo8jD
z9YClcSyPswBTT8BmJtKAWxD8IE5tr3f8A8UBZK+vx3cjRlOqrEXWmZfSDEl9oqS/MszPWsAxS/h
x/XoS2AL7LDMTtcWB63AfHx6zyP5V9bdyesrhBrzDCxYkaVPfpvWLi91TtFLeEQS4dND9tUFWE3u
Uej9sqa/7hQyxP4RbfT3vsQ6SKcVlJLGndD8FDcy/6cif4hzXL3QonXXo6TW1KAl5ewkKIs6lSez
ECEqJBY8kOhe5hChjq9xNPV/kPoi9iacdsmzgQxL3OA0jJc9gEOPUqDslLenVQ4ER1N1rZStpQwS
WqNh1JYsw/D6BReTvOnKQVestaRRORX4pBdEtwS1dwIffow3PO0VyIB0Ga7O7IX/LPUqbvR6m3/6
zfOj0iS1U/FWffETe5sw/5Y3KOw46BdCDUZQ8lNG0ZmgE0rrM7N3qu4EXO+Il2+VOMlSm4gKvjrA
nP24xUA341pyLm+5M6xgb8V3zfq3DeW/cj3BuPSg2HzkFQKLT6zrrK2Kn1mo2LBGZIHrtgLDX4z0
wKtNwDFd8VsVivEMQfngiP6p67JO9oUyUwNQjbnvfNaakPTc8UjuvQUkRvHCEEUGASqGPPkXsCQT
usE6xC9hQHj0JlNwcTai98AJB/fRehgEOkq5vE+In962/62DAKvPGsPjOvlCrGDqWfRkIGiqVfRu
zBFma3I9QaYZuI54a2F/LQQGu4u34gJCxa0sCnnsqfJzgl+j5EKWjoj5LWmP/9F5vE7EqHC+y3MF
GnX7/uH3Y0ZR5oSRVcz2RdlhRMV/MFwdrv3fOrOj22e9w/o1Hl5WpvrXGf+r4+VgmQ4Hhmcla7Cm
mQrHjZfDsWEVvpkMnO0qZqGW1/UYTdcxjPVUSyfSntrNegpCSkYyxl6iIK7XVzQpkCeywK6k+rEf
AC6PZv+mIT1x2wWfx8kN+R4Cgxa47UghovTn4o611mukWrpnhyCedsVYkx6KHzICoaeUt1CgcegW
SDrshCnwpLnfgXNAwIUc6a345SudrGHXMks4au9yXgBLyz1qZ6H7XR5IVQvE7RUvO3ulV+l6jlVT
gL6FMjX+4KsL/90+05mLiovWs++Nnfb5iyFZGRe5yEylPHg2zpR3QFV9h6BSp7C4brwDqCPQFS/P
d4N9zZ1U7H6pUalIgpUGk75ry+ehvIpGewdYt4yT7g27CZR+IJoyqJq1GVkTHerbFOZMpLeg/PMp
9adG0K02jwTtzgzOr8+zcXeyxTqRJ6IaMn1uMwB4ZP+hEndwkeSK2op2QKx4sr7hdEYIgSBJlqtc
oqDrPKsNiUDMnUaA0q/C5puiW3cEQvNQpZ0F8vaCUUIubum/cmGlqKfCIGSfBOtDcFuuZ9jye7qX
k/sbJvEuHd/SKOC9mgunQj47Q67LfLIc/DVsraVyJtZ/I+Hdpzs1Lsz7Yf7jHes8iueSIHN3FcYO
OMRHlvrf/pRRoi0qFFDdBcFn+7lzbh61lrwzA3LPKX95DKF2u5O3oweFyU3yhSNRCnje+ugI0oxv
fb1VcktPNPeTfKRfI52TNBzKg8C5mh/8W9YC8O9WYP2uv8MDA4gZW7I0jD7d7YsmriQBNXXsDEFh
4sCh3YU3Cm4mzEWrNDscOqFwpbbod3i1CJ1rq3u7fz7TinX52tQO7qfpCeffFWWupt/Bfj0o1vYn
wNC8UiC7OQGaJ1TrEN4gGsm61eCv/F5HVNAqjsh4JSudC8ZV6BQgh2eImWeOzZXKpM/hmekZkaXf
VGZYHG5wDyV8NJNyTtpIoxulasGvouAFsvDlD2qtF88XADDQCu+DXXl+3pRD5o5zvoJTGtgjZG7Z
gHKYI/E4gYi2LMvDF47NjVYkAdTdRETLX2MrSFEwr4O0AHpQjH9SBR8fdZbXblsm40SRG53UucHy
xIRh8Maiws9p9loTUBRxMzjmGDUlCXX2Jdd7kpvRTbr6Nhx75NcCVfgdvQlSNLw1qVSIUEc8qTEH
p7E3T/u5isoBSx7uCPqujYNbR43q1cQhhd0p/abv2rbF9vnEGJ2w9k7VMDiDeaLo/Upitfe83CuV
96VTHjI86eC8eic4HTDHXrP7TuwuZ4SC5MoIH1ue6gDgmNYMlrFRB5cszk5malauVjjc87M09Ilt
I4eWfIi7FrZZB4Om8siaHQniLINSERGABVoLuOvwO5Ymttn9MPZX6SOZWd3p/Qch1Tt7aqvBM/pP
pUIAbmRYC+3M0KeyfLTKrnO29fBBFsX49o6CFomPMteHCIxtZxv9HvzIGUN6QO7bC66NzB92TYkM
WRCJ6DOKRL7BIzqTtMYwN1T5Cx1IK1uPw0dsbeI3eEAOuGxxYFlzTAm9IvUJaMK6l5dKDJRjFYKI
zMV8NyeWo9mRqbG3BIP81AbwW7YEu3NcnjvxvUCpMzrLJxZFqB1FGV/Cnf1IdZrO4Z515HaQzd5c
FB9UVkTBAu5BT/pos8AVjSY8hhXgKPVQZpabOIovjEEzQFbf7rmpZjgq4jZduaJqrNq0SfCcneCs
FTg54kgDpfzRy5T1nGWwtvX/oILSyk9ZoMfgCF/EiqvLxzZYiDrXBaevgKBpdDV+IEGsbNyw+suJ
4W6pgXdDeJE87cZrH0fCMuieFtL/GF51lckoYZZfCHovO6Skt3ckkJQ1ts+g4uF9wgTkwzj+dQpg
yCUYgIwQJ/shNsuwxU9vdtjRCvSa9clEa5W08hM4gPYgRh3FNIYtCme55nemRNtbfnZy2ecDb9Pf
1mYd+UHXd/aey8w2i9xq9UKa6RwBcAFSyt9L1IuUo4KQRoRPAwrMvozfy1leJRy9MlDigDuqnkG5
LUtcpuyAW7srEwnYgogQ0iMZ5ckCtEWslDcAdVTEMpV8A72Exrvr2rEWpqQy31ISi9+kdN6lkipT
OYBSjAAUHBtBpIoCBbDwedVPsDJvzsWtJ91dbLEb384TgFsg4wTCobwv2AwB/+NcDKWRWJmGukUr
MpOfcnHYaPtGFd4UtYs3rsd30OYL1R3o3hXdBGDdVq3Xz55UywMEt6zPo+EyhYJog0egj5/MJLpK
FN0W6jDPgoRozYkNcX3F0SsU1ybWwlg3A/xc+bVkNCxApccDEEiTtI702Cl9/p1jpEFV52a2jPme
s+dhO/cMi4WP7dbpCYT0tRhFlj4pyLjPidERRzFY15AhW6HRhe08d2U8+LvDGSmZbDbedlyiDgDZ
eWFBVFS1oDKigMVuy3F0dA9e0sazrxaL7FI18v4TSKXPyS8G8NIbSWvPIhbpVWHzC5Vk7Q2hbV/F
vrJQkHzSrUibUTkFHMckd6+YWS062MPa2pS1AZOw6zAIDA7dJpxtHGAo3PzrdkNjEOGAS1R4PRfq
nGNo1iGZVHp41wn8a9ymukc99i2S/7xRaML5DZWizvyo3c3EdUKp3R1sHYCYcxNIEvr8usywonR2
I7V0K8NaZCrFBDUJo/WAjZwUuneIsidDHZGJj9OfRTUMetz6Tb5H5AwD5SdQKwFrLfzFYY1Gmfrc
Ugb3+OdOmfNfUzrh5/5JFsjQmot2hFp7j3DrBsGv2M4V6E+5fNgRAuyr7KvuGHERg/OOUFyiXA45
ghl9Wrodj6RLKCRIkjDRFoELPP2+eHCkTKGj2dkwlO4RkwFfqjESJflk3rByDbTDxHRTEmYMX6Ax
clv9QtRr933fp5T7Hs5dXanyu5ROrnKWLwVyaMcK+G1n/NaWIzk4rAUz0P806v4hYNGY3PU7aJAR
/jyz1mMKBzly50KSrVY5m08DyIpz/VI16gM5FpqVX3efdCUKycGeEEIc7/WrutapFM1t7YUQdYmG
c9z/xlTKQN66mODxOJOczbN5f6jfGeUp+MYXck4TSYxajl/MN2GgnjwotGGxrqsSpeQ8ZVG31ikP
Fdo20qxuwpyNALfhzGTnns0N7KTEUA3t8N5f3vZdyNXCy3ZbpTGs0WPfNFqrertq+IsOtqsh/GMg
zO+1HJJ2vWIziioAslPk9oWINEOQow2RDrQI4zekrUmgHOpBpQVno3cqlCYUX3CNlvD5AFdzu7wJ
IShJYNYupe6GxAWPZWfRPZ9yv6+SoncIHiUfeAKlFvefYbW3aVOGXEyuchCDOTUeYwdCgIj0O5VI
hHZxMDpw2do1cGTgCTPY+ADdiMXU+WJXYUPEKYePMUN+e5mzYynsFK3WY3qSS7+iagZcUuIibwri
tSZ6PV81WUSP6CY3li2qYYTiXBrjHodlDawTl5zLPgAfg6exEPMfcVyJja1rtI0ssx9BU7P191a3
dmVgFM2bPNWi+++kDRoqE0aLzwjlS1rC5iwWrwIlPTfmOimaoeo5fGFxoENNEbij44iDZX567jS1
asNUN4Z66OFHrMJ+XcrA962giQbSTyLuCpAPdwm9FFE4+sPjnfL0k6WZ7irJHv3jWinYe4o2aJZ9
QeR40Gu6C9OQBmfG1kcw/fBOjpAMAAtXKLECneshF7RGpQEPJOCtLVateO+zHE3fmayaj7YJaElN
GSWp6m4dVyVwHEjabyAnArDqbwDK8yH/8aCd0+rndBWCH1Zmoawy2lud/Hnq4Gg/tXSkNbVzNq1z
Bbh2C7zxWUiF7R7qCtmMsNuZwXUQqhAqtv9OSNE7kC3vzQWXGA2fN05mK98oRZQFeX2HQa60oDle
UhjHEChupX/0oUpTztp4OHXD7kmsREnceZvCKDGCqcRRb2calnxYwR4daghcfXWxpMwvHqcH6ZQp
EnrElpCxsgtI/+Ngvih1jXH+Ml1lClPdCaJ6exBzkFkDSLv3mV1QG1LEpXDeIAJUxoLlf1iT9cl9
DnlvDxTxe8cE9DZ3+S1pnCPEx4NosktE0HlcmlbVALMlvd/aT7XJAykpZsy/3ZQlJp6vxRh9Jcts
jS7/9xzxXiSUxXUKpN0UQdf60L317ZT0TrO8zGnhwDvtdthZE+LKoyM7P3snUi9Y05nzOGh+JRH/
/Kwe48vI24+zCFMUlcx8yEpQvj61RIlMfu5czsZ0M2jMTe/DTi78G/oVF4bfzK7FWEHtLgA7ghox
64unr1LFTj8nXgpy1RzgVO3KncrQrlGUFxRrZ/DZpguQabcfg9lYzEaR7ewEkcSYRm8Q2PnXE9JV
dnIbcBZMGK9vVFLbHm6mgKPyj5NNCTRIObyZby+zjfYIpxcdDV5LEQcNREdu33FSNj4cD35IUydS
ycmZ1KYH7WrFx0OaxajZMJem3M9naTZ17B/qtSFJ/X9EjJmQoNOoX4jqsZ+V1tXv8HWcD35nsP8/
3OY7vLdCFU/7s558C+dwr+Q+cazzb71Srlysf7kcOXwLDqMJ7YbbLwNVT4sJKZK4DjD9vHQubYMl
HZDgnH0JnLf/SxohI6R2C1kP047BiV7UkAUORqJFcIrS3QvQpwNmschZH0Xxt4HAM1Dm4Psbns43
trxHKe9f0+r/0l2SDKR0F60NL4AqDoXMrOW6jcd7k7aj5xSiYTeDju6bEqJNM0bL+It2g2LZhy1g
jzK0GZQeXF2UJYPIutcTEzm8ls1hJ9QM4VrWScbBsV9cGWVP7xQAcrSUkb+ehs393oKovOQUFIid
M+UzlHEkSQ5nKyFadOBhonsKd2hWIvszdEFlekUJQG9peD0hNGIgJXB98bdSG7LGr2U+By/uJ6pS
CnEB3P1ydnHe2EOmLlQAcwz/6yi7lWvDk87nN7saTRDxG+jDvtJRH9hBH4Yme9th3iOILQlJCFs4
RjSVao7Uxm+TCU4XwkmzxThJCi6E5Ry0yt96KRQbn7Krn29laoFIuQqZkPza4agKvhRhxGsjkHeV
tF11CaDYXg64xUCwB46nG2rwPZg1tRe7x9YKluogUXj1k5Yca3WYz41QI8TfyDIirYR6Lo99GvEE
ON74e5AhlNVGLjadfy3foRkxrY0NzuHtUnRftuWjDpIMc0puDsVKJEbHk9rkGxqUnEzZWD26jd9X
j4VdfqvlHykO1WTk3SmHiGFT175INc5DhtIE6WuhSOKz/o8PsglhczZ++/FtOgbrmI3kdz119qo1
ivOAPlw/M+M6loWkl4NBoZJbXjiy41l6C0GNoxSEifuBkIEV3eEVmSKOJvfHFPrY7gSTNyoNwFqb
TO6JLdEgPJX0PrvB1z3IR7gBp+0oib3/n7GYQKgTC0iR+IqB/uOoFqfF3OzZ+kllPXOf3dKZbcUY
bhPwca3kQ/0Lb/+s5gjMm2KwBklbMUmUI4vSlh5Filv3mfBSQQNP9Rc8QQVSlFl4Gm+feXvwWzmA
g0Vczs+WFeeGcUO+EguELTJ48PSiKIuZSzLatzwOb5qTq4EpVC2qJJSIW8526Cr97OjSrVRNUtMI
Kin815jjQ5qOna04VQutjiGzyQfxiP3H3yQhoViKEqrGwhlhY4oXiJcNbpk2YigYLB3NMVllHR1+
TyA5fwWIQzbE+AyRTJL5SXeCDA8w1wGbILoeDzKoFuxRsRsYewCFNEz8mRb9DfEtQwJtNCZFgsFQ
CPSZS7YdtZ5E5WJpFBgeK1bJz1hqdMpzN00X262CvvC8uz8Ot8IH6FzLdtw2qKyEs9/Ja7ZkLcEd
hZaHGLkEgpJDFtslrmAzxXl4wT/F/Rt1O56mQATZ5zcRfGPafOOOcIFTVbaBaLWNcxTSB9yWTsKz
09bSRdPsbnhERZapm6DGttM98m/bHhCY/Vf36pM0sIffczlnaMORQrmwSaqcJNr3MQXWJdtHeWiH
pYYCapWdpzAo3fNDz49a9MsymqesndnhjcFZ8+nw7uubfNLWeWGyuDLcARxfS+1frXoPNDOCUd6r
22vq9PGPyG5qIlQqQh/iEB7YfBsE9KjNnqfQXeuXiyUtcLhmtDHYkNglzXG4jfcIe6bPe8PAWolT
oN9w81SRIYlV/CMO5eiFEiSmKZtZyjvkaQ8tddCjhnaKOQrfTMI4qWWmU18WhUTacAHtC2A9hIaT
KXrPUvdhRNmMaHRO4ZP+iHECfAglHXDFEtri5vzoZ5eLj0b1TKfNBlOfXYyuKDE3nyMor8o+ZJfo
8utH8itWO3yV/1PopKREYJW68+KqJaPd0/SpcVgSkJP/KzfOK0pNGMjDGi8O7Y03sV9q87ts0Q2z
Tfj04McUSFhjcpPvwPrHHxaFjsTePF1wRF13kGg2cu0jpdQ99A/QiEHdYnag+BPPpHM77DRZ6vZ9
L7mKH5ycCu51f5tYS+Cw8sL1hh2YT1CEmLbZrTJ6BDei+IZ4uFRvnkBqJohwD5RMyLo3kVhYaAG3
w+WX2hwn7nfjLPXJmuE8OM1gC4SaJ2YjkGMNy5P36BclhiSpI33RNXuE0NGq2P8Wilnq6JQClY8d
9CBv0aM3wHgOy5EGMBuQ2QRbd/5U7JIWlSBk0tv+R2TfuqHz19OEg36iCkaAH2YtZtGDhFp1nyv2
B3snbvN3xpug+4eOZh8eShvoySJDDCLaqH84CDxDJc9Lmw3XnXckk/CKPvb8zqvpG6472AWWp9pI
lC1d+ewOD2PgG1W5+ewZW2ZxSyxZ2MqbDCQMmCDzwFNvAsutlp0gVxgpcszd9pgGSn5gUUmmJ9py
VUOc5wsOpvgZLxRwOIweoxGFWrCzUzFyYKHt0pkMLy4vB6ctSGerpyAVvazCoiEe43pPXpLbv5OQ
0eWQaki5yz5md92bkWsCnLGDJLZESBLI37wY/rCqsQi3erDKWZVOCO/2cQVKM120fH1lZWV2invk
UU8/Ar6m5maps+MBqbKd2DrZMdEf26q78PblcwIZrkYt0eMvfFrTQi47mAQMZZC72OaNxPtJfcEA
/kWXEbRABtfEjgBUYX7BANsVW40SaOzLn1ElFQAmFfW2SIOLN52LrTZqypYQjLw4637cV1ULFl+I
hKfc7MlMdGF97B4fdlYmrXoF23pNC6Q53flgldJeMKs9Rsz0BbVDCaQDNzT/TE9tVce1LOosAW3x
trWBtDaJdwpRCgxaAN64QJyKXmdC3l6CqW+NH9h1JTJe0rlTGezs6azWO8TShILrkbkIlpcPDRlM
SNa6tR5G2wHX/EbGRkjHYhAYvgxq4tUOJocNGHCUMyAX8wG2d53I3/WhXqD4NA5kYQv8NYQNtk0G
oAkkkQHUrPU4i6Lzoe+edOKONITqz53oVWh/L8BsrTVYpGqcZmMA4GqWgSAm4XXPYnmdfw5Z9S5a
DRHSjCS1uQYFApP3LuR/t/dWV/1PY3FNwbbdUX9iwI7uu5EtX5knej6KfXKBcnItPenJUiEFWROQ
tZ8K9uXiqeaXyKF0Tx4dqy7MNdPp2LuX1cg4KOI/gmT7YsiQMmrLuCr7bkrA/1lzEjmrF1lPeLi+
n9cxt9NJQXWIaUJ3kEiWOudXWiS5taMslA6u7zcz5bDySNwbgxJAlKP5d3Gn9K/0y16OXExIaayf
idxJruDEnVBxH8zEioyOGZ/9mpztLq6lPbfqaAKArznbxaSW260yusGtBp2UZKFgIJKYVOMeNdnu
Rk3ZaFjxYxU5b+jDZwZ6DlM0AH0UIT+cA97CORXaK+yNwRhVf0sJPPecrlgKzC8uoyNtMZPxqRlJ
PJBoSAZFVcm8yJQ4Vuce9aEWvZfSmf2naCVhmqWov2LrZqjsvSc+ucwAUSuPDOt5gnPt14RyJbAW
jp3OWRyZKvh9gOFREldVjHS1+vGOqWovn9+QBQDEnHbnWMuvRztYWFrP3z+/vnxHbBUZODrLHe/K
lu/RoEhM78r7tkitk2DMzQ6h7ZaSP+rZH2qOTsWVVNr+LhUzivhgStzeBrFVfwKRc8qtIH/84uSI
Jrrv09W3/oMpUXpCJa8gjVi/TiGiy7towok6dyfgQamj+CQPVr/eSLZXldpa+AGW5oWw3+FhaEPQ
MO2OYG/0GIC18LStMarorbiik11kZpUl/k02Qs3xZ3djWX6Nge2wzqYuyJxs7eo7E1dMqgz437Tm
KMSSXDNtIuGunU7L3WDbvp5IN4WFZc8kYpSOjFZuT0/GtS1FGL8IPz5D/UONxdUc4gRelyZUibwh
k+8mM291ubvwIvriT+o/Xh6EOzG7QgFd4CnG26orw7P/HySz/R3EvL53B3tpG1+Gvtu+jPFfStgI
xADBjvxf77PzW135cFzoNwEi5oZayenvZxskfpkh1oaNYkrNYyPR5VEh7m79Lxuz+XaJSHDdsT4Y
VEYjkn288S5hPUUkreLx02wtzYalAKHAQuWWq0mSQIpZcqSr3WiXD/auIVUcY2p8WEM8HaGHl3LW
kflXUDe84rjVAC8OsM+ggJJENlQVGvl5v0grFOwl/xJKSTPGDHCBWTQIqcreusHnjLiRgRn5ETQ/
oyhukqwzsPvH/vxkCPJ5I1XJL/HeIpAIFsTjQgekj8jWbu7f7bX2UilvpSURJfAtYEprj4daxylv
e1JUX3zo3y9WyWd0JQ8r69vmxCoNRF4k/DmKDYDzczRruxPHNeiuvHdP2CDV1Nf08R3vBD17MBgY
4N16FjKrcJbji+vDCJEp2x1EhcCJyVXwtaS6K+J5m9iWzGIUb0tLZZruLaOFbvuxvQ1Ni8i37xm9
kDnn6AvthMKvWUmpV/vDkpkhu3IqHnB0X4rZ4WvaZhHtlKhj3qAIPEd5nLf47cv0SzJygDsDIdcx
+nwHXvy/yXELZy1mEUQ1ou2rCiDzWiyowZ3HQCuQXcAFIBdgBCN4CjzZGjy3Gz3wPGRTKL3GFMgr
yX6NNLUYyOyh0Y+wuk3ngY9gvsry0TEDEPvV1YFMKnhvdZ4yzxweWl53WdN80Duj3ElkYh/YuAFZ
g511hMhT01aMx+WChmfUlnJmeA7pVln6doUWSbWRsIavmonGxSj7jSPzO0DMYB+i2OzKu0WpUojL
JZ5duCIOhe0qx/y+kujRcRIc1khtM6qyMhiVcJCWOrzg34Y91CbzuKhRGfpNjVEfXjtXt6w0fKun
xYCsMZMEaJ9dcFsP56F18zLavrjTdbdlOIhDhubWyJE0Mw30e5x6ioJHbE2iS9CB/3LV7GjLCY9z
rZG8434zRAsI+1UXt9qis9uq9cPGSBXwgXAhHA1SPn9lBipUJCL7zDqKe1LAhXWWMILDgOkBPDwe
lbG8psF3IooWhM+xTA8tSo5mYhMelxtGOWLqzNmvX9inMSHvAdf+h0lg2VeVbCMWtJBpFCUD9zi/
gbqGqmyrwNW3NjUiXAfiKudDcv9U/GbtFlLXFevxdikSDkqJPmkYG7UkzVJTwIRRpV9NuaMbzsG9
qB+Tsga2FeIwGPnKuZRR9D/eSW03EyIbhsv6AS3y6qmWJhnh7pKu2uqSrkrxJELBIyKG9taeCfK1
ywE/nHNc9jkhTb0KZZU8EzvzuBVfF/d7RP3lcUbAZxDTAd2MZc+qcUG8dfjkDoszE0k7Tq1CEK2I
cLKEIEaFQxgqohzXLszc3s+Kzna4rN2fK3sRCJDu9Q4xvydwNFHpAMnvXLQeo1w4P4dWGGbVG9xR
wgKlGZGuMWrl5Ja2Nw8IgGupUBNrR4KeMIjgGveWATouAGhb0pmstNAjiELM4Izgh6R/hlIOhsYM
nVsO01e0kpwJaR394nfLewHvyrHiXYe0SzHG9sppnTOksMLzab+O7t+vExVkdVko47et/e23JjNX
Q9UPDpnNiWoAJ5eex6qIVFgiwqNikVIKiomGqgzabVnXhUjf+nrEsyY20G5FJSdNP6V3AY7ZzuCs
1P/chaJHKsSxtBe3sFLa1Hjr8YpksDYeKNyXHcvIvrRPIH6QEY0/uiAkAvwu9+d5LMdLtrYonTxN
XmH00T0tE/qjyATFwqv523KkQDlG6zKNsq/JCp8G0cN74oVLCUNTJ2QXCww+/pD1h4Hd9ywW+Tzb
D+ZT4aLbyD6WTFiHub8UAe8DvInNsYlgCkyBhQsvZ7vnVn57xNlAjOcF39LZrdif2SIAduwGg3lz
0espdwNnRuU7akhbuPG/2TT0iU18YMLsJUX8XWA2SvBaQmaeRxOYHEcLyQfsqHtOPJ8KFaltcNp9
RckgoUAKd8naLQfWN8hyv1MAfuaa/KGv8nyOKSSBSlvx6sjdYDprPrEwMuXxkSmGsAKlwvAVKKSV
TBo4C0UOU9RBYTQ/P4z/Vdv/jpoSt2qIJ4gTUtV828jcfT4wfJjZWoEulYr1d5IspA/ja3T7SDgN
KYr9Gm8IbdcetHLaiZAhNkXWQC0/EgPs4sU4sdFF0UKVS0KqS6NO5fmp1Uw/Xgq+kW6sFe3yeKtU
ic9S3Pr1FionUJVCrk5GBBYquvWWNdIchDOh8IdMbTg0TdJtsyrXj+TNw7w3I0PePGZf63XL+pUj
BJMrk9x1rj5XoImiKS541ElVcpNOGJ+OH09amOr8lXTnse0zLm4JnCR2e5g/rgh1G+bBukRBQVfd
keu837ei0FRqwe9v/cJ+KFnE4+scjqnaJFe9tyY1J/cfH6inaH5tSYkCjcH/V7op9BkUFCzRoMTa
MrqtSxgJ8c6EeeCt4lhZGLWg6jq2KhOXl1QIU9yH+hdRnFTNbSyAqSreDfXbESnyzFswpXBD2bWL
rGDTUAiIhlmbHARTOtlatH08nVjGaNrPh2PgGb6t550iw1U7w/ThAw6kk+2MgK8lTKwMcahx69+m
74EFIHQch37+XrvRoGnCmfkiUrsvNB2AZtnP9be2v4KgXSh+mAte5/fb9PwPcXo3lowgOhOLoe6P
Iuat5gidMRVUT51pZpeMO76Ysvv7BYCCq0cF/fCZgt3u2qHtJ/q1LIHhs2sOqQ9CVYbyRjxmzcm/
I+AIPsDAaUrbqtzLau9oMOXSISDl8ySQKfBNs/qgq6RCy9JMINr+6b0KJVhMqXCzmp0NvU9Pf05K
ASR6haXXyTHBB03RHIEdAHimaZFcDRlh5ItYmW4KDiRalvn7P7FMkisRXI7CpU3f2jjO1VNw6n2T
UJINXaK34j5g8wYxaJ30DAH3/nwLLhmzRLALj3CTnMzMRRMoWTV1+r+1FesJWlWtRkdqTRXj0TIV
CXkN6SE+sty1X+cmwOlowZagxQ4TbcAX629xhEG4psc7NJng6G2U1iji7q6N65HcKSMnpspL4CSf
nhaiJmThqXV9/Duulo17yAU3qqg1STPCY1NvpFUe/DgY4nJkVqUMIsI5lF2dFNOYuQ7mJZh+9o8U
0frLJw6x1CXENN8AxfGFUtceZ26YFxQ9cU5zyWlHbgTAxkMJnoXAzCWdyGEctKiTypXhnINSHKQb
BuPevemwMFzgcYClNB+hP9D3Dxd5PsB/ymos5IX26ud0gEPi21C0LE+uYYVsV+BCkzaMRpP1G7Ni
V9pJ0+IqRiORMcsSD5HAIBjF5Sh91yCjAk1f6YY4SnrfNKOvyMhfIEN46Ir7ydDhStO27ZKT+xxU
a5MQzPaWn/Ek4o7Q03KDVs8DXzrJ4GBCvZbSkyWTBHAWqM2SFWIU9B03LU2ezmvJm71jn2Z4BPFv
oqMPV3Pfn91KQ4cc1YcAmvh8bhMkzpZyPx+NWzAAkwyHqL00jIuWKFZc7dpGu/m4+C05zH3FgnvU
f08U7msc8BrF8Qo/RoIu+PJWvwXklkfvgGLkEjMgd9wwrVJ3rqMTlWL6oHeVEBK2nAY9ABCsoUS2
YrMFkhNh2GDuTE8CSeiuBVKp3//a8RPZzGBzEj5C6W0SCiHPVDy3ncndXYCMMotYbSdxFRhx/w93
0xnT97YrXWEXsd7Ja9hf0Gp16doR2P0T6IfbEP+QfUzstdgSQKbCAInKVls73f8Z8lwLQYeQza6y
kN21YywKNxuemAJJ8JGITZa5x1W93Iph7of3DUbr7ufxSgOKMkQ1OBC2PM/5JOPZi0iuhokwTfgM
tb8vLEtzWZRlkZeea6z1+LoGLVYDFXlkTdloIN5VGdLAPwllZJSdz3VTp7ChSJP3jBDWBUel6BUL
U3A2rOra5zQ+LpT32rhjnJVxWuHiezf7N7bGk2IwSBPm+u1mqwpim8YvWki22OXAP+e0Es7RtMGJ
nXA7bVJi+IXcIOftURKrE11irBi8W5JSV1c9YZsmeKQpa1GVZI+36QshO6HsSDQtYQ4RyxpsGgfU
KY0o47VxRPmIZenfwbUTqa9V90amXGIyIERiAIOzLhD+/qCds57B5z7uAWxvRjthT0dK9iHUczAX
d7IIOIeOJ5mwmGML5shD5Aijw0b63Gu1IMQhGELYjHQHYwuFlFeNGaQWmxTn6k/MbC4uwwZmZJcN
l5p2/srseSE0MZrpCb7OE35ZRHNJH96uIpceEEO9UAh/Cw0cu3hc1fOOjKUZaMiEe5rF6SQvqshy
/Sttl/4WWywg7lA4VD2KjkMZT3DvM+FYxVml0S6AbcNanlJE7X0e46/ZmcCxtvoLHQyvYPLZl3XK
mOMh5bd2xV0PYzshL8jrD7yg0S+CX1Mj70iw+UP2YAZdIKb9/wFb+5HRr4rVzMBCieitOTa2M5R+
TFjYh4xfD9sxbcO1t/rwAqNLFuP9fsg3qKYHKfvNEyFJQyQpxERT8uiAID6bjM9CH271asXz+9o/
p+979GJXqmrvR98P+00ztQa3QdjrtWfbJfBhZP89nOduQnAT0gKYrUG5xKmzt6ooOVSgq5pSnems
sIPGzGdc3c2mF0XB3jhPmsRFOWzJPbMQUUAj2vjO9Y8nrYMRkkQTCGOb9klA5qRXZazd8ql3/N8K
VQUz+WhVee239wQ5RJlCO285rmfKNV4ryxbSPsSGqTXtK3cUcp1BhcpIoZKcbKMaE3/mmn0sQ3HM
I870swW4o5V7fpnA2M+Hta2bItoeIQ5ssEXvwGDDLxe0PYg45KD8278bckpxrdZeXjQD9lmQrhAT
Cra5J/tBMdQDgSXWsbwCZevALrQ4WoMb0PPjyfT9BB/7Ej8sM4e2R9sU50vZtRedBYduWpPD0DE6
TFMgkVscZEWQAQgPuL6j+F5hN+chAbc8imMqXc4mcW1pxvE8P6Lk92NALL5StgyouhlRhX2r/+Es
uQI7ViZl4dQMR4WrO+7LiYje60SfNO6y+UcgziHgfSWJ9Vgd6OzlaYtAqShrPPe2jSeDCWoOcZ+1
2S+fG9k0uJk5p0usEYRDQWA7jqCxBZeq24qkJALvAj8E70r5sh6NXpaq3nQCnGhWHWCVzi9nGTVB
mjkebQcLAt3CSzHkicFjuuLp0DlH2fbw4RBdWl1CV4UHG542B7KTUU4594Zal15DuBuStcRshsBf
ObQX8fHBizYNWGFAdEtUoei8Z8g0B6L3bwKrVUi61V1CIocNjEbJXfsI+6OUWGfDZt3o44QTEPHa
Cte20KTcv+HVwkafj46Oi0P+MVqJtOmczI8lwmt4JaWvrtadN+qGwnKDYfE/8P8+8k11Sz+6oU2Y
zSHpUdkAp1rbbDGBbB9dl9DMTa0r2r/tNSI4PbD9ysnScDJqVxsuJzJxlNF7FxpaH9pHftyBz0pB
AsDrJsuaVgAz/9SWWOy0YYljWW7AAy1UfyfacJHwlRWhtmcuCGlGB7KVdZVzhcy8ZqoMhiUlwVqi
dtKJz9NUC2/z2vLBD2G5Te+cZTqAXnAQmcTQW4VWcslkJSi+TMZRk7zWol2MBQNjXbqWW8NhzVfO
N1PRpPbTXRXk3JywmU3OvnhuljALqPO5wtqzakrqI0sMIzbJlS5ywgsuPx0AylO3FhMF3NRMsueW
GBcdLoipgJhtssly25/aGWN6p/tbiwkxo0NQeU0CJlNBT2tZQIxE/sBtEt3qKxisSA/CRpLhyTK5
nivFk4phu1AZdrP9Fnj7Fsf2znqRZ6APlNFxR8AjzVI6Y++zh/9C1zuJ61U7tqTGsEYDrF3DxnlC
LRor2bnxwfmAVDkABsgXxKTdrhCt5qwnItj3EGiCw/qpjEAvQhWSg7RfIoOIrWm5ldXQr73nI1ff
c210nQ45hJaOeTgoQe7Tgu5uUXClNFAxHzNEc+5koIZoHMy23qBD7fIu+fs/jvexkuq2DzF61p5f
O5Dy266vejItGgL1OvSZDrImd0n+BBVV9RmlR/op2L7x564AOJ+NBl8VMGXkwdbh6kpk4MV87AAm
e47HRemjL6CyOq0ZECjHqdwYKbxH7NrnEixizkyGR816PT2VvVOwvzs0UNRM/+o1JJCHTUJai2tX
ZKKB5njvLIYk2xDlkPLzOCE9ebCcrtRveVc/ogVNcOZjuke13fBD2xYXr+EPtXm086GqYuaBrekb
b0eH3vyB+l10NJzmeXVhFsNEwVYrHGUYSp7XU1n4o0j/eq3/Td25lqIfmcoPdG55gfx+985NtnI8
0tz2WuPyAf2oQUV7m1yC7bZnsa3koUukezt+/zxcnjSnpR2ZvYaTvl+B1CQw0sWaVM/BX9HyizL5
yFb2jcgvvTk0MdJvTq0aQZ8w+zgF8lBBSwsBS9iarVx25dDU4nTyatVriaiKRn+1KIPLOm52+FdR
2ZaML92w3Cy2jJvE6iXpNl5t8RVn/DEUmFlg/jDmQ+nvyFqb0UzNTiXXz8a8pqmxmK+GRKte12T+
Vk90XmzubV0djp1uXNSD2ZQdMbtLiVXOsIevr9uwkqyVi/ot8kSKMcdMZXr8+6tQTZzifYjaAnuV
HxNWYdXKnzx67qEQvvC0GxVygfueoT5/l3iQyiM9w4OawH8w0FoGRrLre/AQVTfMPZpXxh4lz/bR
L9vC4qgjh3pyGG+zBSiTb5V9GV+Tw8RM2xnLAbmDBUyBCfTGFFJTVtZA2tloWWz3Ma53YRlp+z5i
fwDRaKNNx7auHc2HfCabGbwrJZxTPVHT7H1bmxbF73W919lc0B9VLqCRI6NEMqD1mm3mXcLcNinY
zYQUMEhhFbTNjWPipipgVIg6zyx6SwJKJw0ZDbGHIxraLH0YtlZlZ5i0DivBxpm8EpUIddDNyrvJ
qb9eqhrhejuaRS+8sWpzIi2JzwLbloQOoogZEFLa/FwiMMKeGExVoGWekV/NgQ6FXa46fMzY9ir3
xeSZCBxwGstbK7QXXfG/OGjM3cf2pJpaNs34LnCxrok6Ztzs3PiXuUWFOu0Fh8GRc8CmYetm5eWo
TqUPq83QX1U8+TunAaznA6EVKClCqMjDMX2kNeOnHgcnDSlBmsOrIeq8LVimO0L+FjDKGzQK9ghR
U/O5EFKwe+pa3WSv3g7Txz53NLyub+cqpfUB0idatvg3JEymD0XeTiU0JdKY63pg/W+mikz2cmZX
hhNldj2TqvzYFWeKwitQ1xbhKrmjxYYv+LNnc3RkVt3ZZJM7r6/xUqPNon71F7exH3UdwWgH/lZ0
sU7ur6i52W3tJdqstqKfBwUQBfw7MJZ8wORtbu9Z11EgfbGbhQbbMCZu9+yeOCozOYfbHnOqU+hh
vYeQ9Qc+Fz9O4DbPwnsjrR2C/5SXxdvBUb9gbsCiTp7/mF0fX1YE8wrskx93ObhejkBXE7iI9Hti
PnwSTbN9cUmcJZqvQZpxhs4c2RRAYkKrP23I/UkExnsObzM7U8rw5HePvTQh0ho15gubWymsOqZl
D5hAWL133MViif+YGrkYYoJdtkbh0PIam/cwW4DDb5nEBP+rwWAnUHjWsfiU+0T6AupBBkKQL7RP
AaT0xKLBSqq8vN3WBDQi/FtY4cs7mPcjOUqyvsa8vJ1VkioOtNVG8slotMfY60hTDCF94mQr/3KM
SpJklKh/hV93k1OYBgFpAeFt5RwPi3CzgDo9ZeKs6zLbe3/BuQnYK7CIKxjeeqcWzp9OnrWBAbZT
OAq3WS0YZN7mCD3XK+WLEXxZrso3Ew0Wr19yR43xaBPe5w3F3k1S123/IPVG9MKBrcpru7sSKkLB
XX3Zj8bSri5oQrHVN0FdPd9CFQNocPAAi95nxTCadUnQHWtUq5lH2YQlgrlGtesZq2a+rPKQL+No
FaIY9Zgo6ge0OGM9DjtfizufnM/Ppuce3f3ORuS7U9FqC6PaaU9kUNrLb3juVZRyj7fZrBQ59gyi
TItex6cwRSr6NR+9hpBbVs3zma6RQ3fU7HuV7385klULt9XJmXkvXr6zwzoDcgMSsIr+94TT5m/c
Oo87VDM/4HZkio56JfAnitgaeG6AzFO1aWukdJ7pp3nh9swA8YAD4ZF+F4kGb+pQFih3EtAZUo6F
do3Smb3EZ8JuZvbZu9O0cJc1/a5osdOUlUWbVAEWoOCxq5X9NrPywBpuXspHn0JV/sVTaIbmOKGz
IzHphVQmpxwQQEStEpppFm0thN/99FmeyU5C6mTOi5Ay0ajwgMdN02Q/CaLZZ4e2umRc4R4BF+HF
br3VGEGSvxRwqiaYPgkgwq/yS9kG6APKH/q1VXg4HvwXda+QFrMN/X5PDGMMy2eS7mRddXHbXsm3
4KTlC8qbdibphax0eC3O4YT9Ly1FM2bHpugRWWYKYEe9lkygUAVjSp2L7nVLQ3jWgkicGIPR89eq
N1iubOOy5ZtgH7Cb6jmgHfPqUrzyf6F68Otm01O4jELse6VppJw/ulOMnxJwg3RUVmnXHgwhvz0p
4CQ6uDj0Ui3Vcz7UGHesqZWdJabZuXI2bEcktsQ3723kuUmDdE3UGXAON7U2sH69HjXqUMy2hRmB
xPwniNUSYeIWznYuqzwuwnSSA0E6brAfppP2H6O4gkuk2FP/3O5iM+EFd18E0C3bq68kPtvyf6zf
7WadyAXIbsjCOMAsE6HyFo9L+8Ue/9M1GT0VUveYq4Eqyiv2h2chP74KT7MisuCU1osW9kX+Z7fE
/cbmW+NLNH2PB5rJwjCtsKyA57rab5jXqLsHZANi0paX9bCcNNdaAdu1KGqJLP7kPorSy7I15ld6
X427DsXjU94ELbsU1pNDXijI8uHBdiy0999Qu3WQDmqczvE3C4J9/mRd5jkwXgNJdksKnQzzITpK
flTfldqDqnL6bEXG9D6nDT940sg+GVAxm5hUqOX2MQpRUdX0EPBn8TJHKRJTcIN5LWAAEj/92rjM
M0Wgv/psktAjyMBFhmdSbwPI0XHTboT/g6KHsr62XhTE2dbfG2oEwJ/vaUMOhMkWORYWsZm1vy9T
NYce1H+INNA6+1U1oYXFvfZYCG1csJWrnOUUYI0JTqxg0H/o9ytAF2zvAKAEviSAOLBb/V/OdtB8
I6hFmyxVuAG9+lHwmjhRHh0hwmDzvjSa21TaC1pOAPa9s5dSIcqo63tQ371zS4zOnwbLlhY340tO
ryPhtE3cxkj3ifuGpjvpeeqtjQa7/IdVebARV2FU0ipbslP3Qo45kULdXRrlhlTf4ATdt0Ac4HgH
ZMQuqchSAJi30tx7rZ8uBtU7wkW4+pN++DN+ipR1sSf4Wegitm2zw2HdefnEOstkf8xVNZwGvH++
lgl4guFHg9RWTghInY8UZjrbZC9ApuDh/ApTF+DsbQsSFzFb5bG9y3zguDrCeupBA18Lk6DJnH2b
ih8WVGD61M3Yh6VCWqOiySS7z7fTwOWFbpVAr05yjIJkD6FxveHUghxu5hPlezHOiabGJCVW3Bef
LWEH5hgKyQI0ZWlqk//lXgk5Licaxhkh2pycYAFlfZD+Yy7Ca9TX05Ccb8kL/aTT0FxWEH65e6ff
1NN6X55r1yeHotxvM9QHaO/QVvoMK3PfuV5zXo4qDLiw8k+rTo7BrB/3vahPS43fJ0voing8Qk8N
aYpzYpJK+CSaPy4vKWV1TiHiX1i6h2uTMK/JgAFdS11EExyiXDouJez8q8VLk8JSzqt0wD1ZV0T2
cL5gYOvb2U+tIXlL8f5OcgFl9RxK7Pm/7HrcpLyR0KQ1Zyt92C3YMrhxlZSmoujbfKWzmj2p0ivV
auc3HJt6sGUqihAbR/6zKvT1KzQp908WvQmqIeJ89MsVWrY5GVvxnBtefjNpOTEMFNaK/0UBnbf9
hZhu2Mf40c6UtGcdON12bSoosf5D1yKfCOBtpUCqcGsrjVpEzv9tdfk6RmR6LR2zMw+Yo1bxkHaK
bIGtlg4Qtvhe+0auvWbtjhcELNql1kmXtVK5aY3bxwkIn7YnqQU9eL3cO3VGYNuMLnJ0WLHI8JEk
csNTWFpikKSJjw237hPTH1As2GoOaEaZtUQEFZEmky9oL31hdJ9+vdgzT+Dbsn2W1p+fSSI65nhF
oGkxnvRRUBeRzCiNrBLvxG++gccSBO+wtJqV7ZbIuVU0+Sp6M5e6Lgkp8O+o+9RiZMNWxdnosz3m
HuIjF56RboY6ISh2y62wxwP8EgF0MC3kXBzXXOpmC6Xp0OCUpG4EMi9emiNBASN0N3rr+DB5A4/d
ErTktY6vK4NxNGe7ZBg5Y/WcCc98EkbF+znM3qJyQjtxjcTd9ogHdCrZvhY87C+ntMXVmaF/5PWp
tGHVnJ6kOoSkThSJIc63lJ9vG41nMMKSPja8qMgSPrzTGmJGCeO9x8VkURAwk9cIGUCJi2xUTrSM
wf4GPnYTsI6bZXskHiiKYjx5UXfVQ5DWD5WD0/W/ILwpcCo67PGfH5S61P7vVeZKrIwHpru3uXXn
9jT9VjYOyhaLfnmX7+okkeVXXa1MaxQQStVep69R8WLoFiqtWz0yNxTYqtENRFfEdGJAvQOX9kGm
nGHI3pqqiJTXZPxbh5cC/TJCW5l6oCvclOGkuxU8fvDX3hO+mO7Za1K/KwsvvyGHDQdbOQs7gziD
9LXJWXn8QKIWdExtlQI/KLgBbzvtfJXdJWtzcOcpj7YpTX8cHSBmZMVh0y/UKe8m/QhImOzUwofa
ufGN38xsKyQGwVGA7SxDBPx8GAW+BFeC2fHJw9b6gFKw8wxbG8GOP4pFGrZ05GfR9Tvf5MV/YMHq
J0e1l3gGI/CKhSnRnlSKufJ1F4xBMoMUSZzAFA7cWAOOUBxxGOnaopgqLbbpwo0MR3ET+4BHRYQJ
vRp1vqmHnDv/UtVODjX6829jxlyUsPYFE0iio2uubYXtxffw4NbiQoqudKJ+k2Y1RivkLFBVdFB8
hPJlzmz8QiMVkrutB/BD6oTczmk+oOa1afXXx+YWz/5/HoP+ku7fd2JOBrUFS0hLnwm1+ToqAbB4
FS7vTJGy6KSijwxkJ61PIAbiegSosaZPal52b7rbE1HJnImMwpsV1rxDT5qKRzKF1wDSpmNb/sPG
PMbtP2KaBhErqswbfETRT8GvUAXgybQ3SDLCTwHzOLmFRIZOI8bHLTHUpPqeG3cbuGm5HRBK778y
fH1sHFswivE2R4cpQ1qeOBfK7+IPPzeMBPHM4uh7DgblqHw3R6SLrpgFWfk+ruZ//xG8aY+dAf0y
3OZT8CUESoxW3Qp4Ej94i/FyTvOjeKsF+5uONuNe/45I5Oiz4HesAjDlEFaGtt8CDxhcqWO4DIS+
S/PFpKQXTSOd1b0RLT9GPYSf4SPtLm7l81aw0u2YxRQN+B5W9aWskkUHU2m6NkkiWDxpxGrcntyl
de20fkpe6Th/5zd2/LTSRSg8/KnBi4UOdtEqgQXq2Ntv7QhzTg2d+PoHJsNlDzpSgCAFSv+QySeO
sZpJOZvrUlPjipmp9EswYwr19wN2ZtoQ12HzjONB1U1Q2D3+y9A61qDBMyDINQOiEuu0O6AyLYt/
M9b8ckhB47ERLuef3Mw4e/PleqjkahQDkT/iguxHYtIO9Q0v7GlFk2DkRKf7hLWlnY3rY8wS4bWh
abLvsChOnlI9XFcQ3XcL+IO7UHOnrrxomgr50TkGH85NuhPpEaY6MuUb/ifPeqfpZVWnTxya3kT+
anuBbApFXT234XUZoJyOaLzF8UW7Jb8p1IsgaRbW69M+3s7WyyPoK74YF1Z51VkrueAvanxeznn3
LNjFyDNx7fpCtzLbD232FhH7AgID4xSpBrGNzBsvBT7L8r32ECYYh4iRklOByj8hTW7WJagAcKGe
EifViPC4o0bVumusjE8VVyeVNye3s2wfUlwu0pM953cEJg6kPTjBJIDR4yeOrxLqZtGJ54icSDTj
yQGJ+qbOi9wZ5C+xdhdkf7jqHvN0udOKOeGa5DSVZcWsvvCQtWsZX4kHJ+w3cR/k6Im2eU805iEj
eZ/VGVmH34Uhks4tnUQXf1wN2laj1yGEsNCb5sf9XD5f8BhuUFM4cKKWvnpUpGt/aInpVpn5ugEP
HPUYG5q60tHTABchivHjaHaKFFKDSoMWhAfuEGC9eZ1iV5c3f5Jkpf7CAAJ4AdGrh+rYMaEpRoEJ
JnWHbYhDEUWOZ8QZ8+tmTBQBWN6+qwUsLeXpGIuR8m58IjuKponNNlfHY71V9yFIYpqsQSLwqMgs
pNU7laS/9EhyFwN56m/KmXpmyC2DCcQFqu5YFjS3ZKTjVlGDA4HBCCV23muUwMUNmufA3qFZDELL
Mnnijam/EbZtVRRxw4AzGRwT6u8oUllJBT/uoiUw0qJCC4tb+DwhvHGR+2DTa37/zWD1rLyrCX5X
jFPou6EgCCWEWOVc9G5zHFoVlJMX6eSNoJsA8bPTy82gHLw9k/njFIoh9hF54Sn1waXz57AMWX5y
z5l/+NsazQRoommjIxfWA8WfufIYO4jL674VsiT9R9ByWpXoyhs0vsTb3O8DCdbp7+2qTcjKpWvo
GbezlPc3vXlNmMJ0/vCA43bUiLszpiAl00uCvhyrNkfi928NkXfTQip6UX3sSmK965b8Tx3+lBtb
baQ+vl4OjFHiirKyAaV7NkWSONT0fE6WyPp6YSS+QoVp/m3r1QQyH3WWPIDKON3IQP94JbXN9CZh
djAgUOD45Ek8BdLgSllVnujoh/ajTHd/jYLOAGwBn185ymZ4Y4lNGvK07d8gIl7a4uXe8ym5F1ZV
XPfQdSCTCt0ZypZ43Nka8+8EgwKMB9p1MXUz+zB/MZsUFtmJDIj0YYGyXmpcTOswLaRzIe8kb+Dd
BiOMSPT79kuz5GIVVwUPjICBlnnQfvLj4fMAL2LZci6ZfVgmrBkQFJhFte9Np0/hQnJwpvWbhRlb
oj/0rzsLOoXpAb5yu4xIeQ2/Uax2D8EgBpNsY5d/WhN5I+nMPHpnsn2ndJ9ktJjAisipgcMeMSMB
iGtsYpQZbS2yPevNtIKZ39my5GHDJWVVBNNokXfrq+NAcbxVRQW6Au+70toaVXMxnUY0Egzi1h8c
CxIjO4vO/BOarv1BGiZgcAdCrPwIx5SNZ8s4a10MTxhIfVrwuG314S6DrIa8h1Ot3spgfSBa1kVk
2iuVm1WHLwnqhqVfbPNjhb4fmGHE1kxm2iw1Qc1Bq80f+94kiWWrwoegFmJUgKgHy60XdiRrZEaC
blBWx67Tn1HxwiGUH2ThArnzprHhwq2kvw/g/c3HcG77qHsVq0Gs7CB0CU0tWor/XnV86iU0pDZN
8WsXNdfqEV/UeOxre8dFtt3DEGHF2+Qs93p8bjzuqxaDePQkAJC5FR5ICw5pTQuYEqzvs+Kn1UyT
kN37c7C1Z+oJdgtLO2kW8pPnoTRZO03Tz8SJzt82rcJZ0WwHdlUphgTax5tIx3eSSsVk4tX5KQwX
/BDTK8J7aeSjudf8EDsaZISZa7T6T7O9uc5XBjRHY0lPBKWZF4CjcC9SOYhQVTkr+qArpuiZxxqT
vqfVAjyIwS9OwrhjPpuK+tZcf7NtDlBZpGNgSM7UCIxWA9zouz+Hj0sf5torxnVLtE/VetGw90Kh
wGcjIaYdlnOOXDS+PRtL7rfi4ip0z0qUeV1GfoEWxPvtg7JDmZO2ZJ1atRvYrKnpl6ID7bk2ETAC
JLiCPyGNhrN3usXsKFvEEupl2Sr7gX5dLIwpmLBiFTwIoxfBhttiC1cjGWwlQqWzZCmG/QvD4A4B
3Xqjuf+EdA0IZ17sEXVB/tqkD5lTtB2y0UV7hAlWHnwbuiUXphgs0/uSx6bd7djoyXbebeah97yu
+vfnAWcFmH4wK3yUmjsO6SaCoEI0cpIYIO4QKzuM486Ac93VbhhUnGyDH245wACrH3rQXH86fVVa
bpCEbrglRrnBXBVUXnU6eXET46SOO2rI3XHxQ5skRQzgEKqqj+oDnEU1tAuZ+9069IqmEnuh+3uI
UnyER8iVfo0jGR8EXGvr3AuhN9DrRGHYIXkTaJxw+q00Fy1MmxqdC9gZ+StktGYEiJQZ1HiWzFyj
BmOB8fKrswMNpykDvQfwDvzUJOrgh5Pa774V0GxYV3gNuFzWpLEVQNGDb2sglbIWodI6rEj+yYoX
k9cYkjP4wn205B81jdy0FIlRfrvKJRHJuZoDyPNdlMRKLj8KKUd4AlzHl1WJfcx/3KoNpMyMp77A
8ZyloRM1eyLdp7rn9uh74oQCEP4TczvLCEuUYCDjFVI7kOh0GXbDMqjwZ4Fwse36IaaA4XhPpw3u
vBpVwIcr/cRosa+2/3iuIaes4G3Z8GdJ1HuysAy1st4LkRW6SRJqHFl/xTihOmOeNVQI1rq5d7fZ
S9Y4wWuCoO4f+N7Oc6tmw+xUUUvWu2vGSAMqylFLUrhk9GhEPb1xqCisf/fxNvScdAMYdclFQiMr
BfBJBzGhDJxKVo1qXvYZ/f5OngjEMnnfSDcsU6nqtjg/n6P0uGa2wer7TjPni+ekmPagW9khfl4g
9inE2ijRsconxB6TUvDiXRbhSXkPlOOQgg4CjnkovTH76NugnC73J506aN2EwN/IdQVid/xZgksV
Cnz2OUu05xLI22GRB7lEbrupED1bNKD9QVYVwPfYBqC1RfDjG40PCQcQtoHA16FGHWKayxbMGWJo
kmQFIckwlsjRWJqsWrYr2Nis2UL8Y02IE9pC+rQbLDug2u0SHNGv/kkawpX6U6FklD6s8aX1L68v
Ltu3Z+OM6oSohN0MArehDBbUuA5RRWK8SL1CQa3V3QwBl/AmmuflyYs1PfyJ9Gy05atKx9aMVvhz
41TVrxfqWgLRPDp5gx9YkZgGmoKIofTV3jEXBvpJz1pNi9O2HoT4xrmzTKw6oTbbmzbaaJDJ4sDF
JEXZRpSNQ/TWTZVlMkWRFMVIaZxEUT/fVlupZBlfBz11D9DGc5RJQ3tR+4uahUUHTh+4hPLUcok/
TNthVYIsFYFw42X6oqN1T2J3IOxasM/qU1935/mk/JyfAaa0ZdtBZHYOkIXSiKwAJ/NXs6UAEvtf
1H+iY8390uC5HPefedIa8ITJnQmpTUJK1jD+Ay1w8RQx+IChmxXI3d0VUNJFqD9RtieeHMI5xiEQ
ma6/P4C6KpNX/IkIU4uiNiu3+PHDw1ZPRbQhZUqJ+cZanNTy6YT6yySk6dhIQnHTtYi0tjsJNSBh
Lc4V7IAlHAO8yt+eilPd0j2qed34fTcQy5gdGNWsxq4/i+Ay85Ya3kYhaOg8c8I6yVTbPnrl+0Mw
9O4KQt2hLFKEznAg0SwdhvkC5aJAjH696r/v66AXGJWWdHtwf6yzUUtsOHULLyEkyBOu4TS3p8V+
TGOKKF9KDPQv3Xcf+vitT77FIWTpwqh0Nz5edUQ4kd/pCYKHKdXPuJOXjIJjy/byz5pgP1pcPHLt
3ozvB6yJvGC5j0Ms4Ex0zm46r+Oo73hkWvS5GMvGFeFki8K8ZqWun+C4smyFa5oAQ5cr7irjUacr
WdIFPefY13JWRmE1oH/4yjVEQSPzjwu4HkKk01/6bnAwluGzuDOcBKBi+0fdQ1IrKbIghmSyNQmi
tYWtMyM95bwGgC5HGKEwAXMln+sWFY8OUGoUmAWms2mpYJWP0rI2cOln7ffJUGtSANjfs8LQr/zH
8/geGDV9seSx2rChoRfSfYzyQIFFSBJXw+1408r28bh9GxUqP1we0ybx0X7fifvNG9KcfCDvEqRY
zQ4WnCuZTruVjgltSAEuWX4qP0Ec7BsJW3kJUHi1RG97XCFiSneuJfJvfbJBHwzIsaQ7eZ7zu8gu
2lVE+Ox5MVWk3TE1yPSdYGD063SjMdAs3knUksRBhEJjsJE+IgMJ7eoBNeuJwia1oVF3vUFtU4Lp
GL0tCSFwojh6fW+VuFadrGNA9pWaW19j7tRw7P/PwQLQOZ6sSOM5JXCpDbCGBqJW39AvyTdks7xt
F+OWbreV/UJjdo1VnmohFY7BE9eiLyzvJyO+s9wbLj4pMbN+sEPW3VJsJFceANnI4+LGtYT2btYV
jhUXSA8irVGlzEYgDsc+rN8Wr29wiqULPbgJWjz9Y1IOSd5r8RougUzTz5P6xbW6DSosyRx4kqlh
tCDuomsn4xcc3HOKlULzuWw1/sdgD3yra2FZjNKBjN9re1+0ujfGwMkzw9DFcFKV/h83PQbiym9h
NsTl1nfEgLiRQZ8cLq4jDqsZsBYdVeLvhp6WUhEVaHN6bGSpjeEKV7/Drs9jgyRDysvxCEnPxyAO
isi1PcVgL+E+CFSP/e5dbKxxylHHHRGZrGbK111/WSBOpucCgrX+r+EIcvRcGrJPMetoXY0O/ZiC
X1eGVApg1MRmioYkzkPf98pAmyc3NgAvopJtZ1UWPc+k7m0AnbhNS37BHcNjTINWA2QpucmleFp8
0OjOyryBk9k+tVOSjxKpYPRJaTJIaCfTxKml8eGu/xv3PgR93Z8jBzcazlxhDPPBci0k8Cu+8kpJ
wkndjZ1L2j22uxaGPKZxLfvcffpUz62ST/tVqv45Ka+PHpzNvDghNr/9n059saE7lW7VgS3lHoia
IW41nUjs29DDu/XFbHETJEBYNE7pdfdMlFXwnA8bkqOdQJR4h+E1yDw7MZRnfM5YB7aTcGVwaALg
8ZLbMkeLu1ewvVwAbIYRt7KD1gfYcaR8zn82HYbtCeZK6EOGBQu5he/pgokRy+9IomDBb6MeHPuc
zFWiKhvfD9/NbRrLIMvjHgkZpkKqTmd+2fQyjdIFWSLCuQCg14z5lS1LX0yo/sgiPZAqudXzobTc
9w/c0lluMaUpDnY2DwsXEwhL6vc0sXccb4Yb4Mng3c+1wYunjpV/4dja8FmCmw6QkoAMsUOs8Jaj
QusYEcObDemuSwraItDjw+57DlOifEuNI6o9UVfuDQfzGkjk4Ldhd8g9WmE2uBNXfe7s3h9AVHVl
LGGcWSq/x/pM1THj2wXFTlhffZpZnEDwTcKhuiokKfQNNJtxUGY1wbd33Pp5Jo2DleXu3IgJ2AYh
adypkcWZq7GJ4H+hD3zS39u0Byqux9w+ZvrTuKOFsuFSTidi5J3bM7l4UfOqigihBDKDwdL55h1l
pMajAu9TNwV4a0RjDt3E22tOAnd3WqGQx6mLLoZiQSYbEs7c3yIVAGri0FwZj9+F24CUTmjfid6W
qsy5FIe45hRY+XE7PSe+kegFiZa2S8uVsOMA34Mulj9aQTuPkeWoKbNtQUXoeB6+1GeoHZ02sQVZ
qWm36xFsq0a+X/xLJyMu/MnIpo9joCxkZVcK4qmguAiLXMe5ZQprHMKUL7FY8CWo5Xy0IbA7mZE7
G7JSe2ph2Aw7rnTLXYHz0gWhd8qCZMvSTb2+MRHor/dAmYBnrFlUlFOL+/QqFpT5WE57Oh1s8kN+
zLTbc/9+Qkxwv90rISG+R0VJtf/gqehYUNRj/I1xOAiR1m6IZePB0/VAeyMAIzS9dWzxmbaoT80Y
l4l0UZspxTvgeSgr6pTcw15NvQzbWi2/Ja+4bNGmPq594BuR/R4ZLNLQhJ0j+Duu/vn/ItgIhLzr
akitg3V1IDf28Oe/GPK5+zkSSWAb522p65bVpbivKTFoyxzNkGxO4S4OXLTpl8hs58AugwCUVl6b
EIFI77VT/YnNjDH8JkD851461/PNVZlQQDazv3XHwsHjdIk9PNLNVkvXFOD0rFahykJ4X02xiBOy
c72Sy1S0dpsV3iWsKmFIPdzxUqUsr5KeECV1dYYSf4cNEVo6lwZ9IeoH2A7jH+HETjLZ/yzLoS01
egNjlxQ13rYL9ykZgl+wVn3tytV7DOMfBMLUnHUc/f9Ip6kKjiSH4/La4WJVCyD+jNZcKk9o36Sx
4AgTBk4HLWQrt1HMf5Fn9y5RvA1i58osQrDcWzxa6oldK0qQ/onpiT5g4MQl8F2Wr9uk1ej+xDjy
ZuNRL1tUWkVhz4Au6VKHrp39Fl1+oi+ExYejApprUNgQ/MOrXBrHcCk6BK+kbgjVyooVocD/w5Xe
7ZUCMY4+iH+joGRF+NKzRqYVjiYdQlR6TZzLL/rRS4WPO0AOp6khz+h1jtKXgfEfL19S/Kr8jQ+K
2ob3iZK/FzKof9HvRwsJkaOMe9bbC89XYyGdx8gj+eO3PralB16dcnv7U3/FC3E2ocU9HEOASHRc
HP/lA9J5F0WyPHZAf3j7x6r9Rzn2zplB0gFhHEv2iS6fJGOM5f7nKKQm2tIJh9NV+doV3QS5Yzv8
OeQ+xopQREifJjEu7prmWMDRJOBoS6+TLPjknm+dZ6jFaoW+LezRAgJ8lU4lcYFtn4gglYecQewV
Ga9SMqQ2lffxKLhj0FChnb4g+yfPtyN2SyQpQfv1Sm/Go5OuXpPksJAhCIK8KlAaG77o9VY8e8BD
t0e3Ltnan6HFRZx071OdYEI1oV2+1PG31FNPxdJ8T2OTDZ/B3psajJ42KW3D1uJBbC9i92FG1P9A
qNN0K5GDxUekRHrEtcqIhXQjArTbMzgk4u7i4b/trkGjIXKcnnug1R7WSYBHJvI92gU3Zr7o1qC5
2blhlJGodjta/lbbaQ2GKrBT4VoeNCAfKXBDPgpzqLnzLjBsOAo1oJj4vFzf0p7s4mcBn90LZcWa
YkJfvxl4ZNVrCiWpVrowqD7eywh9yo+wJL46ZSYQueyA0vVf4rDP89zVRg3JIp/HWL/xX3AbXDsG
adPhVAftFtmrp2vmRVrQAN1xxbtTKJxR+l2dlokDswcUiOjmFsXA3FoGIUXk/BmGQRcC4N6Ch4vi
PgPbejz0kqJSOesdq8OwfeYFKvey08uqIJ1/cHoWAc43SfWOGxEujaGNo5OMy03XGnYbmSyrnFvy
9hl6Duio1VbUyqaWym2/5DOk234n8b/6mc2WWuLzLqn3VpDEJYuyRRPMmdqyhlcMYENC0vj8Q5Zg
OQaPesWJmz6PN9E4ivEYHMNdzStkjSgrmUMXVnOgxAwXP/aOuzp5hCBYhIoJjgomLWoEjImytXCW
qnga6lTuQVv/vHVfbHryGT4Ne4n0kmqKwyK8xSTSVWO5bgscOFzlaZG4+7qIWT89kREH1yiWA9Xl
qq1CeeK6FX9ZP0a99livlDa0iVaczlrV8wK0uwmMZ8ezXsddVjO6YsYnXhi1n8X4mE5IQdCsfG+N
P4M9Ane9OT95V90bfPV2TJJC19FauFxoA8e7fxc096/Ja6ZZUv8SLGHnHrENMD8Ah1os3q5hKnTe
oTye3/PtDJSeFA42wqCn1E8/uUlusVqW6rGjjEmbD7OxfOYNCpCeHrOLMwVb658nFqyN41bZnxKa
raN8xPTrDJ2A0jEp/jfHAB92z+exUyYguZPSoasaLPRRjzOq3j6XncmDbB8XL4lRI9Pt8wm878WL
s1gcGTfhjGYXT3WBQ+l9xIpADTbFZ59vpR55novmzlliid3AOnXVQW0m0vGgg2WR5ajo5kiDWSnY
d2MwmOpgfqk0Hws/th1JfzsfChS3LQTBeUr6jLnGqO9fW932OLuhZYvyFwq8+Ud6JXd4a7Ah94yh
nCyIlhbcAg9XHDGe2vaHGRn24Wcrn6v12M5wVq2Z44lBk86IaqwSp0OORO6OiUdyk34tpfTc/sHO
O/1I0ktZTfzshj58WvyyW+L0Daf3KXUK0cdW2CzXXHdc4c6jSMOY+u55qSaABB8CnHwmrtR+KJrP
JIc/HASeWteSA6gZN5uaqe475JJs/e0DjYVbrvVFpzHf5ZxN0qVoXqMpyJSzMCI+MVDFd4nNz1Cl
AZRVFh2OKM0L/kO8eM9qnOdUFgeQLwIiRujZnv2r6nHmmxDi0YEYPCFsFqgmyHxD/g2/Mk9T16z8
7I3uGOSUFqPHdQAGxls2p6Or9lMr+S1diRNoihBfSOSFbizvrPgKpUVLF42lsM2RgkdOSBg8yLKu
+C+x9s3/xirrrOn9PO0u1jbv7/bzYKURj8JJ/oE/yrJEEAQdTMw6goGOzmh88YqUlopHSjHZ/Uty
44IiI0/RsauKislzdqbgoYU44ESAQUGyl1NMauJDlpPzIUwFs9EGBWT7BPEeUr1HQVRNTvhah1Cp
adWD/pAFCGOjSN2rr0e3M1TdANOLzYd1tn42H3EW6bvYvts8Kl+WKHgWquXOfbeVrGZ6zWX8qnTU
xIuAxjLMj8WRjJBYsnOgmQ+ZE+bGaul2TIzfe5taBOWYz556yiidGrwUcS74BJJUg28DAjR9M1b+
7KV+CshxUGXZmdj1NW8Z5PsiXxrgJ8+nOgmz44ahMggYPRybfi/haJHqMsiAH3sR1FhLBofq+t2a
ZhCHDp3dKiuBDYjc44fLsZmTcNCclJEUEkrfzv+g2qw2c6H4p1aLIqC9hND10iqAhofhZVYUjR4N
4ZvMwxYjr+h7ddd7Lh33vRtOuZ5DLZI6XLgLyhYkCGCehzxpmDp6sPm6tV5sNc5FQN55zkKV/2ay
SOsuj7PSZDMcoFUPwJZTGMOl86Xtf7W9tOKEtInjhMe3wzol43lshBSo5xLJAjbZoBQNn7WG6gj+
+9/Jq5wXv809c4LRgYETt3+wZGyAdVHG/qJfa3hptkiDBglx1kTB+EVok4fqyfoC0w3Go1hSn8Hi
0Z8edaCYe7m9130pDnj8ttN2cjwfT58bbzJQMACCgAU1LSFNdYMguL6+qR0QykHFGsZD0RHSglAY
WkuKN1L2U7irseyEzzOgrc/k6279mVEHdSPwktavaPmAr9oEV8WUh34wgmdmTgfdsVI7npIHvtK2
DmOJDtGtoUXkKuzE9nuRg5L96zw8saO/zmkr31lSRQQDl0l7aRLOL4hSkEVytooyWZzmFJsLeGqK
HMyIiGHQwbo16Aagoivj1uQ5c2RVGi0QSe6lmf2x+UNQn3feb3xFgvt8JwRbtG6l6gZJMWzpqq53
lNbXzwjW9i07gDqCV9F04sMK4Sc7Bpi0J5nZXAL3VvxI9zWPd0fkpxOAlN6yzZCQWoa9leV20ynr
JieXOeez+P0TLPZifery/JItBpDvOS7NAWB+Lp/Vr94iXIIGtAGPfSkTzUKt/0y2haC80Bmj3BHU
iFxE/hAT9znREVu36BzKyD0dDMdO2fIOHboDn3OmevCiJxCq4h0xdnsgH8gQQ6HN9apEQpmdkpzp
b+VjypwG1jDKMt/R7PmsSBna6FXRcD7oOrpvgMu9r8fyCcBmmyt6SPEIvHQYifcGgcuXMmKH/gVQ
qLMWkIhrFDXPv938F93KvzE83qaYrv9fZgRfqy3PSlt6F9wQPxhxxdi96f7xKLX1bTHvNWgYN/E7
dfUACYU8+KYlvpyIogaoRXjnTmNi/bULowSskwtSCkubpREQBDCDypR1JmHOBafbeXNq2/gCBczq
TsYjvfsFhgkn0MVC4EMBKl8zWbAOgU4LhXRUzbixhFThoBQXOn5V55yZ3mgSe9JAsPiP4fXMYZmi
aRmMof6G2pSBmQvDYr3jcvI/b/jvWvU0bRUM41uKOsfJaW3C/P0syb8yOcokMN0o2XD0TN4kG65+
rAetN8sJeh3RKfxQvapzG1+UnTj2Xd2k9NUE3m+AEMbFLHZiNhlcW2djSXmIzX6x0ZiQIZ3+xAEa
Ox+uEaJWYD6G+MN9pjEmsBSrYOMMcXXHuBk1NQ66LJYwYJyK25eoJAS/uh5p+HjpBwPNvWlXhlOV
HuD0u4BuFxwFVSM0BRCfvtb3Ou/8J7lo0tlD3mssbD4khzbYtyze1wniOjGSKHTOeRhLbyU4RQDD
QpvlVCLySO09hhgRxFyVs+ErSDMndu2BjyxlvkxBbwnRxzHHLowNcBhiCjtUGyr+xK5KoId7kUhI
AFP/d3m0VdyPqqrpRH4l85KCl4ILml6IEcTbXogLABYQDgMLbbrAobOWzs/0GdtgdlP/abiFR1j8
kuDgbZcyftflaYWswfkWr6a/f//jCVB/OhpxnrlHOV1ril81wnWtkq4mZGrYkyzbWD9QrDgpCEGk
9tfv5RFArQ0FqeYYjscsALeOJIP506yjhwFDQ9KB4rndrYjn+DOK1FZ4+OY//1SYVK3au9edn32t
TuvMIzTSjDrTfN9CSYrl9VCipDzPNUnugtLA0/TomPM57R3+9fYSCi9o5HaBRDQqEpWVP1mIL/rb
ZYAHBkiU8dV8QzEE9ta6oEcAYpHU7aZmhNJcMxxHrrn11Z5AYjUSIz+v1YOSdPRT73FPlZsiRmXY
VpXvytOZSz24g+LH9BgNhP+gshdZI5WWM2zu4LthCtf+BjCy7CzRfIgbkQDNjpc7aI652+1+GRVS
eZjupQugqnlGyzItQKvF0kfNISZZEZbrmWjgC4pGCf/WLYmLgVkQwCKGOvb4/VwofsykDpUKC7Ew
jAOVXwMc1frb3Q/uosrkCL00EZ177wXTUAxOshcCk7gqiOsgOJSBzt45hQtd/28M6Tx7q1uqbTT3
YOlNqNEiz12EvnIReftSbayTMChh43JB9duUTodUqEWmCwt1Kf7Vp2se3OEGRn5tGP3S/Ev9wFeu
ED8Z0298Gls0oV2h5ZPv39pJ/bZ4p/hAmtxDi/5cMCM8xsp/qnn24loyqSSeAwK6VWZcaboesbKS
2ZR4zIfNCjM8VimmTD5B0r0LYj1jm4Q1Y06kcKEnhXQMCk70DsK0xaYX37K1eZm+2KV8Mh4wcJuc
dzTi+EE7yUBzQaUYciJW4I+Enpo/dHf71X5wP58vM1ZZXn84maFK2gx0+Q9azOvL6LID0zcuisra
eNYRJVHuDJfdtRqCHrnqkrkncwWOVOEc+5cKaP7PsMntTNzOzrHS0k1ic3Fmk021E0fRVQS/pBbD
uylXfer/kJYJGrGE6QDxFVqII8agptZvQbhv7LsTQa/xeXPL9B9clUaY+pp3rlp0s0ZaAEecEaMk
qBH2VRbs8FLaxdf2avHYG4vnSjRuHORm+HCJYS7eL8J9gsjl18WQHgY4NIhgfjBD1pCHFuxd05EB
nPEiXdTv5PG7YUrK/nPDqOqGIaMQ3Z80Tu7j9x6ipeBAFqt2vKd1PH5bkFE3V+rvsSWBTpLtClAA
RKH1hJ8FyfOwMilQz44d3aIE5Qkt4gXyD5I3BTJYgKqly4F9QfkqeOV+Y9Js4kgUBO9NStFJoCT7
XfnfjsCmt6BkepheRJJVLv36wEWBEdIoRPc2McaOHbcXVg4dSIjxwqqMgeAsJ7J9zEcooMWxDxJV
3qt6XwqmVWiIKxPdO9jXADElSN1H1Wpj1XkABZV5Fb5q2+NhBwni/2M0UyrJXYh/6/X5VnKdDxVF
HZBIWVoZyyxvzK+PX2ep+F0ooEp1SQqO+nQ8tn9jsjxgU6roQQtK6EKwNgdlIssdnwQ5WZuI13rr
UPrPy2yTLMDHNmPnzuM4gPF0nHfChXt6V8bkCSSo5V8EJsv1q9Ml0Pf3NJb6l9yhey8UATwl/mvH
B1lO1Qh2JabT2h5gSZEn/Smx/yU7o/svOCkGLxoaFjfvp9YziCTK5+PKpKpg/hzXrR0Y2ly1ZuT3
pHOswCMwl80QszHG3/nnKc8juKB5h3KuTUCdbCgkpmZXAbA9edpcQY9tTsCG78+PwQxA5rtQJCLa
EVXoasPcFM/2BPf3fTpfHY4OV5aRfQsUQmrsoOACbbNbCX1sfX/ubUeREp+20obvc1M/Ff7MozHM
M4KyVOWdd0I+87eDeYAgOcKGD6xnlC8MINAXzeGOm59iKEX9SKIJfzSEt82Xs3xa+NkdrhaO1RCc
0PQm3WrOTbJpjmvDDDPC171/Oe7Rmg9bdaM/FqLzR2GQcM6auOq/mf7dcN5mzalq/fmZpcutZs32
ak3EaJaQHniCS1RbzhJHnanBQgiEmwIL+Lp7gXiY+Y/DEKsHg287li7BxALRkGU76grwaqAfwlq4
w/BApLO3nKKStRtaV3OqcPkqihIHZykqTyXrM//eO+pJmK6HYjUznemMv9etQxc6cK4n7pPHAV4K
6xZx42yVSShxg2VCoBJD1awt8roQ64YXWevCer4Ka8RUjI7CJYdlMs4GleezLFu8Ad44j2rgSg3H
U2F/xR5qZU0BdCI/MWveJhCwHB8cNgcDYPYLnD0t8dxi3pPpjcVeoi1T6z90sZIVqWZW0YMw4tMB
x75OpOXbmHL22SGpbReDCIogbRuy4RBqkzV1grCjxN6ThWykCUsGIeKr5o2B9OmD4FUCUMg4y6Uw
ijFtNdERiNL4+1dwwS13Cow7CU9eniKgrzc8osTVfszHb16HE2RVrJygRc4k7vf7nnPtHu4Sx/UO
6y3r8p5XRIG96zCDvny3e3L+dsZ8vLEladSGzf19UuDDgtdCYaZXj/rfZSSufvnbXoJUvA+zIvzU
u+4FeOaFcp7eHhHVxbLp0PSNIPZrKBFhaxuH9eaEiKtQUbFDR/jkMw1h8Y+1Zeu+6L4DFd7m99ND
87uM+yTH8wRwgK7ahlN/RN8gojzFlkP/ZsHCPNlnXF2h2PblqetDsSstI1kC9cgjFz9qpWHHp2ah
IBncbkUjKAjAUboLEtCAKEe4+v7imSir+G0goI/v1GyuFRR5uRAhAn0nIq8nrBIVCskiru0fsrSY
9wkV5+WQuRt32MJ1JsF6exlmqHR5R1eAq8urmTomiFSEXGmkDLwiiRXHg0wkVY6LIbhSM1wRng7A
UriuSqwLtDo+qRRSYGeR63Of9pIoSJvI8TGw9IL4x8KrB7Lj5bN4Ah6OCG0U7zhRno6abo6B0pQe
nXyUPSxNVppbQwwQ63JogpO8Wdp0ovYTVlVlIL6PTq4gz3Et9h2CYAH8/RgqOwAPFwYnEaS8RKSv
VzlPhypvqP/ypmv0XO1YyEY5Ihggtm17La6pDUfsTckj+iTxpf5Z3FPlKftRT7V2Q28CBtsc6Rmd
I2QzNdjXEwCURCEm7bWMeuZDPQzLcydbH+IWZF4+gF0oi9pqbrgo7b1ldj4g/WzZtkOdwiboD01U
deGMYF0vTk8+/DFaIVpFeedkEhIYHVEF5Xe26MbLYJ68EUxPoY0SSTbU+p3nATWoI7Sd0w3Fumi4
AgF34gPxumEsEo48WZ0CJh57WWLYVXd/p1g9qCAsQKFkITLqwdZFW1mN3WFZ/5JUCBLJ+u2SVi9S
cuggRWO4T9OYeUjrQlPRxG3EE/TqoYhr7Yki3oIZ3NIHMw2mqUXjofO4cgsahOIXyDbux37NgaJu
pSlZMHe8FAbyB+tXldDoguKHvXOF0B7BBT3amKA0qduGAR8BSxachJFk3mntwB6Mmt4oMlXqrf2r
Fn1jYQLT75o6QezqN1F26Lc6SBGOmaQ01/nX6yyamhc2Y/3oUUwkB8wjQ9dkMrUVuixf4YeY42nA
fmDo46ecZpOQm+0nBdSu0CwYQLsdFf0gRIxuuyC+O04hB1Pjky5/7C31iB1yYAGfz4VBeZvTo3NJ
ex+JqeHG8KE8bISs5uZC3dKgIEUOHWctaQ/u44Ys00yqrVCpDhMorUDpqwv5wQkClzC/ybydcTsf
POZK3mCilGuhSlgVyws2q2hnaJSvbcJ2Ot9XMuR0DJb1FE3A5bc1aa6qpfa8Kn/c8Sui1Fi2LZbF
WykRCA3fMddzFPHxkFaHiZfTvG3/5a8GnA8hOnDacL1CMWsl8w787hZKUaCQVNz9oG/yVhnvVm7D
qPYZZiuWSJv+aVbcVAmbP8Nwj0cd50dNq0YoYttIsNTgOaQdlaairTJ56toh/9/1+5Lh/OgFCsSj
AJ2CyDw4om8BhQplOyfQZAD12nbuYu91OiIm6ZnA2IIuR5bOPWm1NBEY8Nm0nOQn1IDFf4kQZqdc
9+Id5F/7jMbCSY0X0QhHxxsztgRF3X3VuasFe5G2lWQsVTxvgjijosnWzPgOn1cULrdds/QyHAqO
FtXoDY9dPX1gzIfAwjMG5Z/gj6FUvrG5vSIaa9AeCExIXC5kkk9MQ4vya14EZF9xCJfkdKI/Z2sl
GlklB4NcDXJQKUBuK1qN61vFPRUeq8cAqfiS4Y6dRyxjyFEEejnDTL7moW+0SJr4anWuDrvuAB8C
cb3NLG3dxREOiH9dzozEP9fmfR18Ybb3O/da5hFfXXs/CfwXR3Tv8k65ayhJ8VotD1C3dS+nim5X
obXBNvDJ7/NoxLXkdhrk5Rm2ZoU+66Haj6HCM9GhBVtYpqXBJjzDTwH/oRoxFJ8nWNnnsoAxhUSB
T7FAtjlKovnPZ1ShcaHt8QJB1gQGpzOvQ9/TFEESIe88sgWyvMnN+nKVdMbqE40yMhtOYRN1SMpL
WLkmYLspiTPdkzy0K+2Hps9pxsLBeDmbITrGOGPnCpUkftJrU3jEH7Y1GbqB9h4koRFV+X3QzIwJ
1I8fAnqTr82GNepgGqk+Bl1tU0EyuqDO73xJQEliSN9Xz8d8cWpusDOsBySW6J6ph7h+NYQ4ySpc
gOlK0TyfZKcV+KC81+GVUlohmPQzDbGp3WUm6bGD2EMasT1lU7Zsj0PLNRKJuconkfrF+RhZVEci
pIaH9zHUVFeR8K+IfVv2IILejf5dDxV/iG59nUYhH+4r1PrL51K3SoL6KIqyY/2/Frnhnhf5ecpF
5Dwm+LtAfPzXSO2K4quUddzegNar6UTpKYLPIs8A/8N7K3X/MLwSHC+0LPGwOD6Izygfwj+PeBEi
cCu0YDTH2ric5uG9PFX6DVOLeuHjOhZ/431d/xxyky1PC0xwD+cPPbvbZNx8MqM7xGloZooctj6h
E4FRncSoRXdO1ICyV8XXEP1IiK7I9ZWryTtU16+K46LLHjbOkEkyX0ofF/5F6FtDwg+T0aJO+l3q
GitvUNo/cOrnJXNNG8ke+Ysl7V3kHUQSj3sHWIaeSSj76+USsnzl82D3Yh4sCA2dZpviZXCMPtN3
wsZFEDxpJGwnjKUGsDi5ETpPhfSftFCTQqfQ76NIjk4iO+fk81cbDYJhWFutN0d+qTjTeZ6kZ+X7
oCnqnHiyizN7Kr3Gp4OawpgYOAKY0CVIXZpbUIm+a/nX7XIiqpDa/m+I9jsodHTKQ+9wp5DqwDYk
sDJqPsWRv3kAp94dakdr8Sgi5Lhgg9q+W5nKIO5HCR5UnMTWXDurxFd3s+dXJae2N72ZXF5MkEaB
YDY8sh+uiCCOxVp55nywRR4/N/jELMvPAH1kU4vKoRKuJqXAsNU5fKU92GTvFJoAPIQZVUbRTbiu
VFjwaYP15P3jzACEYW943uS175f66ShjAt67ZurwRMqQ8LdA/18eGmPbMw3GAWHVfZXG1SonhQi1
SifFYR+pyDZ6zGR6L0YhfihIfOGBqszxgGo/GoFm0Np9p8va3OFkqXajpDZsHzo2matyWSDJsW9v
FDtzDi1JpKgzWCPMf2FwTr/7TIK0T6M3uJOlnO2v+Nsvuwv0cKZY15zGPt3f9j0YcMOyj1Rr8e3D
KFS9cGj0nXAHJKCF2U43djRAUlzhF2+Bqtb772vR+Cv9fJ7sCda+05TAc9V8R+QFfu/DsrByQaIf
eiR+3G+ia0BFEgluXGF0R4vRwaPvfIUvs7zwFuUk4o8l3vjSO7WfALm41XcUu78QQYNDanaZoTQx
hFv1jrFH35d3ccVL9SBP6hV2roOX1E+ZV/apllJPH//ASCSEu08J5eBckunePv4a+1+gbfYJ+Wfz
oDBiM0E7uVhCnoZgI7zjLfnOB47BlZXoHNEr2ySQFvPt7WJcJbjUjqgNgLoQsFG1rtddOGkQFZbe
ZDe9Im6JLzN9VgUMYNcp5NYbimaDq+hz+tKOzUkcbk4TWZbiPQ9Kuqs3D+u40Mbcn7szO14mXhFP
40GmY6/SEwgzuRvgYvHv/uCpP+4d5VppfpXCJQJS2sKd0/jv5GHToHPMK6lHulNyfCTrSkn2EESY
Kl5dlNBw/6J49YW8tgKy4mDHtIpEAQlaLIBqEQnX0Pj0GJE2pHICxTRKARMg1XNk/9PRG6ZXUhLu
6Chi0sNkf2yXhq9nbq6+D26LkQip3XaiJCE7ssgfjhV8mC65+ENVTM+zk1i8dt8tbXCVIEqYAgtQ
uMlHF4I9TNNDHVodzY3MV7WiowKQlXlvW+UcQlmijDoHUuovlGKnNwKMuDN1Uyr5tZYHZNLEcz5/
1CyBiBBA/RhFXNyvL0ZlDOWB9odAeTPPBtZLiVV6r9XfPfy4pPHc7meGWPi0q5qtpCQ8VqvKOzdr
Pwx+72FZvsBya7gBomYTfatlf+PkT6VVHsCXB0NgfMQ8U7jc53KfT2hJ4/jN/eruHdpmjN1MIGG0
w83LRHJtn37B+VcP59N61X9Zp4Dfb1Wou2h0OtOEjvdubeuVU7ufh5UF+Rs017l5YcROaCcK7wtT
PjXvFuFaZGrdY77rx5uCinbM+L3Pr1AOFHSFbw7dWQnb/Ffb+kbAYdrkuPGQGnjl7Ix5i1ql1ci6
1x5yFh6ueitzZy08p/Cyo0q4P1BYQ4MkSjnI8bcWD7R/2ULF6jfC6jho2cn0t3Kse+hpoO//8sEp
gp1GpP03oEsT1zM5qQyshXVhDF5cluxHlZoRIcTk92Mki6FrYe0vTlEntizSQJU6MikLvRs2bVf7
Ij6CepSFCbS9wHCLKVugE+qAioDpTEll8lnuEVdo8tqxhLBC4I9rzGVrn1AtnBwl0E+Wuzt32djS
bwrMJDL3ttrP6h3RzaFQK/C7+mjh9BCDs9wAV43AiisdKQllv3J0Il7ip5AJC91ngCYRPqS38r3e
IEXV5GWlALfHPYGexMVH+ulFwxf7dVww6xKCLHKS7nojz5eXkdekBr8gudoPguAKjDuXEQj2u/Vb
pK4Y+1WP7tbqSnukANKxWdxFFredyitXKBXjpVERjhmniX7LjuFis7pebwcsGgBPqb+imcbOCLzF
2H6zltdDDybQS+cTSn5fcsDS775auQmmC438u+z4aHDYvYewnE3ZQRmosPScQcZ5BK5GRfwcV1Fd
Oj7COrjrZ1/y8mcL2jGV2hsGKu2nWEGwQx5jAq2LzCZYW/bdRUE7MpcZh31+Rn2F2meqE0qcFhW8
WTa0K7Yayzel0QGz7YELEeog/PHitR2rfGRgWvNCrhlY5irYMz6mFY3bqgo5W00Z/acWu41ktw4e
oBh55HNX1dVHQYYkwHEprM7FZ97fxbv0hbPp3GSNpy7WaVmokbhbWPQrsC2lIbix7LdW9Dg9psMH
EVuaModJlvSxZhuCh1npH4xOedk10/qUUYzVzBFmb2SjlmQJqnR4sEvfOgEQ88sYD+Qe/5XLjGli
7i7coTNM5i8lm4ZKvsnmBLw31FdzJqgEMf/EjUNZ2rJwjWXZ98XXAKCaBxhR7qefB5GFvjWB0VSb
XOQr0hZbWtDCElJLDZi3apX6OjUvvDh4hv6rsSJ3RIvBXE7+LUjMRLk8EnUO8EKDqbYggTp/nsO8
eWR7dYa6sSs1zInAnIahjwksw1xoPJVYV6nG3IIfmoUG4q+joLDtXdbHLNTn0m6B/R+pRcA9E9ZY
HE4q0ZZZZGCn0i4RzYZ7Qa8q6ZkKPCWmkXjMq6ZTARSQIvsIfhvTRpMWTXja7QiU03n9R/QLH0ie
9Euw+z9CZCOHk/E34Xzg61i23Ucvw7vShYe54q1pNy0XoUrwZ147ey0l41d+iHf2ojPq/HGVaw3m
3S6TaW5lhA5Na2hubz+UP+I/cAxTkjos5lSK7RoSDdW9Zqj09A4xIzRAUiwf00f+oX0/hYv2jZP8
3fZV2LHD3N7l1n8KGviM+IaFXbzuey7+E4GxporrJgOzjYW0T96kVqTasgjLUcrJzOpQx04gnLX/
HMdF0d1YjzsX3FUYbj0dYoYiB6/8w/qz4vUPz4hQ6gAUdpmGj6o2gCCK/Z9oBLdAK/Htd+3LXz5Y
yI9tAgiIF91yHooaEpT9dPOvJdfSoEkVAjSDvUS5dnghBuTxNcQnndGtRuEIa+guYYGe8fRsL9WR
UjxeBF9mmwdkuYT/lo+PjS1yRQxHhKiyYTu55cL+QEr+Ngf3EUhfdNb1/uP+y3emn38SMXVuke6u
a4L94d0hUVerZdmGYVeKkM9qTiKYBucZzqGPjZbjsfUHNgcEafwpC1MJtPGwGi5ytzTnnuIso9Ru
RyWWGAFDdyXM8pgJcp9/iHQKe0AXGnHOLzvTM6jfpqL+2w5v1Hvelwhle3pWZaaVMLdIBsdyfeeN
ElwYQNhqxKIXnn3vQ9Ipb9Hp3Kg8ShKnia6F5qByvH9YUb1dd4oyxzhchw1p52v+AugcSULP/pOt
G7EWkzPWRQJhKn0EL8exWdUx7ipCtfRo5rHN5g5zmcwB6CIneVFThu1iosDAxavlsu2zr0MXPfDV
BsDDkaNF8qVdgoI4JZ2x8JTmPLTSCVj7vRaJyKa12CduaDSVbxWzFogZuE71szZAIM6zuC3PPRPR
sI0+rhmRuU9cWrXz0LzCU/mbip4a7nKTx/Guxu6nv7R0Y/qEyr/bsS7RQOfYUAHyEm5BrCQWh2Ro
Nvd97a0MBxk0zymyfoAmrXA5AK9X8GsHS0QcQTdNmmizgjB9JwVOY/93icpsZCIic50Wy/K8+gUk
+tLokk9dF0MsFCIWP/woAarZdCf8pRvNvuNptAAsSIOtQeh4BksTi/wqCSbBM1/WtxwPEpz0npXN
F8UJrUqa5udXqKzkrUtw7QJq+GGt++Snd+F9MO6ALJwxbMSWdT2XlYE18zn+JLmsyG3+M/w4hbaR
d16fySnjXgF3arAwNeTqxFyG+5iuEPpWq2e+bpfNlGpwc8Mg3Sh+jSiZru6mms4qVf9zFbI9V8nD
U7+YC8UbkicL6MXArZuPBerMPQSt7im+XKE0k2rtD4LOhuEbe7lEZ1HF6vkC49RJ8+/WFpiM5hRk
HyO/8cnqzah0xGVbnIzpWZzHxgX0NurUCIg5ukScr+S6CQ6iSdZwGnDGH4ptg7+Kp3xmWP3VafBU
3IXOS5GfWzNuGKzxDDwGobjzZsixrIvtswDW9pxLDRgS/Qp7hiIVPe+aNNqLRJeCuPX7tT5OwGmr
NVUXYoGLRtKsDnktuCf24OxNsTeQTk+3t7l4YNJDNCzCIwyuSGYKPfcpNm8ialowvMeya1n9Zc+z
4Uj37LVHbimQDHD0V3NBugAhO2E5wre+t4hx20NJ4F6Igncqr+QsVCexHbnTlVGy1BDAuVaJuW0K
VbRmoLromD2juZIs8HiDeQY+SrF8GyuINFIxRMNyVPyc/QFUcU6aNXJWOwpW97uRcZ8SvYBiH7Vl
2Rdv1R9lazazJrrpsU/X5iiStkm0RRGvlusKCqt5TNsJ4HERZ0Aq0sitfs7tcGs8GY+r2JBwub9v
9i+enfE5c4DEjsg2d1joeE5rjwRGITUBmN/HBAoT03vkGvKdl1HyWSfDOvyldb+/t0djEqRFt/xr
tTPbKaM06CTuN4Up7byqfExSk2SFjJVNR2KcJyAcf4U5Y5eGibY7bqCH5O4kcEJHT3Wuzgpfn1os
u8NNguo/Jh9TLRVPbkwt6jESPXrtVzP6BoPMvbXkOXmFQm1Fk/QzTq7U1tKq13DzzRi9qvx7l2xG
gEJpose8Gos2pZ6YLWaF9M7PJmxKd7MJqtHQB4a5fOIMAPlRlEIvEE5n0CMegO4IS1y06X1zGI3B
83s9kHc/3IKIdFygKclyc/Vh7fbw1ZD9fpsnGLb1diezdDsSkh1DoO9GFaNi0d1amul0ASUpCmwW
uWcUwkgQ6VY59giCtausKW/ot7ZL4tmXqvhr+KRrf7/sXu0iz/JuQFM1QzQQSGY352b5to+tkjI/
aIz0Be1fPnMH43QhIrzmjaRE/pIr+PNy7wwY3afkxW/NVPo7DEhUvNp39UQL6hiL5lnyZKNzyYlT
XeQl2AEMgzjyhjd6V+WcsFoMA6ZI2HVOuFVhGBySp9F83fNgb7nIHQG6TQ0WzgRrcTuhxXks1xko
mCW1MqVe7fAoKi6xsB2QamH7SXE7Apas+AWdiSPhGclRytopH+upsLBFuXQBDXdtwms0b4e9icUL
mVOVlbgRG8Az4ZKFSwyp1CGKVj25bIAfe+iUJgA/iImkuFOMYY6/cBOx4xCABXXAKwW5yD/GhUUg
8FhU/PB4Nc4vuTHT4cGjo7EohS083qNtKPhg4YtQVnlMfcDmwkZdHmBphDqdivn085Y2+jhaqTCx
YLvzdHz4/8fT5sSScCHhfFbTaMyPlwhxMOA/iTiYo7c+mVDzcWSs2My33ywyWxPE4TiTWW8eR7Hd
EJOa4Krg/KlWtcAROJD73tsyOfPJl1JXRbNzGyYTQZKgPKJj0K1mniV4GfUFc0tGGbusOJ2i5vvR
HUabMwJ4uHBQKGmJSuTBDoqvLhILXLEy/WyJ9khtiITZYRPCbHIK4LNYoAd7H7TnkrDv09924lDK
d6FTH6nZXiMf1W/JK22kXN7MUUaiShmT2GS51tK9UHCYsOc81hRKESjbZRc4eMMwlggzTYWy8ffi
yqPMD7KqkaVIotCEtXQuWtSNfIDlqzqvIrJOXfcVmPZiH96ucVEXl55DTc8hR3koCVJV2LCxoy9U
2M8su/DH9T6LRQMEkosT5ne+mArkvOEcZFo/9hr/c6Kw+7jc5MuT6Oko0OTB2257BPjBvayb8nhh
12EtZa7Dk6xf+5sc4cXGUPY/BuDOYwbHEnNvfHmy5l6EVzuDTCBtjpXDgrgUxYbcmR+wdoL0mq3s
pm1Lv73JmOoLOyJ7qSCPKCA28CPtrW/w1rWK1O74Hfh4/WYHxRI9eZmOG7Ir77MmgUcpD/r/i6AS
esWx+Iu+OmGR3xWfc3v5Aqb03l2fzul4dWWgnmqEmqNzp12oCmQk/h3S3LHSz36RtS1hSijUGNyU
4rk4skbwD65W3xes/LoZ4x2g+M/I0nN039YFkaTPdURacRmoYnUBPOmMCDRbfs0NuC2+OpqT/OuX
67GNqNd0flC1jZpxRHzYMMc695b60bWWUxn+FYKZoLi66HJWRqvVn0igZJdi59K+oefjvRAvRhT0
Xdf4xiB5xnV9dQoFWfI9nJHN0hF1MMyuSP+qh4wnvs4C6hW+oamZy7RPb91cd3z+0lNaBizuC7Yq
SkqFb+okC1W1BjaH5PnDdDNULADXKao9U9ObeN1WVqclqqzdGKc34gPGNJ/jJ4iacIn8VuO/c7GI
CgFkZfvcLezqc7yDJc8KmdCHxwXd/2cYDq1ikS1dFTGJuMQgKO3Z3EzyncypPa22GAYeQ21RXpDB
B5h9wefcY7CclvdtGaRY7CAdYppSpXHaFZLphwiay33qBNIrUvSP/C904imQCa1eRhT+1UfvuTT/
FDwOYKIubKMejB1wGtReyadVPgFGb2fhQyEe+FPNKUOEZpaSgkxvTemo1QpD2HbTH3HnYUJ0SRou
WKybhZ5ZVHS6c8CMpbjDoNNlJtqcjIC+IUMIxGR0pUoDRQfylJdh+nQKT7JUMmVjFKx/NmrHsU2X
4Qh2W2lxjieWDRfuLBX7SXh6NTJuyjpgao9OEoTu7KDXPxGg9QWH5/U7GdpovvXJIwrmDMPHSdjq
1TMSjfxr5Pyz/9PASIsjMI3/lvkX+UqK1S9kqzYPaNeFbFEUT+TEqMlsYimmF2F+eR2X0s0awC3v
B/2cY8/CbZgzZd6Ku9e64xT8MKUfx1VTyMS8B/CXwZPcq6B4tGylMYhhb980w+ERiNq8un/om5qn
Wpuj/4cl11p5Z3t2z5qWiLW9RdE6FnfCrQsSg2IzQ1RqpkLOSO/3uzQtzAP1ugbaVjEWy/OMaLoP
mVrLAnh1Zp6t4ljSsG5TyXVMeqDK1mQBxEG3bk4cxQqjxN1LWrFMmQPNmYhuZb+tq8jwJVZtap55
zztAqqB5biKMInm7uxS/bOuvKAz1dSFB5/9zaogbwEJT/ljT3c3v73mMckVh2ddRyGz8rmZO44F4
SOGF7DTzZYLww6fvGhrHegf17Mb++f6qmdDiGYiL4iT0uq1pYUKKqut3SwIJLT5/Ef7co59bJuUk
GAjjMcIKC8eAa/1rTyeREXkwQYwfXRj+y+wL19SQ8558XOwW4gustzAWMEdGG+wW9TG/E7LACcNv
4kcjUgJJxJ64JvNa3wZdd5id8QCtpM7GZN8ISdIja+63i3Uoqgk5V2GBKwBa4uxbEiPhysMSPSt7
yeIHrHUH3RzJYnVZTfpvUw8VTLZyLUoezImbQJuWFuvWiJeNFwwvI4FoaTn9Mmi7DBHEIW/URcWI
/tIa0tFfqU9VxbXTZNO+VzXB2WC6Obzu4xOMAWT5baJqcUnk+u9t+wIE4w2jLyPcLmf9A9ckFnwR
kB3zaDztD3ilnRD0YbkQGPLojafUJP8nIDixZsE4sz79VQ81AfpdxBUwm1oh11GJCIbg0LHnixru
uNi6z3GfUKETi0HJWx+1wkFVqaGq3lXg6l5RtFjKMJjh5U0TE57jQWBsAK8+R/T+WlwkdnehgFoV
jPvvpsDqjCEa1noqnLNpzYiDHpOegifK4xYUsw2lgS0RdcDOcoE7YXada5a5ZeizGPriM3ienVKQ
Bs59GtMMTQ4bSNU9QKFxrsU9V9wGLHgy0lR5xOitQ8IZbIR2DCGP//vL9yTK7UcIGUwupwKJqhh6
RmlDbqrpnKS1rMCqYsFLfKi9/2lt1rk4iLdtkTkT9DlDVYHrRcyqg+MVp6xcjri3Ti+UElx7E0DP
rZwSJO9Q9RE4aMvyYU3vMMHx9RbCwJeR/GBWfn39wfGMKJbtD+K7utWuflVnE0yhtR6ouXq5Ck1i
813H26ltIKGRshemXX2gHpo0T+rOQSe/CGkR3znURPHfSP21OPhA4+4B+LLKBSlO/+xCtXD6tiM3
OmPZxvFRkDcfxe+4zwdoHHAPN5jvddfmrqRVM7V96zEpC+zR4c89yfcOi9uZ7D932gHt9pqw02Wz
vPAka0cEKPb3QH/VwHb4cRohTBIUtUIjNhtAIqeGq7HVlZ1cfAgWyXQ5gqDQFQbNyRk0Xn+93yTB
kkgfnbXFJvvh7qBG2bi7UJ6nMkpRIKvLS9W37rfSrFJTCAlYEsPaY+QnFxEeQpPeZvgMfadQh2tP
Xtr7/IhrLO38IhAGH7LaeAyaunDlauoEg7KpOar4uiKZH8ZLTKJ/3Zwgly7c2S7b0/vls1iV8O8B
3jyC7m3skBnhsbi82Q9WiY+Y8NDT7sIy6e+oPfGLgZ7xt4Xf4/7bgF35BVA/i4aw5yFTJocFFTqZ
bfjAWYImgg8xMapgdVGhyMp962L3+PsWQmyH7IKYwT67wW8o6VF3sIbfMXIl/BF3gsMZ4AAWwVph
sadtnchPmsK6bzYODsUyqI/bQPpph62Mj++yFRT4FvFb+Q803LRyI34r4RJGnou0+sHniiButUxa
1PMLNDic8oykcLbupkw6/e3IpQbb0OeOszzNd1kLb3OXk2GrA1N0VCj2lZRSkeSBBm2K5y+g4fZb
p75Ds3c0SW5EJTvg3JxiL34CDEwCKR3M2fdxXFxDyuLAxzmEf0t0/nmXaSMlib5FL7eF19fkCt2P
V39WpTZ75Ab/WlCReApo09Egmf+l6UcP+D4c6bwBBGoEocYpVPEsPAgufVRarwl/JHUHBwDEEd5G
gUMVKMh+/35YwRBlaMtZB2bUFFQAShp5JWE/pcDrJsuBzfApHQBkxsDt6XbfYxLYLvJz7Ne55DsZ
iDMFDQdeTFHVnWdC++Ugy2YDYhUvpCNfxRyNdTrPRfbkUkpC/FCVeyAYbv5LMDYqOQZlF2TohTQI
jzaWTxcNlIrGf0thFOxLBHYPb6u+z2MLpbQr9RkH6bUJqPWs/WuowSqX4bkkE6zwGsT+uCTVQLWG
0e1nQduut0fhIOJdW5PUAjauwJWHnaAdkS7iFT7XPM9G7l4ppYvOUS1HigUnjSY1MO/Qk85rBfFQ
xiEOUuGQVRRwwRVhfD05cAjbh8wpSLpOT59MKZ18m2rMSi8HnSzmGwooyPX3gGhg0ngkKySQ+i1/
XQ9eUsNfZkL+KDN7JU/pA885TdZXN4u/hSRDyOUUQqX1ZK/zggff2cQ3GnCjz72Fgto8NgjqKUFJ
V9UgfB4S3eEwgZWPqdKRLy01hZDfW8+MordQ7lsrI+/QSrTnamEbDh8z4TwCp6aGYEUYMyBIVsfG
OKsGiH4cnfA21W3349uQhP6KuSNu69pI/khRNsUae++jWQO0mzMWQ3MkTuqWF7xRUif9JL1cdPkN
ZLmMI0bDD24xeuh17dNId0/84d9hnOGY5v2ZiFrJv0ox0Q9WUppBuiVHxqcKWfUb8Cr8PnIhP7zv
75qgIv+fbFn394IZkgTHAEHMQQLJO47ngw6IIjRgWvGV+eM5Qk6T44g8C8Amo/ye4saMQBYoEHfk
eqC59La0RtgxPmqaFhuMLm25r4QtqDdOqibSBCttZhRna7Ivm03PLNfoAqIhobehIHKU79GOzhLv
abQEl3SpVHyGlY3KhV6B32ymj0Da5xlOMMrmtREKeorFmeL6ktra3Z7rYQv8w8xY1hXPkxSvN+Oc
4lVGIFglXMOOWoX/wE+9HmVp1OnJKV2n9huo7aKVi0mvDedqxdzJDwBaxaQDtSLmTEgbWKr48t2r
gYMdb6pdBpLMZ1+BTRk/+6ORRqpI6htH34OYryFkwIjEruXpE0TdxrcYaY8Nr//zgbaCT6zqSztE
bdxLXwD9+0h+JFIaf5RLzsGAt1MahNf8sdAOH/6rdbS1eg1MA3aJ3ViHuzv06xg7k2aRL1B6eQhP
P+KggR6u/h+UaTgzqSJfA5i7IVZ7RCSfPSF4J4cxkVFnsuMxTee3kVMNXepyKpc08zyHEvaYXO1R
nkdEUvZSudr/K7osV/pVS8pOJilYcIqLvcR9CoNCMxBGPaO5IoEa3lvz/0SR0LebFpifXCZBvPk9
sIz+GhSCelw19y6NUFCae2qfNVQ0+2biP98P59eGIpGZve5hmgvFOqQJnj40CRIvCrWYMgfi9RJf
TtEsrphzPgV0Y1Xug1AUUUDA75ysZ9vVy5rp0Nq38wH/zwjsTAsdL1uA3jUIqqkHtprhdMDvYKgp
5TbaVFZ2QGXvytAHoX/4XYAVmqkGNCmUfV/CgNok6ITwpMobXfUWkNrlQKVbCt9sEA4Me5Z2TQyO
dISmcE/m/LmwInIqOLa1CEEFckEIg9pfQPsAQvi4VsYcBVZZRWcahq4y1r/vYDuIfiC/qigP2h3I
h7wX0UMqsYyVe2YZz8Y/aNHulkVRMmfwz0/VfDpf994sFE/WLaN+zGQ6lVG5nE7k6YJ1FTgue6jG
CSiKQvquB1TYxJwZOIiChPgkRIR4piRSuINbGisy6a5noBA8NkAhaTg+abfN1//A8Qn/gn+V8ywa
zxNSGxdIrM7qmN205CgrITMr5V9chZjOB5ggLLME+s17VVyfStyxz+jLQ8jhjk6D12OJ2TCxVryf
oGYkH2KMcr+MVGixQifu6gIDBqq6kJyqAhvyWOx5ZjPa6nklrfzx9RQb11UdO1V/z7EWg6nD4Zs7
aZp6Art2MgSLMvGveTkJzwwkfLo/bEvz3jRXLkQI6/viejFxnggAuryEKT8iurxDCNH4oTo1V6Wr
cnH1seFylOlM+H5rIhouRX1lBIIwacZ2j+PjGtiVLfpIFj3Iz8ATX0P6H4p7j9xP6LG+OLuQaiYp
tfrO2zZjpOWWf4CnCkkjpMSk/QqF/zKtnJBzcpcBdQw/Jp4svdVJAk2F4I2+Lh74vkqwG2YNCD73
/w+9Z/maAbf+GiRmJXCtmLDKJxKiw35d3601DVA8pb5nQAmO9yaWps8xNw6EVZgIX1ZK/yiaIjVr
CiBjwdclI7unq2X+DGH3zG4p+l8B01xKFoT+jN3IQ98f+hFcK8QrT8o4fnFxncsnJNqNV07speSf
JFwTosTJ6jkNdxPlTYYLhle5ZF2e8iIEsDtJts4Ned9I9C6H0qya4QmK9EcPaVn+1wd7eMeBm13M
K7ODpPTUgup+xKNUl3XC6osk8Qmc1jx2P0fzg3j/RgXIyFtX+z9+jdeQuT6W7kzb8QpqrNk+Df9G
miU1dC4o42iSkjURx5lXvGAk0ubZ6bd2z0z/waCMnwIam1QJ0WYHGQWXjekJZVUTJYPZr1iFGw5a
LWU46xczpUEAViWRILje99JdY6TEyC6ZLVo9u8J3zhcY8qJoYqF7ZckkxJBO+PqKRhQAfUyDDWxf
DoBkDBav8UB2dveGvvQqU2SxipQkpvZ4vOOxyHgqs5seJUQLKaf3fWVCkoXY8PXyhHgW4JNJhVc2
TXm3udV16VDWDBMw7NUM1pR9MzFzmy+u4EC+A12K6BVTl8Tr1NCy9dDr89+n14f475JNF1Lv6EhC
B98ex979ZTyK/+YgfVxfQxAX/+1y2iyhZRaPOjJzDCJBxj6O5QnYVsFv38Y7fMdIZQrHhIqQ6cwb
qhIyKPoLhJV/TztwF9YEK1fidcQTfLYROrOw96Z9obReQghbzY2V7Oa81ipsiTwhOrRjB+2dGLro
xmRY8xjf49kweq33wlw2HRreOQIg7npvjToocxW3bu+5LM1VAZxEcZW8tap3DttPjUtK5Rr06Gq+
/xhyCNue8z9bjCxFsUysv46T/u9h/1o/dZcd8rno2+zxQ08unLFkd2Cb6sG8G16fccq0839Us5Qw
52G2dnf4JBlb+r/1N6nOgzNET3TttmKfQWaEBPEaJ6/aLNVTqHlIX9kB+8rOdeq8ADWu9e7OQ6oH
NOZ0CPqZcNpIRp/oosY2RlLamnViix43BuUcnpeKtfxTvNzgI+gO39Aoo7rXjnfr35aoVyrdSA9A
sFSlTArvUjJXA+W7gueNQqu099lpHmpH1f7EpbyX/kOZm3kTze+dnC0GDUn15/gbfmh/brlh8YIj
aV0R9SnhfQKWKp5fwUgdJF9dz1pEAzH79xVKvE3AnbHpH97rQmFpzHa6KWK4M+trXt9tJtF6q+a3
rqbKB4RyKUGb1PjyuQqYn64Y2NKSCVkZ87niEIqZ+OksoL55j3qyKRCvyMNYrUdTZIrkHnph/XYy
GWAM21OG3XkZ6b1Dv48YGxTmBrFjLQ5a4YZVeC/0jxOxm8cZBkCBumG2vJHND9V+QYikuD0raLuV
Tk78X6YNuhDg/m8sr1+svPWOX7dBiB6rsvQiBAqicHYDH4gxmhRPS06AhPnNhlq3dIdudgp9JuqW
e5/QmySK7k/On49AjHsjhWFhP6kMOPixDptnUg3Veekr19RjZLHRb6CMGaAf+eDPW8aH2CoKQvPU
ykzUz17ypWmnNkN70Bqy9de+w7CinpVbFhLDXIsaASiT7nmCWuGovBphI58ksYs3z+5bPoljRSn6
C7PON5s6ceQ1F2vYpHCtx7IjQxaltOrVdrGgMgKeES1dkGrqpGKlwk2nYDNNjG/emK92UQnJ+m/T
N+vZwLrhGlIFuXAf2n3ODeZYA3wM9scbacWRg72tpoTAZhZLH/nQhQ0CoNBpDTnQ/TI26kBsNUMC
pV/Axil6cVYAkqGgkxFPhfcD7hR+xHT1C6Fr2+qvQp4e/5eJxT6EEzK63kmZ8Ad4+/zHPXy0tzVv
Q5UVt0KkOxAIbhsToOJYsKnwPD2VU8GBXi1IWNaZw65R/HX12LedF2rC+KKbuIaOd+laW8Ac2foo
R0FGgTKjrzPVVvLmckNCF2pTdIXdOYlLqpvpFCGR8OkMUMifHWbenZTX7EAuWsQlzpcSFe6f91Mk
FVPYQ7mPS4B7FuwAty8USPln/ameVb/fDzLLJNtivYoTyBmOgYEFu7Rs+D0PdPVtZd0jEZAvqBW7
rE+JWjmloyxTK+JVo/oyhFFGIzfUoUbgxrm9gCu0RZC9PDLG0OYdErhSRll4+0l9IrP5pBmFBorK
EKJSoiT4TS6g1bhrRjtUqJVhSCIPW2iS87S/mfoMoSZyc0S34NQ69CNeuET66lBx2z3qXAlQjR6X
OrmBVdk2+KqHB0tcLmmmTknt28ZidNTD6qXufcVU+SzuqyUlISGKyWYZcaR5CMnrQdsEByaHHb8+
GTAdBhiUiC3e/B1UPqzkV7PNb8xVkddv6yf+R9VikiLH5Ehv819aajlIItcbj0iKX9Pv79NOzTQI
3tCwUHKYOGF58Pqu+pjuo+6SxGPFWa4snJ5+ygolzs3ipiAFfiHgCbAmd2z8uSuZfFnwP/PSA3I0
RifoqsDOJoCKEQcyQ9ouUODFK9/2vbveNPf+tcEvXSMPk8j3w13bZVdy6W7cQ82dNyjE4ZX242Xo
nIeziHLqR3DaUjSEwudf4/qTnWhM5Sy6I2ClkofVxZFTMymbUGjEARIwtrf9zzxPXMyirWbUKeZM
5WkKQ4BGnWEPFQuwkXHCY62/c66ZMgVLsp9ZnJqY9TuU87mxyElCh+cELYH9xBPK+VTX68E8d84M
YQBbkxOaBEUeVGuWZZGRYD7eb1i0uzZXJiXapNvAO8PtMU3bljHsFF47zfzrcqTxhLyOFxGU7ELF
XZIcZBMO+8lld+EQOvvChHRQvNxaapOyIcF3TLtSMOIbrTd0e6ZmoniX51k2P8AkhMVV+mNAU2zQ
buX7odfqxT1xHXIE+GLO9+MYcUorzn7fF8WSgAP7DkotoY+0FoYYOp8XNtitSB5a+U2EOyLjFu0P
3KQU3s99cA5jP3B0PBRmKpszRGW/ZQHybPl4gGcFeMqqIz0JSLFcSJ279GLnEBsmqGDPU9KIZW44
QfcCnCfF78mOTOgiSl1/3geqTGf+jbTq1snx8WDi6EY2LCDIzqfkiq4gevF+tl6TI4xeMYCh/CC3
RCvuZ1NabS60AJprSCaw44Zz7IEAvB5B/he0oFnNtLHFLtacwIm5vqedGAIYn+nfHICc0+/Sv2Ug
xw6g0zOEowbcsm6CPGlEDSP5ggGQ942Ko6fqxVDoBAm1lJYuJxas7NwpU3D89rK59S5jJW0bf/tR
sKDzAFT0YUN6jX2zXA7zyY1WRiD1dQxjPSgJf/tdxIoQtC+lj6bk0yEfa7SzlshvliN+bviWFJbO
znXqxMJ7nF0LTzJfrUgya9lqHRaAYtEYbRMWwkD+dV8WJWgy9ZVRnRtj+7SoYz0zPJkxeRibnTro
bRdUAnH2TgteZR8hDN+Mg/xEWZDgZym/g3OCwDQIAL0BTD3uFl3gQwKSsVMBMKXfJOJlpN+EbMif
56vjoaRmBbvtyUyZ04LAqlTYkzaG4lHBwc2BhqRaH8FguZxLL5p76JnBzTweZstzM/IpAcpL3yxh
Pw+hQgF4pOPwY2heSEMrXF8dQzGW+PmOTwyiO5HuPwzyRkR3sfLAmrCRF4PE+QnL8BL7wyWYO91o
R+kGIw9t1IfBh3+uWVTDey53kJnVp2hYN7SJrpwB/0OMAB6oOdfSoErNYI25dN59F2iP5uiBPHKV
whxtCGGqsNm/LzkyFJABX3jCbiS9hnI+kYB5qbxsZIkkiEsBcRjLL1ornbLMAQUjdkONx1GZFwqG
YXypkLWWootPj+aUdmgccClmp8v9Gk05DmZnoixqvhlsI8YKDeRrNXjXNFB3Rxz90NZr3gXtxHmz
qYSZjqgB4cYQsvAQ8ZaMzoLIDXr4ONaYgtg3AnlwOnrmWvyQN67mw1PKIewCzqr8SvTmnufKmpzk
FwdGitQ7oVUBqwffq+KjppUMItVCs7jQFSVpEIIh8gOCxzSYGV/9g2jYKAdUDAlFjbKzUeudyXr+
3jqFjcyIG7ujpj/jzrtPsPEPXgZnOB4JdQmQr+hEKFPxDtxiNsjOj4ryC89r4V5g8YwlGIGIMQu4
ygcENrF6ZHmpICfd8nHQ6YRwshZtOFXXv3W66NZ+46meHWFrCA9UsunsiJPpQRnFm5aPsTX45mGb
xqGQLpbXlu3QpB6FvK9OmXnW9c/AP5SjaEQs+4sJ9cvsX3ynM7OP1zDxaBX+ECK/AsnqnKRfiAqw
coklLVWtMS/xPHjC3ci+0/ChAHnAnZfwB/g4j1GQ6FZp8nagquoFqGkhPUiGVqBWDdIoL3Je92aE
3TBbNx2ZQXMgDIOig64veuSYMEnL+ZiWAfK5XpCM7IX09shWOhYxZCAFDGC0cc/2P1zXJpa/C2u3
g73DWdxvm4dbZ3wGoQik4Zi1T+NB+f7QozFNJHcxJPKBdACJkkBK8oFJmONlINqCd+5CrFDJVzVA
VYYhClzxTdiBVN7T+CF74bdMukSQu41xuIVgMg9fMdoFmaP8h1nS9UY9E/JGMWjot9fnd5VKI1EF
UMBI83Qp8eDsYYF2fkHyb/xqLZSgFn0hnDfPwJM+9TyQQvTu0anPhtQQ/5khfqXPS15u6Em3JZy6
/vjyHbMjn1zW44YID2suIfGwYTzAFWCYruOmNH7wU1uDMZRgKLf1nCHhcAjKVg6s5Gs1Oq2EGt9k
VYlqeTyO/wayv02iiYlmxhbCurp9hoVwm6jX8OAsuDG0t1ropmDW3FVfKs/cCPabJBqsOvJr3ZF2
sqVmCBwwzEmDalloOSuyWjvUJ6gKai+1pRuLqsiUafk0TnCkBiIQ58jc5W/LFGbRRDnyTzDAlv2q
so9wQ6ea87539M9HzvPMa/zYS7waWVO0x2mJ9f9xsD129f1Ew+qNIQXcvQdlHt53uxx/Thpl8m+m
YGSmGbOVFwzFqEvivJyfHu/z+Xnes5+HgKoqvr4Mkj+oQLUr/w43/CvWBHzvkv1rc0bBie6kBW0K
5Ue7r4VxocJNf3zHK+Lv5ER2QKnk5bkVlscuIxyksWKEXQJArlrhHlmwVGHWSGOUtWeE9Kzvo5Xz
whpbPHm3+DV+zyXtBCQ6Le6472CK2PIPp7A2rHBLqTxdVpyBxcbEvdTFk/nu5c/3dMk5fRH7+UtW
bcaH4Bm4M+w+xLFquOXyit8wWhS3uKUpvZT6+aYlQDMmZnDeia6YcNjt3HXryMTW0liTWy8qmhkA
fOqMa4A8c6b4feP0dIH0/k+LuKnDljtIWz8WvS2aNo+xo+Q2ph8DWkfQK3pT+sjz84rrlcmKZuJu
nY7fK9FxL0UYQdwMxn8pCybRwjUbT1v5W+51pTK8sXmbmbZon+ETZzbwpNst8rLkBkW/XM3zInGD
C1yPs7gzqpc2ffJOyUew19YyQ0evbZcFUiCHN+ZwU5NNlGLKBfKH94rL5BnJ6+tnLE678qidtnio
mnDsDKhJuyMX653bIchSs6qiQwcX6vTQVhWPOQun57/IOmkqjp0dNn4xRTNmqHrHjR36Jlq1S/kv
cbqX63vgvWexb1E+xRa4vyjP0LiBPTH0vsNW/A/qTaG+klJ/PKv7HZeTSAnxdzSNokONG2Nx9Fh/
cIvbIRhfENKCkHj/b2JIo4sBlYkE72n4E7ckmoypESJKhrvaB5wHsEcCb8P95HyLRotJw4nqzmBH
qUg2fsKK0vhrCHOYGvgTdFEweWCht2joVrBjLVxTV9f7/xnBxJX3D8Kg9RQRW4lIQtDVftGBBcno
H4o6wktJOCML0ov4NnpfxFn8q1fqUZCCg2Ts0lj8sRMTS+Dhw4eaRdO4zCTkkd16QiZuKsS9nKdN
Khn7RtOQhZDYBk/FYLvoCShypJGpRr9n6YdxH6fkcOIxKB6/eN0SYCgR9+D0+HPNRXu1EZ57EPll
u9q+ESs/yWwFJDApvprfGooUNSFh6GJwESX78DELoZmmL3YBlQugI8yY03HItKf0S1VJVH5fhf4x
7gSn/nRRD243M6xD0mvZrK/iMu3cpm6EF7NWtAXjUCa4zXIQ8Z5kwDODzj7R4YBmAQleqV+mPPjY
FF6kg54UnFBAou5vF0OmOY0yvzTfLa7OvaY0IU6DG5rIfjyCSSbqluZVVF8hWy7wqkgLZ5fWvPcy
rt3ZhC3iD4yR99clUK8qR9O4r+MQMVTuQ2DjdOPE7eLX3wd0j/RF1XKadmdtBHWKtbqA3dQyu6vX
mjyWtKwMUdD81kYd95iVjIustfEkgxnA6b3LlJXI49BrLztVnVSxrtuEPqjpTW7d0GIg2ZjISBwX
m3i0/ryWa0HHA2xKR22UyyZZ0GKWYOLTO5fi/7+fR4Pd2BagxGcZIjxmsdCv5K4VV+1rg4vDeCgy
3qfceHN7druK30BaXAjJOBfVDdJeHiIdQdOfg/hYVsIYHgQ8rw467YX56ffh/jqQq5DVizG1YLLD
bEk2d+Rii2cGEqFGwbNLCG+hdqL5WcFw9F4hlSzhkxTbyOVZF8OrY7gG3EbPpcIyu5QS8YOBcZxA
ztwC4lq50HUlc/snVThSPAJGUcCnqNgBAn84oMexI5SVclVkO/8qvMRQ1dIVm1dOStVBrBMm6YlW
niFWRCnrnLU5LsRc7OF+mttFZ8rMblPCGRFkT8MNyK3SyDofv0X0n5DWLfAwbZxyrIPyNu5T1Nx/
m6aExboQO/Qk59eB61xspH7As/3HUVSYm4UgK/hxsXzJD2cfixecSO6pATtaoNOVJEv7Eh38yaV+
7Qq+pT9ErfVeXEGMfOXhz2p/AGZSlhIEXH1nxaKyuCetnlel7hJjODr6T1ME4YEXWmf2zsPoHRWU
1r4/dSaToopyDpzmDy/YLLu5r9M15xR6FPtPe+sxmcv+5mkxFsrfXcS31jp71+iXVhjTv3yei3Kt
LGxflTYnet4DkpOf55qdfWNyzygjsGld8DcbxKX1LRQzm34kfqLSRKxn8+t8fyeMb/lkc4p8gTbB
eovsye/FI9szeclh+GgmyHzoGPprmpKh5w/ACFGw4AVtovmS52bKscPAB8r/8w3Y22T/JVbxbxhi
M9KiYCYg1UD1LXWVhpGnm/TMIhsfv9T5QYxCvNNrs/PvGEWZYmWmP9WXy9CCKFFuKuQ/MuT8e1l5
EeR9mi0Uy02K+TwomSYja1Ivs8Du7TgoBD1CUEqkguubIdBLAdpyKcKxwyUGOmXf4zKKc1/zyrne
SFuzeL2qykvwDJGSGvFpffyRLH8joMkshX+q7gXAJJBtHWeeWJfNHQLAQj2AQTGQOcWrh1RsBFiq
nYrO8JvMA/ZuyGBLvcwDBWNy9HC23OzF/FQf52d6MhwKFXx7hDx27shueRz2d8YYQVub4jRagdq8
nJnI2t4m4xemzrJb/SMFeHzEXjtJB/SZSlLzqJGHKfdt6iOuij7/FxOzURm3qSm7epy7L10n+BLf
DTEllUJANa9b6JZYpsLAnh8Ao2oLNd/EZ8S3xteqVZ7EXAS4rjXRuKNP7a2eSz000pTK+LMPMNEg
8zs3GbpAOFS+xhuF7FRTaCGV4i0Z5rXqKct4Igz5AbQQIHhMJtmH60PZdmFSS/LrVy5XcsUH5gTc
LTj3v1wYPNQOS5WdG3vuj7PwwmHx01dssVLnM+u3+wXxY2kbVyrrlPuQHl5o7CqQYqmsrweV2vSn
BISc7IukQbyheor5BJ+5hdUPUJ9djJUjKMOtJDBmPNlizT1r5SyzI3Og7AkGajUbUrUBdQPN6AXF
wTMIKhRQSTUCFNhIilkebglglyCehKGTLvUN/wSuswD04/CkMQPhDrdAPIXQ9w3TeRSQX/IZOgjP
q7Jw0yVHzDS9LnrPYinLa7/5s5lctvAUt81MIR33eLDEkrBDMF+EdOBAr/l453C7UxJP2aAQAdeu
rfzCbG5yoWHqvv6ELEfR9IAYLhzopf/llpk1o5qPVo8AinF4NR0+tdTMBvhoPHaVIuZyeXXRcKEC
L1ofdfElK8zHVPJTnGuLS+LiNGabvr8gWffuXkLfy1Ukh1uJuPv/y76BaNJtEguQ3QkAOfXflbhq
GlFbQjuSP/bSclS35YM2RsD9+9HZWX5do9Isue2t45RJIy/NgQOBUSEb81YN8RBkS2cZWo0Y//p/
+0hHGe25eZjAJqZgmzpkU0POcuVzaOOghAwzC1zhYFlUWownijU5pPJgmttKVtve1mreethn8LcY
z5CvztHALHQ6YYQUZH/RSwZEyNBOM+AA6hFh6QEoNFcebjPs/BPx7xIKdzVZXaFhmCoC7Kd+WSd/
jVw6FUuO748DPmFVwHrMHxs3nXm4UwCAi++M7XRO23yTO3/1BndUUxlYurSJ4SFzG6W+iNlQ2/to
EOyz1C/fYs5AiGW9L5jVjm053osKvdc0ovhR+tUq3pKFYTPvzRMu6wvcS9IcxhyPCntCSMTkutF+
Km9kFezZhEju4Gbvai/vSLfxAHeBpgvD6t5pTdnHFqGFjLZnOhJnvijuSnWb3qBzJbYpxbLdSL94
E629pSjAAVaKlSlOvxv12JzwTQLBqrW60P4MfRDFADBHl7osIQnMrAQljHDB4b830Ds8FkaZyW9x
kDnAAsPtY7K1ItF/3Me5ApHkPzUPdVGkPP9o3EDLHPp7xrHZmfZw/TLEmlONdLq9eGqBhUXlm/Zi
aQdidPLq8vCegZikFxONCd2Prh2+dTJ2gzZSGH2AqkgxgrMw5B31SjCs4Au+rWXDzmQZHfgnqzQe
unS20BmwL074R5IpfN5x6qldLw3t+W9A+2Wg47RWHcp5sFAWxCHuY7N86x0+7pPSBTf3m3N/CYam
MTHhS3qsiv3CLViGAlSVHZ8VSRJs/DuS40v5WjvoR9DstaljabLcwRDxLlZ2nMEkoTWeGcN8dRjh
rpcxNecORzcImHXBmFj0zHYNWXxJZQL8s84bTjcFUDC9aLGkzIPAvDvdupF9q/lFUZrHTi6PvEzR
JaCUXgPoOXCddi2gJHlcpqelqbD9YlrwmtTcwZA7BUWv0NS4gIpFkLW7WbcI/tBCs6sau1rkQRy3
0OyJlNRFcfrKbhyJbxfYUYjTLhd+TkAThf7sQD7Tk2qj3H6CuUamYPyhE6MCYEt/IOLWpUPxaPP8
UYQ40PPbTD7Zxc2Qphb/PRCPNO1f3BB0z4pskBWDMNlXMhSQ9UHXk5k0YZ8eNuoPbAeuWOyG/655
x1aY9QcYRnbe7tnDc/torFWF2SiF9Qyvu0IypxgfeyRowkwWE06/NVkwM04y8+IAVrMf76A4tGsO
hlePcUf0h/2v/5APaK6wF8nTQWoygpOnOJjzYNzaFLdFGSjhgwJzq9Rt1dYOHQyuiBn2pBdnihD/
NWEzUudq9qmTMEgDGbXw1xtRNUnteKUkemV2zBkByPZvVDQD0NOOvoZx5ODLzbnc5R1ra2gg0Wnf
gToB27gA2Khq8TSjQUuqW1chzGEzEqvMOqqFD+4YZB3Z7WNIH/hFmqDn+qB1fOUVKqlPfwoVYtMk
cyTh/POWr0Bk8JjASXqhKgY8RPCVQzIRH8HaR+SkfU1gaZLWLrEy3GvDhn0lf6svjlDLGbreXL33
srjAEHvfpWDMCnKTwOIpo+tjUiBI0igZZAHB0BowIocYuySg200zFO712f7wnkoQ60yccgmpC6gA
c/U54nT4c2ih7wvKZmiSUQqo76Yrzg7ymuITZnY5G5oyLx2ftp59yNKkeTk6RpxTr6QPKpiZ/ZSt
8uQfwhlUoudx/rLR28GSnc9CQ2mhJdqhOUzshBxBhvq/rW0UHxQM/xAO6Kju3ra07QNk+UGhusNH
oHM0q9q/q4H31NjNzW2HjzNy4nqvaZJsxB1HUFrzVuOvNtwU3rTl91HzKXYFQZygI30JRLxrDUXR
1KzKagdAf58Yvwil/3/VLdPyQq3GNqaIvyvgIlOiZIbRLZtjc8nEGu4khbWUmNusjVE4iuBLcxa8
oBIZDLgdPFF1MRd7q2fzP1ZMid+XoUqUTEvRyRBci2X8MX1Ahzwn2m84fFUVowBcjTg+ZxSl6LRC
t9/ND/sXLm9ptbRhJHvDpuBvux8B0M+FSwQa/qhiSEANOGT68XpRZkBRYBoO6FN1EzBD/aPI8Sz0
L/xc/uxJnQRhPiWWnaXnF6xqvLJBJZ490OFvJl6tR8CmWmn15zWd00FpigRsa4uOUnsPvOmVGAcp
mOu6ZNoDUywk8mypjBudlwBOEbPECreIk7Fh3sNrONMeOWSHd9FMsFKiPn61B8wPaQ67APsXXDoH
JiY8glMSVA1KjgSn4BCAGKvPfqNngOq83OEHLPQUmokohv1P+hE1917x0w5zobAw4Uc8OU14Ynzv
T536JVmmJEQe4hpncX3jQaNmm4PNvSGWnc1Mih0wME+g4kXs5kAPXv12xm1h0DW9djG1k8QtgNNk
rWL4WiWAjBEmLg2Da9fQQRceognS07hK0wdah0BR9OuYgZYE6VRi0ZCFZhVzbJNDCBQkD852dQXH
VMNnlrqu9P/WCWhEUcis1cYI1MLpFA6CLwjMhOSFnGQu+PoPdG2cf3AoRbi+/+HMXKfq7Cuqsekd
OHeqfCSMmT5oskOmNbuJEkckms3V8pVoUOJ0f0yNJ1uO84V9k7aF8NZ1jaJnFPk8AO0iY9oSPrJf
91hnOYv8MmKYbNrTGFJtJlMa7UGnjAUTTVu02xk7bX/uTOvji4HZtDEm0MgsUwh7JASXKWhUaz7p
EjY16ZkBI59eLPKMKdVXMObc67tUyvXHgW358I/W3tFERNVfW0HwrSPZXomPNTrM4fQgrtFeYp/I
J4LMaRy44WJI2ifIW89AmAYcmISjeZxl+d4wNbqBJoEZ6iCfP9gX3tufoCkeTm7DAVJdcOt5niIn
6LIJgpNOp6YSqjVg6gYEv5fixn+OBmB05P9WTuKzGEowSH0uQ12kml8r4jM5eCg08ttMdqQh396Q
RXr4UPCbGTuY1ZSxpnw/DpWRg6FRoVN9ju7cv+MJLkbFg5VPCyJhRl1/qcSwtUObyhRFZNtQKXgf
i51HRr8N6p5ayWevP/LVcr/ZiKhQNy/XpFk/bC2sIv1Av3IPwaBymPXFKn/Fvr94Lmz3nxQCOOb6
56zqIJ3yaZ+rgQfS6XZM1+67Fkb60cfyF8WrjQH1o9VUTCnfoLJtL5VDTWyOchNIV0L2YMDiw93l
lfgK4WH+JoUOO7ehLkXel0cZtU+PXlq9zGWPKFSatLecJjCLl87VKWniDwxyQYZsHnsxp64JsdlH
jkht5Lc9V0SIAYaHkNRcC5TjO1Z5yoFJok7ksMhWt0mBq5UKUduMBzCrDqS68eBA2PYaQN+ce8rm
nA+2rWkFz+AhHa5uRhkO3JgKOzbgKapYpBljSGZ4QMUN2Y+BBouZcxGJXQDt6HphkJ9N9jKRhFKx
L0WhjPAsthAtDUB5+tNKXPBn9V4anuUBLQOR3LrGQSHOzuujCGoeGA0xrK4DOpNGFRszYFXqv66+
uBidjLbVdYcEC3W5MxG7dy/JAHw8D5PFEsQwx6RhiMNvZPEBr1ZU+7T6wLSmHxGKvyZ3qvEuw8Lx
LodFVep+7z11+aidhJe6fbhT73vlMHf+UToe5ClVlAxsxpIMTGTWbqMufhT/BUBN+c1zeg9U2e1u
DUnV2LZb9k99IViH3kq8esj/83as1CYY4IEOyqyvoQYHojYY6rNe1bgc76zOhww19Ea1mP74eonJ
cuBYCa7cLL3nk6Z+Iv2vIB2SaKUhz6gBNydgnJvAleahHt2w5JcQK87DJx4bWVtRZukKTtIEYwb2
OWjEGESdFa5xqtiMHOPCtj44h71CGtFuj9znAPUMiDVdFWiZWxmqmELsvP0NtVImmjQTNS2CskJX
/jmW1LrZnAJPJ1zPaUN74v6n85AGKNhdMdIbbGOVLIWQO3nqgF2AQsoauciH83eGwW+odfOULQSM
2gNwbVjHAKCzATaEvdGmCG3wBXmhAWJQM42xXysu+vtPEfulPopA8MDu2HSp6dSk+KtJC8bUs0P7
pvX2EDIo1JxE2Heqd37DI2vTuESZ09PvI3oGChESm/TvEvBiV1EFkzTjljhxe0cll6xR2Lsp7eL6
4e8e0DZhnP+fDPWBEf8tErtKGraNv19OhqzDCc9Vby+yqiLVBrJDAO08HMH3hypmyiXIKoMBuKfT
T/qmxh2RvZSm0U+u4+ZOrERoXiwUifOQmL+8HBpV3f4aFmit8R1DHV3xhWsl/i+ypbNdRYUUSKGL
/jfD8yZ/9/IYtBTK9mz6QbxagCkrEYB0znBybAjiglLKkh1Dxjb3oucgWlSYeiqIMWbxBVM5hg8N
EoNZz8Uhs71LUOQMwQJoyRahLvkkma4JS7CmDDIbQMLOBllOmGt9I3C76vfMHxIE/P0XRsRzRllw
D4PEcWqNU8mxyXG98xK/6gxRRxOix4eZCM5Mdmj6Lhr5bKrd4HZe0LEIwR6rnLldFd0MYh32hDmA
0XjZwbua9m9V8gfZuZFZHR9G+j/4hqI82QMfIhxJg1thz3yuJRJTjbVJUddRb6malNdyf/PTEEF4
oLemw/AkH952nnmbyfKEgctS7uIjn/qO2F+ZCU81WLC9RJ2LPLcSs4nS6MmbT5rl3rKoFmXtW8SX
BxKdFddzBXgDZzFpsfQPGze1NVL0QTTMPs07iKKKnCOjZf70X+Xhl9Z+pSiDGvXVs1IpxoX2HOzU
vtyomxtLO8MxPVkhLFPdrt84nkJL4c3NE4fX7X0bmgIb/Sqbbko9ai6Pm9JnHzMFmJqeqSiEJG7f
L5mDtoyX9DspztfA3qrvqJ+rNWnC9kDS4AlRmqcVQQeAdQKGsGMXq3D+bMatOJrVoJ9jV9YwHUcE
xOrZUsacdeVSmx2quKZF847rlhZtoPYv6BmN0NiejsZ+BRTggRMaeVwC1Z5q9hhhb9+1X0MfJF4G
3lMfr0Akrsrj3iEtj9k81GE+7leENIV1UTI5ko3Z14rjbNnn5cbHoGLgQuKU5KwSqFjg2AlpaZ80
mqGUGovwO6ZlQDI2EEpUehsL8UaLvpsmRBpvXmT+aWDaOW8bptjvFOcnUeicnEDWBlV2kwJwcbZ2
u3jD8yFUaixFZpiYHbE9fsHa+QVtF5buEprDMWL6N/yYI9oD9CQNyImYD7K7sRKCK0W10lHyfw/3
vLJkSYNpoj6QaFt+JkU1Kv+fLy4FGOusI7R/ImGRieD1Jbr0jlSd/FZF9lNE2Yk6TXkn/kLIYmMg
VhkU71mU5PluQz03vimcFPPZzOLncZoCs8WvGD5IPNyTIxPb7swjp4Qxwaae22r5ARWc9/2VC1Ob
vG/uRiwL8EyazGdvWYcKiseT79S6H5o8x2tXDiI66UHOHo+gS63jMxeMvz1JIQBcroQOHKqxqzSq
EQRyq1FPXM+AJbyxnNpt7e5QJ1nlfUf8HNuIdfVKWTENQSdlkhojG3N5r7LUKnt8/4xPnJ77blej
AfdVhO/L+Sx2o44joPGQN0rRf/cWJHoIvUQU5QzNz2kJmRF5WpS8RNXiF2k615aVz24Ajgf6LdMt
48FeX666j9rMGIu1GUr0ozF047asbyNn/3CTYKYN9eEDnOqpowQ35BuOv6eFwwfDZyHZkV+hFKwj
McaiyjY6ofVDEULzcp8BbsUu+jz8ENyyj38mP84c0E27kpWh4zWZY8GiNY0mxC81eC7C/32a6CYm
Snu38KxNQ+NxzVF9SP06DrBFZGFw5Oe89TYiCWGtABJOq714mM60JUBeZ8OIOn+Sj6mbn246gIOH
pYx7F2nUJVolpSlTMnVymcwmQtkO6HSX0gnlsEql2v1e8PM1LiT02PM4o9i0fqM38BvZPGQXP7WA
dVZC5GMmVIYNnQaj3zTrjmEHiAfaCr+yjvgXvA0utrbrS119+gA8hCCaboCfSNXdNkHbR3+HGTu3
aBSo3ePIV9J8sJrDOrpmpx6xZX1RM+nTHohpZWtSMicZHSCI68Hb3lDqO/BSVu2La5qhp9OjGrLD
qEzEfwQJZDgyGZ0DXj2ryS/rETrXZxi3Wh9OPlvfES8CBLjTfCWG+cMG6pdIhNd33laqc6qC/buR
2UbyjA44A/bK55JEviuByUNF0izbjMAVulF+o+Z9yRTbnYab+s/E+PcKlwgU09v2dqjnHGMvV8Tp
zf7L/GODr/yde/b3/KeEGogT1y7XBvtDGtQL022cXkQIVHgmWp53eRfCWgK9zWYNgvd0yLoRpbF+
S2DKeiBwtLA5AH/lc8ud65/2/uS0qMOqVIkTgX3bkYwhcnX6dep4DPVX5WV9eWDH+K6LELv+Cyy3
RfuNk8SELncLTotFNIWsrhFlkZBOsWCUrOheEtD8Bfw7E/Ir8tbJz4XaQJ6CiJAJcdYLQAsTnrl8
njhu5YnR7YN23afzbHXDTWmQ+ShABZEGyAJohEvXOdGsAXBznXU6WzLMTe42F+UqmMu3mSFVbVMf
pS2Pz8Yc8AVWCMALKXSTck/mwCOrlZjUAbos/I3XCqZitCaOrthUmTi8pSSRn5/JDmn5R+gsV3e7
8oezZpKSSVbOdJsDn6NuE0XDSsSQ/iCi9NC7G+m3l7O11bFmekXhn17M0K8IDsvS0HagxZ3MsJjG
RMUoViLL8j+wedMUfFoj66JOlpinFqgrGtWSjIb8nYbtRGQi3kafTekC5ypRWwlHpuBhc+iIe5HF
C3v+b97FU3i+/ta0mbi7JZAAhT4OJE86e59+VUZhDq3MunW35S3NDYHaoYLRcedEsNCOwTc4i7BJ
yUeXPddhfEVqzAMCq1pN1jJZrTHZqUaS2intdnkwQi2MRevcAy5h8pdyivnBMRKzbosXTVixcEJX
GTGVyUORvV/RjnL5uu8ZQdz0bNNL0yagolOXzYg/tV19RwVdExi92ItMr0RHsBtpssZBStUz73Gs
L5U4Rzt1j+SsVsjbZJUhXq3zsav3XBhkClQ6ZEHvvRhrkgL/5KXm+VaG5HtRn01T0jU8krNsw4E0
OxBqH1AUtijSgMU3EJqGHNtXurymnJD1I3DrUJIIOoU1Q9hzV1PaE2wzKYIf1lwHZSfMICYRUpX6
W77zAa4DIWJN3DMCCno0UM7WBK03QZi8DTboXYIn8YTvo3JqbhFRxOU8vJ7sMXHmJ0G5A2YU5z+n
zhBZHoPNMS50riGi5oU/TgtQdpleou41oadUuyH+CC3krFC25QPftJdaf3nrPJnvooghr+I7MDNO
e7KJtOn0KktWm3n97YXGeX5FyvbAX+5CaMyXOpe2smWjWcQiBx76KesiKcAi4JC8TWZcmKGB8sN3
xS00DmQn9fGGlRlAkLO6OyWKnxnaw4cJWZ4LTO/xjnBYQZJrColRPIo9NmL3JQGerFhA0n4ECjTp
OFYI7jauB0a+JhdV6H15DLTXHA9r/M/GKTD44olsKbGVn9xTBnC+XA3Yp1lJzJL8WPvTEB7VVv9o
jk6BEr5QZmQQfGBH6nZaeKAv/1NG/7aZ3mZBVREBRsz/6Vkazajm8349nrmFzIgqThXRVeEezKZe
iQwj9dhMCKLf7N6gD6J47Hg8JMfFL4tLRVRg0xpO/UHKSpuNDkpfsS8TPvwVM+ziTchocdoT/VKu
cSBNeEgXHErqRDmgwBGtlf3QwnnRfHZoQ3LJh1k/Ze426kZm6gkHOtQgOCW1QxuGN2tRrGemTYiD
dIRvG7urXK6BJcYq+wGXK26D6rPw8oZwTpX5DSnU41vnF137L1yWDpk42ysbQoNQZdjAlzF0o9yG
ZzRLpy7LkCjGh5cBWMnkWARbVFxC/OpdROQyHwwnstXBfJPIGKctWpcTfWiKN20dADQSdGrKL6gp
R+h1hPV0Z73CqOYBgTsRVZHoBoMvn5XDdQRJKj6awgV81/7VsZJtekaRizu/o01wmD7sqSWcqnlS
ZUGm6qG44HpwHqaAlS0jmKULbwAsiB9tnRejvxu9BHbsJNSswb/2E/+g9qwhfX86CWPDUdZ1T8GV
eLPJkwh+UqsAbggSOVMK3kmQXEQH8Tjy6nueCAM4VTHFuq2PjtpXmIpuiEr/5pm7/4oaeBlgThxf
0R7lPbaTivDbGD7gVX4fRWRfG0wVg6rD7lJPQEBoMIBAcuuPHKNvZnilTjeSW3pJ14lyGH/W/+S9
TEd8dGR4k6y+parFBrrTy0Ocz/4Jyyj1FtY/FUbVDy7Wxj4CU+IAXq43XKr/Lw5AzE/c7YVigo1Q
E3beW8vFE4J5vFPSaSoU/cDDNVzmaqygTkYxV1SqDxykbTEI5j5T6kw3buSPrqs2TIQIfpTFdwtv
pRau/1731FdkoVkhN9M1fQw/slRWsD9bNFWv86S2Q+Ws3vVLwwLXGVdmVMOYJTX3N+6mEE2/AMxB
QYP4tBwOVIlFyzJX+bGmAJ9iugt0C0bw84jg+ckuR8Qwem/RKb6dEObndgyprQ86wHLVx31YXtGy
oYe3kUFynYtuCV4AOY4hQe5pUtI9ZCKVKECOBvwoE4OmYdWNl6nCK5+mSvZ6pzQ0euAM8OEOIfm0
ckQjnq4IzwgtycvjyQfkvKHFJ4SuNQPQ0eXcXSbCYSoKsuZiylXue2Y45pTOsxGVCCyVfoA1nUJS
ekOCjfNDD7Op9tW9cXWSxzvEG5WPvQ3F8qWbaxp2sWibB59CBJ8rapU/92+v2O1UYkQ1MY12IeSG
2RvoE3NoaVUWBlaNYqeITQGr3fvHlF2nGbA9oNKA876DMLaECmOM7CCSNGvdFc0C+QAr/pEG6MSr
KvvLdk0s+rBQOEriGpZlZcBOFRWkTGYKTgswM2couOrPX9AEnTq1F8HAfNnVEZMmbuYPSohT8MVR
pXUvxK6Gp07M9JSmlsHW1/xoFrXOo3olqsQdB9CGXKDuoa2MNvndTfUOU2qCcXn1mtWlT91SHPco
41IZyvdFe2SdKzaIIHqjpK4mWaXRz8NHPqUnzPiUcXdiBhkKfA2cF52o0mfaxP5D/5npJvxrRLjI
nz/JejL4t0NTuskYMq/VcisWdCoVobH2jBzbqJUVH1fE/qkO+8pB5q1jTulGti0zHTJUIbgUP4x5
8qF1c5IYDknQaSJnB4fgxmKpZlZo760b9mz5ZN2BZ8MvKpsJmV6r3Cz5kWCKdt5KLDiIE+wQ469T
sJgRvzvShSaTYyIehIIFd2ztoYI5VPli0HNkCRfAWqedGoovhdPqqIjsyrWZNlDa/bHBt63qnrry
NafquK274ey9dE0gd8/9Q1Q5vgEtpGquGV5NzjVOilC5Q4mWSpAxsAnEvJI4Y3UbFo2dmLANmj4m
ApT72yskJYJV/WbeJIQyODtOl6m1cmjwl4N0jQCc4n8XNgduGP1Z07DeN8QdIitUDz2tWM/R7tr5
9zpusLfwNbex/x1J4Fkl+o8b+0UOvX7mS3OPYtskpTcNtRTUqdi7NeiOb4V6jn1PEh525cu87LUx
NUmp8jAKbtvq9RBa6ao9iYT2ID7ZBanPrBWba1LUQc8LveIkphznkZapAxiryoswFBcDkXWs5z9O
7Sc1QP5D/NB9f5dVI+2ieAuvJuwLYzQymP5/Wy7dXyCtEQpG4JBnqhaZUEC06Cr0WuxQBPg1N2qc
5zSBIMtZ3iZMMzWFxq0tuQGW//RHV6AFdChs/O0rihJ/s3eOmbUW71Q0iuAXKHtrji3/s+Rd1Ri5
F5gfbd/GVwqbCk5uPL/RJLWRk/o/cju3TsVAYJ/uzP60lzuY5ZQ1LCUUHx2EkY4+YVpck9OSpFtA
H9YuoJ76bzL1RxX7sCFPh+SbvB3gJhPnyO70HJvnKWvkcGMe35WlWKM2XMjjZ53DKFlccQn3oPmh
Hptftr/sPTkZO7A/7H/0r2f9ptvHE8C5s6qzanfB1BGjqg7gg41EgcvK5sYzrNsUITZzgVQLOGqW
DP4HbyNhclylP5xE9H3IOktj6Ff3RjfZpKfeFVQREc8T+ev7UsKzKUVkTpaZlDL/fyQGhfYRX47K
4vH1VJdRMWISEKbDCH0VbCNQnYnURnGkbDlqxfu3IUI7Ynk9tG6n2vLRfTuVE0Q2I+TGDEUQonJd
87ao/OpOi6Bl88n7e/Du+CDjFDptFAuSqBotjyRolJNKXIJLwpzf8ya2onMA+xmpiMHeco8Z0EUJ
12CxvEGMe8XBv7gtIcrm+mzguCyWfqAGZp+jIipUT1+zgBu08WINMCu/zSUQhcUCNoTDMvRepyJe
DO1QmZ5MW6bt82zb0epCzLB+4GOU/YGpgy96/4DKidgP4xJ4Eu/eiTvZI91i8fr7pGBYvjjFPloQ
9afQyqCyiZ8H6TtU0L+GIQh+a13/jDVp3JGuYFBTB8UiAgpchjG68m3jUrnnMfaFo0Ua5SbHKTo1
7dVdAT1sl8JDpJ5KWbt3jJoPdPFIFaCFaKNXXNMqdcRCwyxoYH2XO655ux7Wpbxnmx0xy2lnBAHl
4UTy3TAfjVJil8HQf88o7FrNRT4NZ/ZgeLritkK5SpSxQAQrE8QOOUqq63XblGdtBD4bey3Nfdyt
YpSE9TnzP0PvCyHekwIzyZ60gIQDZi3k/pYBSY3svDPEnuXrkMrSYvXLzg5y0ZVSNiR56owp29cn
ZzYXuuiVno2Ck4rOJYNvYY8Al0BY8LPkeO59MJWjzRq9d8ziJfDtb/GQ4R47lTDwxCqqQ16ao2cl
6gVVzlxg2k12slsiM8fSUyP+be0b6oklEOLX18STG/K+IQM03A1wjnvkuRE2ZJrLKKuknTkvUhWc
X1NrSqBSli0Ot1eALwIF2XT2pIgJ7kxzQxAdltzh9Gz7ja/jZjJSATJo+dspre0i54yElSATfeoF
GHP3XguOkqlpsocHp0Lq29c8W5Mc75Xadu/oYt5ApXyKvRDbN68ircP1OHSnGyZy3JjrfCGc3MFc
VrEnK1+crzuBPzRDBi17drcrzKiQyvMZxZd2WpaKUf/HB96pGmuGZi+2kaWCWGFk2X9h8VYVdj9H
Fjes1RWR9ciXogrA8BZDYLeMIjFouTEGlSwSLkKDvmdOZhAGj9gIJ+tEgoHl3JrwT1tTB870r0Is
ATZYMAxu1yJdWxwKDU5FmoMtofFNL9fF3SNwFlBkLdKyzr157FtmnymNfkTaMbmrPhSByyMk+Dea
K6Jz3Y86HCru51U8DOrwvNYzuqayiypLDCtzHWQ9yzoV/Bpu8cRZ8RBnF35ynoKQvRWdg81OEYgJ
m2xG8kK0DXsFGi1WTt/7yZLqvJKPVjPb1QIrQa4QG1kwidS6ttezuKOtopihZ/jVQUSLDLTGXrZq
Oycy81mnE9qU3nhjFSM14t3fkyWMy+3EFtDGTLOWQRPi28rbodonKDuq8KKhcgxFuJbAYO6nGK9C
7Ar7IMTkCJ7kf7BZb2hDOd3fXi0duYQXlWJoxgZRc/pieQuKl30++P/cVSer7vpTRkiDAx9bBjww
vslc8I+ArHGjA+8Wd8dqFxISqWXmasGQUz9SyMG0421qRYDjj7IzHFfhIAHWpgLQeNQV4WkdH1bJ
DDROXHaGeUkTieT2MA0FDMmW6eDXMVAPHfZdFpFNp36veDkG+JgkDr/D6JXFbzEU8v5XYK92FGiW
Z+BCAthIsX86RtjJmV6T0QyYkJIRZP8x+fbMBAN5m3QhBKpy8ZyuRwoW+1Sv/frKXYgM017bKZ/I
0ekO1vFe3zEl13pNbHq3kpWzxPmaPAoFcm6rkHEWtjAPtsC9R42QSvUE1pDgmM06yP1TGcKy8y4s
74zM+ZQ2txkZqhu9FLf+QTuIoIVlock6WiAK/Eay0UCSL/+za6NXqvZstL6PtBFzTgXkqubj+v/l
RexFo8qVTiSvv1d2hvNwt/IKh+ZNerzejpqb7EyW824ZFxCGIjAZjvF7CfCdaunrkstseNtU0uZT
oqCOoxAMYEISNjRnFg4ggS4tB69TatOu5Y9wW9wEl81UqoASIhw0DHJHdNXxXnAYk/Y29qEFXMAh
BU1/NsdOAFZpwhkSdxQko0HMMVM+Ny7UWijBVP//9p4GfbzRrts+dfNuvYLJLtdFy04zFn+0mVwf
N4igFeRQZnmLJe3m50dec2FPNw7J1IN7PRbVz7a6ZA7YnyRUySCH4FgTr/39dHxNRw9j4BPQ+cTX
FCdWSTuZ0JXjAhAGwFjQ6EZWd4PzMnd07tlvlwcMEag2hv0X2gmbKyBTUyvxgcyCs0r9nhw3ZcKP
JsVMsYm7XpYMtpzd6E18K+5SswYJ2MDSbHKmC4KXq3XLxZq6pa2a1gdHodiobLao3vB75ywjjrNu
WXTjMKOSqMiayt8+S7aSVU43E4KDahJ7c/ZZ8WkpOAePIDOprWaZ2LxV/zNeAyioA+Jca9kdhHLD
Ve51ILb0ptUBULmZsv30ux3E1i2BfsZyCa1A2NsfeJ5CuufJdq8hOjbakPiNWpb6NWv440uptWpq
CLH3D1GvaloHrM+bNrdafLui3VsuVJ+vWST+j8LQyLmTR86l6kLtpsBAIXBek56m9J3wHZSyxNwR
3NNf0qNipEPqiwMQg6ZoTps3WNWF18J5yF6T9XbHkJeL8jLJXVt5mBkzXdofhZUoX8accd5kthOu
8nOJHiblKsq+RE8nMV8xGu4EJhF3LXgKCuXadSM3uRI17Z4hm0jEq7cr3g3nSu4G8SNL5/EnPajU
rWGl/Cx703K3/me7l+iT7YkwA7u3Fk/WG/tvtlo7XLek9YcBOjI18y4GR+v3v3TOqTFNwRXHuEjF
unlkGte0Kk/14V9aMA+cMOsL9zom4zVrA9xSH204PNHdf1LV3WQdu0avXF/iPrpkr2xlsg9woAoL
l+MW4KrLfUhhQ7CrzMquhk6w678P+8PadBaEsFGoWSDsToheP8ZYmOHrs8QxHl7WdehezhxHrPI9
lIHAXwe5zh/c4TSWDIPlgXcZjP+4Nu2l8hAIWzHu1Wo72O2NwCQguDU8TqFoGtJ6J4XBIWnk9zsw
JaPXAnCEIplK4KoIaauQML8iOK1lCvHfL2f5QI8bDVVanAfZT2hTcT6kf3qyn4xZPPyY7mb0XEIR
Q1wuSz+tcYMAemuQy0oox0j006ry23hnufArfytzPoFEDr63sfdR9i7XdrUXhQ5KPr9tc2wdkd6o
b6woxSxFFEoWdVgKFOGwrNiV4NL3d232zQ4xmS35N1qLAlGGJmP85oOYEsa8uyIDsFv5PNx/8cnU
mgj1NkdXzxqmYnTVWjPle9qY3ZjC54qwDw6IgoCV3IfHSTl+VWKe74YbS7ta2CfkMrXxPgiNgSon
+5gaOX6pyj9YRShU5gUZtk5cX9f0FsxxMUcA6pvBXzE3Ogwy6QCxMYPPoZNlMdf2JvPzFfv3BqIG
StWTFtquFJf8f4RNawLxtegHIn8ezaXC+ZIJs/7uKvI7EqZiY2GJgFNxDi0Ah5tbplX8adZ6+6uZ
b1eJJRyjORVxahpmMw8eUqzYd0VNChe7Omxm6LKdiT8YZRouLZDQHWV50mml7dT0cMbdA7ap2XTd
gIb827gyUdZg9AUbcgNDBUC3v1GvdIFE5kLjsMqI+S1hXUuem9UngwCJ+/0pW3Nk9sOeuPx92ILT
lzgRgXdqm+8/X2hHh7+hr377UgfduGl1sqWyYTlyjnicwkmd8HcnxdQckTcWbpiEF8Lnqr+jOi6V
NQ4RZfWeUkSji9TapHHjyL/evdzM6Kj+p61/o+bmSQNEkR91Fyx7RS4NyTU1nMbJPvzTZLYmAjo1
kl4RfB5PWOpTRcgULtd4E74gHB1omEmifDNL8qElVuy5tAAa/5EDgRnvEMcYdhZgIHTBvPScR8n9
j/+6j0oS+aSPFsLCBnrkXFZ09j68ObEPDQGhPMJHsgiik0afld9rBrlBBeXgqV6wTQ38AqsTCeqF
6TL2+PecspVvakocjksE2SJsnay5k2qy4skx4IgIgM57vNzZoHcHK0Uc6T/NadwWRSYT9V91VwNS
+PWIGf8eKlfruzlLRqqb7Zwdr6k0lEUUTUBE6IweC2hgeXMpaiuBRO/RoErBBuTmzVQsI3EzOWfw
PTALARP3V1rqyoa68y/iC7llflzPe/MhGSUYzossmSOAFnNf6BOlFgBvZusFtIGWg/gXT5BfvOxP
DeeR1jXynNH3sEtvO0zXdpjRJ6lhmh/d7AnGJbNj0YPjvyJU4AKe/7Xa/s1UTXBQmPBxkInBAR6b
hbNSmlEVnD8lHOJjdDMEZbo32ECUGWQFlNCPFFT6DhAnNB2zHe+ARCtdvnQmFAWAp+/BTFiUPaby
zB2bYb9sI6v+KzLuJ4/oVUUCaLxN6LV8OAb0m9uv1FLx5ExGDaQIHhAtjPZ8mP2r69NGFcmWW15G
etOz3v31iYyc6FyFEpTE3TkXNj8hS+zreK8l4JskoeK4WbqxG3mKD95CP1tq/6nn+/h+bN91kPTT
ED1xoo1pzB/WTwIvUiDWlEr9Pk/CRDo2rvqz/laX1Ox8a1f5mND+1Wn8I3tfHaF4VlAKQiNNBHT6
gEM6wQtY41551IDDRyOA1pY5zBhkxUjPPBXWo5LEAHKhsEaLTMVFWxPSn4niWvFFqpWrLSV7FELW
spWo8ldaNIPQEXmumuLkJrUQqsij3Y8T5AukU85CFo2zGHDwgrNrpX7I2EVcetaLcE57odGIofZY
GUkAf5Rw/xCoWKhFeBzx81Sid4bMhbcbQSHY5hwT2qLi2i9w25N6u6DTn57zpf6OX/MAovaY7wwk
izUbS13U8zP0M5lEmVYZ8W6eFAcUK0anvOgNdvFepIEIxQIa0Aq0h5l+CM1wSg2T+Kz+8wveEqrG
fQT2oFGNaKNixhBNg2i6yOKQ5LMLsesG3mWwOMuwmRFNpjX53NV8pWncuuRdLg1uEJtk3R7D1zud
ZE5pw55+oxWkKNUK0D6+/aSmx+jo5D4Vbl64jMaXpUJayLVFxAOFfB81sXtDgA7sHDToXrIXkscw
y0oBBNBi7pWTt6RGkhAibF/CQOTgpYe99C30fdq4k788p3r6SKdeMzqAxTf1b3fmSr+2xMPQp1ox
EudxZmHXZ6Ny9ce9MIr2g2ZpHfyrKevb51BB7Jh6VPmHaNrDDqHGlXgvoKxX1555Wm1k/L9OnXIh
qB8RZkxBxoDQc8dI9kGzxyEHjwAS0PpyuktwnKazLCx97uNb9ZXiHk1cXSFdRY+DuLPSbZ7Ayv1t
8ySSl9k5mtYzXWD2IZ9zhfNVgzUEUOV0DkwThX1qlvK7iYoZ5wRMhzQ/Y8ZUvkqPKh4oymH2bE7w
ojSpe5ZsM/+c62cAOz6laQYP4p+GqjCDePhUE2fGh7Xp04tkuAYd+jIY8rPyD0uZgC9AmlG+ZGe8
bpux/P8BxcapSBy3vKdLQ6rU/SXNv7v2DN/QtZfGZf4xATSsI8iqdgK3e1SFYckOEAydpWGxbUvp
sn2M5/G/P6g1tKVEkpry+isaqMBR3ofhJLUjkmJbbyVmafL71/U8q41viWS+LsdJQBJxogmh4JwJ
pxzkL6MExZz5+8v+7y/6spvjqOQ4Vg8o9CHmY+uiBJs3uAqJ14gHibEPqT1av5BfpyvLXLI5CBqk
s4V7uu34tP33aHDjiqEyRO6X2QNKsUpzd4Gm9hbQ7hhR0F0w392FLc9KM37LvT9d+YG9CKCo0tM+
/rJE0hIkGARvjTum316TYYkdE3aB/r79Dx7yf6pidUkL1Z+eFBNzkOsR1716geKZwIQ14IHlupyp
wsKx36cu1yexiuvaDY8XAnfSegFVC+IA26ewEazy7lKiEe1ptZ3xZBXr5MbZBQ60d5Pa+1Yfs5U1
rcLL9AnukiMlOuB3da4x0kRzLCuemRRwJ2med2b5d1DuOnZAbPvpjWp1nz3EwzNeHCYEQ5LCKBL0
RKc0grBGhw20cnvl81+0HQJMT/efaTYO76onN2Z7BHK/r0GZX/IzGk201NLnXJfkgNcsyHTxvFA0
dBjlOIFxniEc6wJC93AqLMgOSwu9kazN0rD/8m27vHEa9/w+FISWOQWO2j0S2wIWUlbU5mhlMEGb
1aaejtf9Gi6HXu7IuqgHmHseKoL6x4BVSryPIAJKCgCfyQLtmgpgZi/XGXjiBiz9+l9vPGyfskNr
4gyhTFLKm4XMppgMB7y20lm2bB8zZPpm0Gem2dHzNa4c1F0CBdlCTR9xBeIxDZGJhI1WZ0ciLQvy
lhDB04ZwWqCNK+TOtmFTDy+2oxSkrpE2YNiDXWdIsTTkWGbmxpbXWi4G0cswcYRE8ZZNs2ARFNMi
ZLUvVCehrxTw3O67RRHE1A/pEwq+qa1PPKiwhp4H0Oj+Gj1KNLYGChwCYbvszUNICuBnhWdJehpR
q/XmAo40FvlmovweVAw42hZYR71x+2VeE/7IGSqs7/zvPIhg9q7c5fOTM2I+p8+O6QJRu3tv+nl/
ap2uJyWkb5ZnPJ1ZRlQcGAJ4MnDRDcVEC8zQmTYiZUNtM6JCzNVbqdGFSKLFnAF7YOFFJ/5omsZL
0CPP7obPIVx4n0A6QMjuZj28WLYOSu/NdrO0xX3pA6gUwJAXi1w6DfHdG/UCX+ef4AIdfbDPFYLz
EhkQgHUrtbKK6arFLDiSqIyJ6pDOVWV4k70nxLliH0ACQTM1Ojio/yVqImioJ9ahofM0SNUUtqzF
9orOs5/vzdVl5BIpDisMjObp9nf3cBUw8UFAB1FYCa63FkJQURjwDgE+slCKgU1l7CzDo/34BotK
/xBdvcko4gMlfrV7gUwJxrJZWTsvU2PArmEriam0NDmutg20eFid6n8sPXFfew9eifNN8DF5Lcu1
ND4pJQAMdC6mHm6QTOBnzDhSKCVN5xSdd58S32IRFGWa1Fbw+oauXybIOJR0hmSvwWBUxlg/qylw
GK0c7prycr0f4rKWILZLcrM4kKCRKX/UqjmFnRxFWXKCgZvgyWrnEBSRl6x3KEioI4hDpFEMLgWI
7LGRgoiPThpjijd4Rek6PB+kZ4kSwkW1rMYveyft4JZ3V7h9kmBDbmoypEoR7uHwLgO9lELnU5jF
ZleiZ2Zl9SBPZtYu7rJ78hTZK5k5dm7PxFT3gkoTfMqGJpdMYWTduzenQUx3eXgzrrgXPTjrY8Jq
OvHE+x68+c20cmFiqcWpb6JoOg9wsyekD2569FZ3bAptot58wdS1BnaEHas58lJ550FgT3MgPoT/
wMpfH7vYNloCaW24HOD1oSM7aIBbf1BCG/cmHYJLSl3KT38YZusLaFZA1NdrGzg7dDdDmrFAjbDe
sFvpsBodCKgG6kSqNyKRIqa9mMh1hTxNaP2o1Zr5Jr5zanQf7DBwO+W7LHNHvPTzBEJUwImN4Wj7
7vJjNk1jAHNf1dnud39A2B7e8eLxPFQnP9MFz1nnrXqNqVDh6Ko+Qm6Qj9uvxskbH8vdafgRQmLb
2r2obhatwBtF8+gfPb0EnwQfdH3Sif6Lkugfm6Hg/tEbKo6Mrn1pYS5/fKV7PCNORc/4cjibdkfI
B77x9cDPP06mWcO7SYOUcF11wK+7j1DiuZmNq2AmkXW5Kquuhiri1PENVF41WytuBzhQonY8NI5T
WpAJr+H+MbQMB+AWDfnXggrkZ38MueB5D2p+VUKyIQd8GsxA1O8HVlejrGMsCFuGHpLYwOP3BMKr
i5fKBXm4P59CszmEwHjyS+eN0QbqvwprGdT3fu1gk0yryjz3e/JL2jHIGruBSRdFyB+FMZh2HGZd
oL0luZVHzP1FEXmt/wAMV2/RleR6KIQFiW0xAAQ6iBGC6sbhKuud5GoD6tlT5UCQ+NIbt0+l7uTu
9I3VVubZ1Bt04lDSxHcOX+2ZHRu7MN5Kq1IOHmCeFhrkJjx/t+GJyZ62gbgOLDx+Ec1StCPZVlqG
JfPj4ndfl/6GvqCCIn7b2blmzQdu6qhG3QHdsf+S/j4eGhY81lJqJGR+v2zhyN9SgyLbYM0/JCmT
ms+RkmASt0eSmM+Pd6IVPxEZ+GExx+QlpQKX1/bcRJXCx+CH+Ikun8gAmxP5zHF5xB88QCdgrrg5
os1Ra7///clFMPJaWZRH9ty4foJbN8wenZLvrrv3USkfAjcWYp0MFEREQykb6FRGNdeWCT/RjYYP
7mEqlj/kw5er0RMdzY6R9ZV8F/rhlFR+wj+dLwsiq9ZlhcUJcbsS6k3ShqKB+iOpYOpbh/FutfqU
OlFC3KaBZggze1phnMrNvQWV5TdfHBhuybrYg3oZCNg/3X2T+/+cdF+3NMa/6FVThvRuhuIuOL4S
utXf1LPcA5QgsbjmPh9GmlEJK7eXRJ8ntc0YhlKg7uMvPJWNEMHUTewlq3apGF+hNmUoQg99FYUM
5UG1QAmIaxbQ9Z3iLqLQ31fDtROuSpX3Y6EZcCYD9yoJdzj09GFKD60Csi7CLfxnf8e0iK0WpiZ3
kLdxPSOU+vEKPm88dP0fxW2wlvoqY9tymzuqAfrUklE2sMo0N+B54dU5d6J0o4wrJwLhfuT2F2MA
nkzv6lQuxEg7Vc3AXlUOMKp23KWJncXqIRLaPgcz3zqcYPjEcuwCpZPoBwSPg/HeWA6rf5sktpsM
9LmdnOkl5VW6A2qVj9kvyXIMTvaY1UFJyfqwVNck6ffiWzi0CN7SALKxmK/0yQDGZVeChl08m1YR
4sl0n0nXxiTtWaD2Cper5FzQr8fYLGV9pawSaRo+m1NHCcFC5gM7RarqXF0B/wncDGmF57mCIIn+
pPwfvOwgXAD7sSL5XU7xqPr0jcQXdNDxyUi51IwsUfxHcigqyTdhfcyIUK4hD0D9BGOAH0rcF4kZ
W8+Vr2kHRc/PeSvat5KkpMwwKPyWQ7n69q9r5YZ4ONhMIUF9EWfTS76kOgf0+K3xg78UAWPljEkG
dnBXtafQVmnxZd5ukn1z0Ck9QNjtolmOS/eMptmSdVVLRKwZ3rbnTbFjdz3ZmIIzAigjRIGHJEoT
7S2uzvBQge+YvZYv7PbEA+H/M8N+kFTb3sm3xYRlwytPx4zhgqSkxWJtg/52cPNaE6qWnoZD4xgU
GffL9gAqU3Itk1vkwSJNVljuwsiNj2wQ95B4VgraYytLV3gCdkEX7iEDZXRD3duLYsoOpn3nSIPZ
q9WrgXUVdpKEn1/B2ig7V7lnbTrLrSKwwTZLrzhmdCHSxRgttCTVy4dPVrgubWZRid2cqzp7Tvfl
lC7llBeWaPkKDUoKjWcDXMiDRhw0eiUgKM0exsSkHY78Z2icorASQO0tya0axf858903Eb6PLpHh
sWtAJQzPw6H2PwgrsgmEfAG02TCMkJ8MxXWe2wQXa1Z708rfdRJNhZNvmATtbs61BMNrsI9GmLOi
IB91HXGxy2Ctd/Kee9EFtZ0k/e6oMpXWbm1Ncdk24KOMlMbB9dRUM7I53xRlAhOXaWCEfGQDvshc
9JFuPxJ71gniMVUt9FtdzcP24GoywQqjEOOvNhnbRaNDS+uTYph+lj0Yd8X67roSh+pykiHTVoyS
tNcnjoRaXWVFOtZNavQ3oSqVEriS8KRwyS5rESVI8C3Ol4uzmYmdKeLisDt7y1+jnPlLbkc0YzAF
sL++S/EHhZiiixzURo0cb/aWBE57wu+gDpkuU3nyMiJ9sQumvr/kZex+Atqh0P583GjeNWfl2rF6
DbUHnk5GVpXzMYqMfVoL21D1/apeUXKIkYBTf+hGwgWxdHoCAiu5VeHsrMahYg9HVFqxbd8MoQtU
zZbBNXRLvLvWGU+4b+MhBfvCzCZRu2NaOM5OUW1AS2S8jJqQpko3w6XfQEkWdDxhml+GAXQlRU/R
zmbnuROO3gAkb9X5gZnwXOpyo1UrogOMPXVf/X/Tw5rqJ282SE++VL/YW6xTlaiaChu4Eb/WWGJ4
htWeVh/j0gBHkJlLPSKYJ5Jq3NBHj7BcEvFE6Hz55H/L/ywzJ2Lduql55qwEVDOzy26HIa5U0aW3
TGoo7jWRR50YEesnvZp0lUv2u0e8a+tIA/KZu5IZAlRtucQ6eZ1oE/x0rPCuRPanU53ixLvrYNBO
WGq7l+zMZgxdGDl93b8n1By/8H6RETNivdOOVfn4dyiDi5wdKFEd3/97vNhxnUxmzG4SP+JwljT2
thZTDtIqrN4kVHHNf6FT6XcS+0UrxLdp4QzvptvL2mpPAJ4lakS5Ja54s1iTQilvRpel6aMN4yqg
O60M9vcW91ii2LlQSrVfxgx0hP6y+umz3Engu2fRHMhqjLikkrpp7LjF0Pb7tVoD44CklfgPlDpD
v+jK2arAUY3en7fWbKKp2HxQZeHUHqLq9vLBe3xEd/ItvYWgIznV82scj9m4oNT5KD6KrhzWuXrJ
0ggCwNhIXkk2aBwolNX/yVFpci6YlWNcKeRo3y5MrNtPsqvwTq8pvKvntd05x+KTfXdf8BFXZBCa
4XyNNFWrm4mQ0tGoWkTuE4pWmTAMqp2AYme89C8FuE7TXQvK4XA8uGIWTIA9YM7bK2s5gFHYDwOl
qgi2JhWhve6WTMGTb1RcJ2DtLsbOHWjFDiR/OThLZJi1ztlv6IBAWcYCiOJJ19IHD5xBYzgVBIoT
VBv6oWGFW0R+iPRrHW9DsqzHbE9wxUctabNrDGcVFDnlMEfRTKGMTGsQ1BV/JuzvL5MG3WIXV9e7
6RdjUPTKlcupDfT4OdmvKH3uqG/D3sAIeEJmT8PD8i06Na90uIzBK1Cidl2ciya+52yVla/TJG8s
u5sJzj/Toqz3LBZUdEmgdQlz9vjAuSDAldhdgVvaJkUR6cb0K+Ldb9lnpg3nllFBJOo0zWHAQJ3Y
SA0n1UmAP3yrPjxTFzx1nNygMmuw1VaAgOSTZQn3u7oIy8pe1Ae3qBwcWdmzPjn4zIMcAloOmDTQ
ktJuRDR0x6qKiJ7nZ8LB+0Lm8jPQWIhWeSKMTszWWh6dDPZB4YfVSGQSxzsh5HuAzwWb4p1nuSa3
i7clE7q9CAkfp7/gbu5oShUGcPsYqEO3WIxww/gYGK880LptSw7Q6FWhPgmVXLKGTsBoj5E9WkJv
3uKeFEtpj3Sjs/HNn8XPNbxXs7G8H8OZdJ5GTv3ygcXRzw/iFJlEys5xmMvBB9d3N28iwC3mYH44
HSiwuYIk9IXneZxtTEOY1dug2A229QwW3YUdfIR6sl+yc0D6CnLfzj3mGrze3eLoWjzLYjqrEJX0
WolDuZ7teWl7ikpn5K73VtU9Ex2+WTv4wFn95NErtMxQMeDYS4HTCepRJKLGOM+8j8/U4JzAJ03Y
dvop8UGfy56zwCFMSQnK8TqDOcbFLkFeA50WL81lnuuh0q5Ysjutc3693juIQZ1abSV/4qBfs427
TIT3okGKiutA6jCB0heL+7gFba+9jWju3c/6UzGGYaaP0xoEH3c4U0tfnFmQraZysyl1FkAeqDTE
KtCD9MIqf9Va0b6C1RcEIThGVb74GZvTpTco3dsFBq099pJDRFFwkcf/N/OwY/4cTeivUs0HMNuq
l1dzWAMFmBG74Q5OnCQ+6iglCSa6Okljuje9O17AcDfShzFj7oaNrfWXZcOGqz3BTAeJoZooerCb
NNKbJvvG0pE2e1KHVlRb2kIneW0LraXhferJ2zn5PiwzgSbRkiezqqHKEJpQWmWsTGGfONIIgp7z
BpeNpzF+28Xke5lVFP6Ad8lJZuqGTFXQ9H6zmha/5oj/dHErEBt0urdLpwtKH19wjFfQi8rMlcyC
RO4ziqh93MP//1PgM0V+QRuFcObWo7LmDMGM5iXzky6J2QwKMHFg/MO1Gdn8g6qOqlIRpXh4OSp1
VcMUr0L6hrSlUXg0wNk4XpvF/dAIJbmVHsl+FOthW3aAkF5IZdmYopuejCmvwvBwba59IAUAaFCp
ComDnvwWMgguODyJUR8Oqw0eeJkR6/9PzLEoXfAIJQJ55oSIsZYAS4YyN+Po5u94wYJrVIMhARtr
js9oVxNz71XoXbb4DHs7MaNLyCbYqxAHfPEt4lapJwsQTGlU0GAKeirpl/hSW/9G67EP6xVzAMLB
vRpr0PUyiUvOdQ5MXTL7+zExtUYbJOhnwmgamsEcivATSeNMTag21O4twcDhUvW5KuwIcHnZ7R0b
9x2UeGAzR16fbE+tcIVUvOyb3gdgMgvpnkG9WKJ8NCH2GqBUuDdzFT48jrEdzj2d2uQ/Ykva5982
Epxgsq1t0s0PxcJCLeNFwxBBO2eY6cWvHbVc+sQMlPuUNWRavQUJ7Wd0hlGkUzEUrIj5pXaYSsSC
ZNqrERZ/eLj9KNbgeh5twy4Ou1F39HHYLqyTSfGWI4tvcx+XCKtOqubaf0arG931G7YhfSxHRUPM
wObz5I7k4kskSGAO8YDlUaphtqY9QGkqDIT0+uo9CMOAqDlFnTJs2CFX42/xL+nuK1VRG23OEMok
LcOG1zxQ5DXIHKmm/OWnVXBVaGU49LQuyNGXPOfBAsKBgkauIsxe9X3M7dyaY3ZrW+y9IjJI3bJG
PiJqt7ZP013H41XabpvT6et4MOF3qCTiKx3vgOHpMVC89gazdlbhlV/dEgYQqBqjXzzbc+TUNSGu
yXwmL7o9dqPhh1kxFIB13UXSkcco/9+6+3HLHoylf1M72fN7b3BSS5d/ReAo3WJtsjfA1w5yeXvG
44500yNGF8w3aNu1D64LEfWqHsT0yoZ0EpVxN8Paeq734VQvH/LgCRNLAP5zQ3BAwYYJUgWcjHr0
JGzAsg36d6+vjfJL5lW3ymgTZuo0NK7pT+CJ1qj2BtW8ZGxhj/904H2YY4UfwtZw82Q/vYSEk2jI
GAuE6jODg5FTGr0v6SolmBUkpitpWXIlaW4Jsbr7hzUvLbpSKv3tzkAxC39hSHfH5HtJtMFYyIVs
yQaSUxAPLjtBPFx/XkDVkuUspTwGj8GysQdA8cWkWZ8DddvQNagCVqjNXZMx81wt1SzYCBgeQ7p2
kQQIBp7Ht/GmJ/xxsgTFT1Qmbomlmo8HUoqtpp15n6jHqwxZcmY//fhy9WsXdz9RaH430rKbtA/k
STNqLmXpyRuVK6wFhpaQC9enFAaYA6W6T1ipQDZvvAoE+y16HzrrUP28ZXxW5HKwQ/sFmXWidNFr
x/IMPAqcTceIbxjS7QiawnnEbp+5yOkVti3FBqqucE1lEnrOOwf/yJq9QMjZ8/+9WMP5KbvDep3o
kLUyGO5yfHiSTVUkF5OpVtjCeiqTH2Ty+HXogrml6UCu9W47fzAh8b6woU9rpUH7VM0eEBhHHeOt
8I5Tv1HH24+Jie1/qkMa2+F2ZFAYtGh1+Qqf2PV2eSA6OXXsqlZZk+vxU+IbnrCD7opchdGjOHdh
atewSFbBT+liNmz5hR3Xy9xXXQ2GQg7g+XAUWC/DuxYrY3Rp3CzRAzdw1jYwhDF0DfrzGEfeM8CQ
2Hn5KADbDd0vc7JQ3NHSpo1D8/bdYxMiDsjWTnR+FMJ2c8rRcNep6RYVH5ZaNSqplV2uV61hpM7a
0kQs8QjibXhjwFndsq1S/QBw3uYul0UoYRuLVhY63Ud/DGau6T+OFDyFgWrDujKVrCFwfbELfe+z
tOf4gtEMH6TFyaGwqiWgRWeCC1JkAVAUA3V+J+TNCe+x+O55qBEicZ4O0dOmFNdfG+mYnFxuPLy7
P5FC6KIH1y0cD9xTg5wlFHTIlxDq3VmCUns9M87/A4kaq99amH1gL8wjpLjtz5gu7Ip6URb5D/ca
Zwr4IxIvaSeXRZJfMGprz90i6RxdvsFGGL/IqvbjXQZYCOZ4qxNzhBF2SLVUFCySRl/FVJNCvdHC
EWWvLor6LWufkrt5srLo+LPVwlmVeGgPo5daD9pydvF5fZaAxaRtrTZROE1VGOVqDwglo0ehC57p
buokkixyKqOvhl4AlGS7YBhG+XbiXBlLiqGmfFkt46/SCS/QROXvhPjqt+4NihFyUOoTMDi5Qfuq
1hkidfdIZk78qg5y8u5Sefc7GgwdxV1D487WzOECXtTbwUstyKLbHDrQqmu+aRGzUInM2rh7XUng
lBsy8fZPgLWmE+5oax3vhqOZ5zTnGQAuvg9d+qq9oq6C8PrOFls4OCu2FEhFHRDfzk2sgfCnRyc+
uRTGfEPSfjnLeerOi5DyMXnL2ePIwMKiJhyDHOSD8cmmd4HHt8dc8Hwesb+1AC5syAdFVJT++UdJ
FdmGOpPAbYjduek+B5vCndLmnhjkb2OY/3Mi6ehK+Br0WgVDfExA3cD+1ZGtfWuW0gJo2Ok5Vlhi
UpX2V4Riz8QYC63ILaC4dM/4NGN03aKd+SJVUElX+iKqJBgbQZ+/xFxUMuGmDdCdITIVPwkV7CM0
MXUjnEoJbzv7ybcq2FRJW6hqE0mHx5ut9sybhnYVgkfiSd9rzgo3wgzg5YR30/V2AewiHuqNdzBS
EgpgJRiJWv1rmdKAiM0LkAqWN242PPeAEuXXFvcGp7xDjgk5vUCvN/GwPwrMejOsBDv3ReiRG+6l
W5hVV7qk+w+GdiKTFFPJHwap6+LUsSP9CaSeSkzRjTkYzeoPAhDJX5Z10tE8T4czHKVenoTPsqEn
vtZDs/SRQw/XvXf7VzHQEp5n5wEijB5lFnEOuWRfl2+Znz/WUkA0N7fqDxswp0OYiLhRuNNT+Krf
hIxNhEoDz8k8VkbpV1P/Mb37a6mtCHBJHVA0vYDCBVzPwo8ChZBOGRL3B9YMQ1mct5qA6W3xI+5b
khvLi/iwRmSA0Y0w9pPDXcSehOLQPN6VV3SqylFkyy38XgXr5idyHxtj8na7dl8eEu9bcCATDpgB
Vq85hayqG14Vu9KM031MQk2Pq1pO8FgORjDeTaV7grgbla1TDEL6y/t8Ru4o8QXGj38phrMwfGUH
EDpLR5GHVirc1Xyaolw4XRLuE9JQDf3a6w4zUYjSKn9J39qwnuwo71Oh8HN+zbSWxpAmBPd4zO+I
Ir9brhctVsHmdlQjNIMz6XOEIhKyhzYvL8dkQart2oSw8fDjEGFHWUbpz/jRD3TXb4qRZm/0POiC
A8FCchWepNN3MZVBPLUA9OwSa98kkTvrzVCPTl4rE2OAXN2Mz9CCJD/ZdBBMUXgHlW69kFhSSgLa
sb+LqwPQMvY0eq0vWFrKNvvytO7OiL5cJsLRSDiRRskSbAC99YzYY2vbNAl9rjshGdw+LQxaSpgO
TXYKaor3+kvK2HmRnmC47KBPsCt1uAboHCW7vYGBBGc3TZtg9Iu5R8U7zv/16WM+GeaMLKUGtsTW
9RKbKRjzTS596LJwG880HL/Rvxgo3Lxwdfh40uL1Oz0El1S1H8Er0TfGGINLhIPlhye+qCpYC67e
0I2ue0t0Ye+W0FTSwU6uOVChYR/g5cB/LtvdXyFA5YhaXFMvu7Kg78gV8VWtB/z9ExjEtSXaqWiP
wjVh+YyMgsmtVI485a1CcDK81hsHe00edP4OHi+Idr1YuFrLr1ObkehrOzaFc+wJGnj8TorGPT0A
CU4AMHw5PSXvq49EISW+E1AxD2qJY+IbePAg42AZ67tXFaZ/Vi3k8N2TlvxmPnDxgp1wxlbHqmWE
ub1N8U3dllZZAYwH6DtOmPsxkMhvs82qbjvpHq/I2zXS6pFNdICUd+0ndRSNFtJPcNBTqDYsHqUu
TilkXcbCVuJMbnqcrKavDPVobq8H9O2HBU7hGkRRgfevgQ9nM1qmwyDENXicWfWroEKK/FRxJXRH
yLwqqDkBH9upWeiElIufDdTW/y/Zt//W8WAmRXTLO+crXv/cVeKMWg/4iUBYWDhiR5+ZMLbymUPP
7paUHRnzKm51xaBeTyViTZAJ3luDvtxlOaz9lenb/izendDHgLZRj8NKeyMKa6+7cH7JJ0BZdnNt
T7uQAdIS1VXpLJtKZdrJdOmcq3WsPvGKD6sl/hcEbvIz/e78Re9VZWpNAM3s4eMNKSP/7VaeGOmT
+/oQwcVxH0f5jX9L+b5lId2ITSCaP5p8Bt4HXNGgpDQK+0knPX+uhGzimx0QiUaxswD0jrWCupo9
z56cClI5i/q07JGxEXddwq5lDV9kwZthHoPm31qtgd9borJrz1RDNkrXi91MUTh0C/3FUJ17GEAl
iFht5fXSItvWYMIPaKvBkyS6eyxo2vwEEDqxzZ4QkKQ9s9KwwJUNK7H0DquXzho4vYoDqWCQ9NbM
YLqgD4BQVjamwbRPuuhDcce3lMofLNnjpTC3TiAVUilFkz0hTNOU8UHBVLctQzzqM7W09vSthMgI
hetAaBwTSvEnPLGVyYOtedTX29k6T0SOdNNVmwgWGlndDgPhFIP8fxwG71ZKqqy+OHBHu9Xrxac5
ZU9P7f7k9fyNvfc35BybUsrxiJsbQlijkZMFBvsojHjgCjJPjOs05FcUuf8eRLcW/8WyHO7vmul/
QH+B4EXIxzSyrDsD6gFlENe0lWa2ChRcYKdICEShg0XeqYB/clgwcWfyfqRv46QRK2quYGBfPlJH
oLdHtipxAHua6XYFsgDRcpen/8EHw66KzSiunUBaTqi/2yndSgF0+0zRr8lR2S4a54IRE8l4biy/
sMXhUuqmcI+RRm+VXFJNEaaMCCW2njpTIc1HmvXyAgzFQ1K4itbQ3TXEosVaFtQsC4zIFm2LQqn1
O+uv1jmG/kgEjwoQXFCZz+3ykbQy1ZzxzrZS0rPqkQQn6qH0xRRVuFKCOcQxmbVK9BDd1CZcfte1
WIw+j7wjS9tQKJ0oQ4XG8lpflIWQ26Ye1jRx5BaE3FbzoUsDZZQSe1ecgVHyH4NI5dGcUlS67t3p
qWDNdLhQI6wcpTufUrLX2DNf/PiJIooHfq+Ah+K4CycGPjmetZW+FU1eKF86a0N7l6OGgcegIIjh
ihTnPscgxWVRi8YXJKKRaB0PoG73Qs7QTCbvCx2VItmzXEAGx3zSmROM9k3FX+FBkL07J2U5xAS1
eAjrygmPfzpLKOT+TAXCpcoN9KlZltnWQN/Zofa4e2Vz9kZxCfL0dVNLezYWQqQYtrwaiX0J1rsw
8p2hM3WWeNSlLkxUhGpNxIyoCTAHxyUjTqIWUasnUVbR3k2jwKR9qqLGLyQRks7TOYuudSsLKzOw
JFOWzG6xNzo8WcwcK5W6yP/8KBByWzm4iDyvdvuxFeDBDCtLGFLtMWJXicx3MBEzKFy/owTH3mPc
FXOK72bu+/7Ti1X601UmndH7GCGmBkLC1B0iIk89+Hpxmd9BleccNpNrMsLuMbTFBvZt6XXS8eHT
r1qhGKO8E03Uwc+tHJJoWEfmrFkqRSVUGiiEqhvwh6rcL+Y31sGejFsmlwlhLpa659CEm+LqACK1
8L3B+Y1J5QhXi4fu7rMVCi7d7ziICMffIfzYm2NXtBhszHd0DJMcoh597kyjoRknl0JUA5nrLqXM
G63IDQbsbvaNt3roDS2xeu1v5MuwraIsFDOkUG8miy+60gwkvxhswsw9fd77ruByrK4PRl1Za/jd
wYDxibgGyCxntWf2nzSiDXOl48Hf+LLZbM5DZut9ymQgHAuomERKJrgh4efeLoMtixWOhfbITFfK
bOZYte6mXh4hIgCulP3UvflcGJFtYErYgecYKw42qADr8RIA7Co9HYYsMZp1cXgJRSpUUBt8rYYH
7Ls/gvJIUA7XHzFHoxTKm358zDDuFDmOmVO/a5P1Min4y30aKmICdLPzOmf3BEsD3FEPK4cyFA8I
m8GoGbIALe92ArLm/xnTsd8UJMFiZn6tPpLyiCUGu6RWXI3pkodg/6ZncYvcnKdZBfcxNCk2xovi
z6Wuk81ksltOjNs14dg4+w0a1Xrm6cLooEaO/NmZ1QcuxcMNpi+XIRv+j6eP9hejbqBoHVmG2OlI
dznv3JyVcaB5VQIVjCLGWcC8DnpH9zTbw2ZYj+BvvW22rTRoALTVWWNNTefA8Gl66z0edRjVxPGC
C5A2pybm6dFd9GIQ863Gyf1sMVncG+80ausqhDR24tKd1O5Ro5QTunRgTPD+7RP3/g6q2mibq6GW
4nbIfu+Sk26+jnMkdBTD9I5afFyrnlT4VlSZbQT15fBhgN9SMOeFzCRf7QyrisEFTJZ9ZkLfGI4c
ImuOC4XBvb733aCuyiI7QL1euiNPg7o3bchuEJIpo5fDbUqqZfiZ27bl1iEjX7VRScepEYWTTj3m
N32RuOx3N+SfnLNWxnVDW6aRpnfko3b2pNzbMqegVrFrQrybYpRcQyKIBWc7ertpnDNbdOnTj8Cn
XByxXn/Vj01uOd5AhaQmFn+0U7UrGoCmKvqaLd3Kfi5MCtov2dC3K3Qyp1j/I6bu/JjIvxrz0bOf
L7J2D6m/s3mrFfyVuk1cVCXG2Pxu+xUEhAfKOmLaJ5cbA0Z6Ph95Sak/i4JIA1Ew8xKACsXo0Tpq
LilbD7yAIsdwaI3uSxXdgA/kmp5C17zhISSAQ39L4BjosYYsH+0IlfKjwgTPHg3xRx6Y3QMZgFxe
G8WBPTc7DvwxldD8JKalWa0Jl2SEu3OdO/EkLl1eI5c5/EcaIZMG/HA02S840WbtyjmUu/N46/sC
PNgxgJHpRVxhJyj+ccJMdqs6r8fDcw9QAPf/c0VXsbpi3iVhlCsvFjR/EWF5t9q20Q+UDYB4woY4
FCpDEtM4vdsxup3iDqcZxIhR/wVzifERTLdhQHoTQoCYTLydJH7T4rcQYzQzI7aWDKfnDYjAcRnB
AF8tTlTQmAqW/f3ZCI5jsHt2W4JrrWPFvBSMh+67iDHpYW7sx2+5HQEEtAyi9hjmjUAiDT6CJ+e7
JEZCMVFLMV552hFXEQXBwlW0xadGRxrI9d6S58i2UKTM4CL8zJycvyr5Vrv6c1+fAVC9dhP72dg3
6cXjqaEcbPXj5VA6qUwf0XWgFjactECGszJfRc9vaivcBanJ0i6TGudPAvnV74o5j5s1untY+XGS
ZiXcIbd7vAIAQph3F7KtbodaB48/+JcWCMs5TquAbaE9kr/OrxfC7LsuS+TeWvb9XOVg80BMsZ5Y
N8v3TFzgm0i5VGly2Bca7flyjscXsxJDcrXsp6tjZakCUBpbb1/YqD+JQY3Q7c4fScyB67P1qZkA
f7HgWlPyaoxS1bIE76Sz/zdBkBthGzL/BaYhbU6PCRMyak24qCP0SmXbJsvwf8OTZTZAQbuXu+WR
HZc4riY82iVVHro2+439h3xVqV5d3ulNEzJMO6KyOiAMObF6fFMKP3oZH+qCSjcj1ZH0knECrUDL
HPmoVuy22RX32/Eibp7ENqLPGq44374EWxidLEJT0xnOvsDmZeMdsqjYqB5ybCAs27ijA4uPJ1q2
h3E5DMugLiVC+lEdJFYp0flUJc56+gcxE4OKRMmsZ6HjHLFfLii2kRLQ2+iEb0UQ9XpQDKwaJcgj
rEyzqt43sdqKQVLysXov9KGotAv/Yub04wMkjGvIohJxO/Ti20xKu/dLT0kMdGorwjQw/M6F7MAb
1/MOcuHzcyVrhgrJDLh3uDxWBzBIm+T0lTgssOLF9zSsHdsDozYmR44NAq8YwBKHawN4pDkm94X/
gaAj9J3dki/56OUSTXtEwcCR3Fm/RbfG9vG4+JxWVc29sKbw1Ldsj+38emO0WJHs8TtaALCPg/WX
gGMdXYwRQ6tWH7l11ZfS5L06KL0bsk7EN3iczT0eljxaxiqvg7gcVxCeR6bAM7tSBMgqXj3XqZ6H
BbMJYALnayrHiU1Vl0z7WLC3g5AiYGazZw/tPTJtK+WChF/oYTX2f0RUwirG6+WQrPVg7Iqb+uNR
4n378z0LSe/xSZJyYs1bPwPqF8cClhWngGO90XRnZGabv0Fz9bOe9EBqwr6r+Lgs19HG9OdcXzKo
HV/p3Yjthbiy4rZOfkxQZTm1dbYj3njeQ4asc18wSS0k1ZLHr8txvat1552T/W5LDLz/jsuMJ3j5
LoICPQIGQRo5tuJBlZn0xJJygZ2nwJ5CUA1evf5qUidqDjUF7iWCpt4UhVSIae/CBcXdQCeZw8P7
vS2gU4c+pn9MMh3qvZK52rIu6HJgPlJCPu9rf8MlsKe9uvNJVEkmYJzDGbYmaiwHVZ0MikFnNK52
KB2CMyu9yhvI0QsW2S7bmHJjU2HLBRXZJn+apkK0G5YFBKEZtjZBmmFzsv86iqn6J5Fjt8RSnlvz
TUcyo29LBmd75TX74B01lhKWJP/HrjBhL6na2iGoQUd2FpudK2w/oWaBRkOeXTUkcfKUg7yl0iqF
2PTn7sUKa32To2Jc0ybztjqhHMyjKPlfZh48R0qy+B/aros+8sCIIGeBaAWD3K3ffqHZ+DPKt9jT
ptkr4jonfitRB3x1xDZ3Vc+XiKrmDAeVXEeLNvJYQSR5ne/MfkoSv9HFIplE8LqFa1IQRg/kJaPI
wJkU7JMY0G/qiLtUUz2hOg5UMEM51nGVi2QSS3kXWnx8qoRHTmbMZzVhdiwt03Xi1Q2ZxP1Dx3P7
a31IFhjdm+2OppFNhbwlO0KiTJNkZ5E0mcKk+61FmoK3ryTe7XVp/FkEW2PG0Ab7bJkEVhvsUIjp
+cGb4ay8rJjYwex6/XYnBXng3Rdp6YtJQS8RzjYW7v1dAXxskjgORrwlmx0pc+lA+pphkadcgLBB
ls3jO+uc/a4RPW04wLk35RtoeyLGy3XwxTZ9A4/KDbrXlHvd2BJtoSILNq677mG0D7d6T3t+O2pS
d/oSvNaL+WCHRD5A6GdL2hR1wtWQnP+e9fggCo+oH5Ywwheigjw0AjOjeE/cvKGzTT2Aa+1fUYJr
B/ZJNTPDM8hFvq/uDUOwCofPl2bO1ZP2n3jAUfodIyEO3UXFdDyv66ODRGZamJWkH0bkzDApAhEp
D9hVmv6jVpCYUCvapArHAL4loEX2/NbnYCyzh2zUKe4dxtfqDjfdrgCkn+LD/pvjpuYJkoPc4wvJ
XOTRUjTbmRc889ZQfkja4VSpY+E7BlUUzrqHzfJGNXh+gNJxdMT55ZerN1bK06MqlFsEXPX3YCFg
0tzoKod376anuK1vXPVhzoNjni3TbpbgMKFG7GVRgy/6UTmdpPkzcNHXpwdwlPzq8gxKJwhyKp7f
wa3oYmmMidKiHJbxWBZUTYcxCa+QcMtTgoues/WcC3cmuOHLXlusLvyi72YPT3xioepn3neloZ5t
q9spYwMEjpu8Q3mWXmhe4DzXaR49FYAi9H4AjmIOwWTMW6JGNIQUqKblE5d/RRbVZy/xOpPDYxoa
RrC7PEeDMVssZ+d/JQ3t8w3lkXUYEtLOpuo/06n1aRHM281ImSl29mRfONrAUJfbiM5KANhtn+tG
zw4eIiLwsWgyfWTEQwiJ//AqavPV5jX5CLnYpzaq5U/iDq8oeWTDo1QkmVBksrqzgfpgdw8I8CD7
iM3VndliQeHBJhfIhDYpaoWmY61aObZU11j9G3XrdmhHCmRpQKLoLxYHaH5FiMv4ZTebi1qBiWWG
TkRIbO+AQLfmzljo3MdsZ9Vlq7oEbwFf+U/uA344cH20aM+FLAy783os3+2JzCBQDLemh44SCujl
rFtGdx1sIYPxu4ICkKekh/FbVqUpilF7rseJxSJr27RJtVAnMoNFfl1JPTAzVPba+9OXP+zSVWoV
3fcHS6U5aycYGbG/m9wk14q5OpMJYgdF7r6xbZesz+0fXSj0wVBAg2yg2DRkzndc4HU/EyNy21je
NvmOVZTvdoUUgncJv+lUY6svS9Ifb2kNiA13FpEjgMapTDG50rW6e/rimCDXDkbMY+5TyfwlZgWe
1BSrG0ynS8t09FqKTqr0N7CvOoK+QCO5divaZ5zyPuhD6FXdErnqSmyeHYB/6jA5LzF2p20eGz0y
qFMznN0ovzPd87/0WuXiFu6CogVS+MiPc+EM6hI2fjJswTmyvzS52YY8jmX6UKksChLOsx0FJZJt
aOkeAdnNeWEfbzg6o3nwOX0jqxayMtozoWQSbvLg2yq5aqW8MjH4cgliqqA3mBohJvaY3bEQDbUQ
Ps390VxiA5/Y5Y+PoNJsp/4BubQsqrnbrbOUTr8rvUFVqSfSK7ij6mh0Ck+VNA+rEDNc/9dv+nS5
73TQwk7jkJ275lP5im0U9VK6q2vqLpn1WHVx8x4XLNpHqMLzrGVzlm89El8XSTJeVYcIwZGMxMEo
hRJY5xgB6llYTU0joMtVUrs0tJT6DM5Te4Ls605ZdAOPaeAuB/4H3Hh++XmETG7RJ2HfyGT4xXFi
b4uMk75cFid7frOC+utn9+IKdxs5yPY3xaV5sKZw97iT5jRe5fE4/OAaQr5dMXE8FZNiaHdqCvsw
uJnj9n5My2ET7HwFunjcnjV0fP5ebSPFx/iMy8SBtiPCgyfzGEx5l8mu20FYWFxiLkDVPbQozwqr
Z8dOPyPJYEToN/BLdOOSYMeAueyXRVeVZisFw07jQmPQ/GqGhi57XdsN1ChOpX+od4JVdqYzHTJf
s0S0iUMsxeM5WEXFqU3KMp8YAt0jEzdcNs8MZacDAgjOYkkEZd3jnA+s50Pw5wcl7l60QlQrcyVE
UUl5pnqdVCK+XA+z+KQjYqEbVYzrWuiH9eUK5fGY38yX5R1YIqhtjx361HN+hd6+taijfjA4yCTZ
s/Z+Lo9KGLwwnBaK/u9PkMSNZv2voOu+/9aQ8HjDay7FPZzvTvcNDUFTES7C4V7pANTgdpLN0zSi
S3lnaISLH/KfnzuvBLJs/c6fPXNBVhON+YReekF+ZR+633sTReICww11Yj6r0ozNwdwDibaOPsCJ
568/fIrFmHT1Kye4kukgFyK7AUGbuOT7sIOlcgr7gPzmaWsIP0o+8na8mdHWFXPx/MYox4IhXfWI
We9o81HtZISDU3CxRmhWfo4Qu9FF/X/bmJ9BwI7KeajVNcXU18e2x2XC0Oj8WYNTDLspZXVik2lQ
7jp7owK6Px+IjUY6I+dtZ7W5W9lzfQ6YyHvI/t4j7Rl2BZkxyKyEGXj6eNbc68AYMulwkhp9ij1x
AXQJ2Zyx+koESVeRDJPCEugPwvwYP98TWt6i+o6xLf1/uQprstlj9787+iVWnh5PXy7tVXQO8Mx3
GJgl7zi2lIm7CLR2/VKxmcFVZ9mZJau5mH1lHJndaf8GWfHps4HxaQWRY1iVLE2ynUi2dsEXHadq
gWiKkyiKkLI4MJIbg53UjDwYLqW4WNPtitmNXOG/VLbzFjWghYqV8Iuf0xvA25uKHRLx+j/xSigr
mlgCqm1rrSc5ByDeoP36kV+t1mC0P+bnWgEEeAFo7sStvYjuuSwhKfTh+//tEjh1Mhd2SqihOvGA
jGF0HaPUdLtDxI0Z638tJaNC306lRj5XM713F+p9RC58xhMkHH2mtjmPtsbUpxSxoC7NHK8kOiKx
G4XUfNQJMR+Yt2eblX24MceB9/UwkwIr/xF1ubkYYDQUkVk1sxiHopKjlQ3sAKsHYzxLLfx7SsH4
HcGUS8Gqh3boRxAGWlM5TlmpIF0xe65gGRWdg4PqisW5WaU/yZWJV03JebariPqhpDX+mTOTSfPh
tOH6s358adZMhp7wkalLUztvTpqRB/L7TwclNFOhMVH5eV0ePk/ZFFFSp8sqL+OieQv+VHJZnGuj
uSweEm/xq42gbwF8tRIsmuRDbY13rEV1+hqoOavnEh0FRzzV+8oLcfL2LhPD7/AApN4pSgiIVV+U
b1gYel5xfDl8zLwkSK/NDYa+Y8ZdZ26BNP6o3WzEVYlDrhmdTQS7PPLYOiYk6w1guziKVmZiZUKX
YsnFBGiugiGXDUDEkMLXtd4LYzuy4PsNxazKZvShKqKF2Ay604vXsStBttHh30WXV1rLvUK29AkZ
hPEfEfl0n9vX6fyxFt7qIQ8P2uDQucjBvOMHaVRimFDcqTQFiIzokw/62sKdLd9rh6uFXOQucuQl
IvDukStNB4OHE/zBHiboT5wLZKRLoFZGNaIQMb48ZfXYT0SdaMelD8XH8EYHz5Qhq4G3NNIQj4D0
9VdrgC2j7SPGs1zr8cjnuhDeYpcPaCq+SbR8B0/C7ChA2l7dJcI9cv+XM0WYZNXeftQuFM0rkd5S
pHUsktgGEKb4J2fSSflAaoeeKvJkiHfGcBFosHUs6m9f1oIvyLTfMj+JXWoV129sO0yWLTBY4F0b
gzR7RWByTUfnKUsMErZPS+vta26o/2C0Ww6SK0Ob2eg/wqAXt46iafoEM775WJBmzO6iMGz54276
/gfBlx0+WT74nrzunkkGy7qAGlw8ErCDCVTBpoMCNej36kYX239ed51DKyMgas+gnw1KSRn5ZS3P
jcycN/eN0GIKIkhVz+cp9NkpwX2N/jpta8BGvLRYhejw+oprIxirB2Mj5DCI0b/3gl0EsY371jEt
6hQMb6nrOGhsQL/C2QBcKZnGvtJomuIC1fKYZJBlVExt6zhgPeDOZruyFY1+nYJhjR7192vK0X64
9Z8H5alp06AYAXi9UPr1Sg9fM87WIeanWgomfc/hTq3+lw22x1L12RiRkztNYML/J9fh2uuAVoQe
GDjFxsIt6cOjizszzAcNBONFIZz0y3xZBkA8VquGzDM0LMMsRc30cuyCNswxX7hUzGmreFSvzZTz
f0pH/dy0hvH+s4gorfg7JQjoggnzNWplOfVQkbaDxUyIudMo/NWolsEhQj4PvPPtxuy3HuKxmpi3
YQ8ztK7TLG8tqcZMf2QQQW4B9qHOTNlijHv/V8uP3D+FJg7Ig2jPQG0Z5azd5n0jiWqC+QNj8EqN
8qYztmiz/lY4Y6Pd+b9bt8VuumrG3Ic3Sn3kA8easi/QNsH62kB8/SYor2qXN+pey+lMDVb+Uesm
WhFwGjTjZQny5RQRp64XIVdDE7jPorA0yWTaf3icWb+lw4S64mMday8Nda+kW5ViaEAyK9xjZ49C
BWr0DonVpym6jHtDm/9qpYMMNUA4KZv6Ee796jdtOTCjb1LH/QJXXlDnnGxl5vHG4WR1Knaa9AeM
csPIkTAuBEA700rVdquwK7BLRdBLHgqC6qPs23RxFJiLgIFMT9aGnr7xd0lDo0Ug96t5cr8t7G9f
oo9bVW4L4y7tpcv3svtIkVWDBBCbH8rohkxRbKpp0Y9sLOEN+4YhX9qTKSGuW1EixX8Lo6ER0dcH
LopGZ+hLwlWdj/F/oZCo6XaEYeK4ZSiXbRFvvCkBxZlaqR8+waGbP6ttEpNutVXrLgCyKr8Pp1Mm
EKhoVjbEUpT0UBwoCbsqSa6WUKL/3GtAH9MLS6aaVquZo4pFEC3Xg+u3oikY+i8pS8dIIBbcx6mN
Z9YyD6Ky6dgEeEQMkjyyNNEe1HvVCBzkTb9LEhww+R86mibahG4KgguP/Lowbki2bdaKg2nraw1F
ufhu5DB5HCG6OQhQMdb3I/RNjN+uGxd5A6GQ4A7EPQE/+jl/XMAlJFMFKY2wvCZNuPlh7PD7R8dG
QH8kOkyAeG8fdnRekxdtOQhs1fFuXkU4XjASp4ZkPnDXltCZweSFqaor8lpqTUqBx+KuBcAQiglv
DLBcDWlXjJCsKQjApTAk8oousdCloUWdjNikkDcXSUkl6PrbfPIevfkxhe1m1s1TztZYcsnrTib2
3aQQLSty/8yYJ1ab34tRCbCM0fRli8W+j5IKsy3c5ysSDvfuX9XSWopmZMxsG3VfKK2HBwwul47G
zFkPSTIxsttMdzHl82kGfqL/K3E67BMvqzpzgad4c8h+u5vmUUc3ni4K3mOmWYWNwx2L9yhAXEYK
EBSZGXiXf/NOT+pgkkcDqBqNdhXOh/myFIdp3u2fvzrn8G7StrxAAcmGZ78xNvnvZMiQ2m7isdg1
2/Czdx9wEUmG3z1OCkrCK+BI56A4dJHOi35wkBxhFpNPW8BF2cpTLmubKyhn6xWz1F8RE2mzoea0
jBKC8llGi9RtkQ/sHxFUGBPF3uR7Nm+vcYUBUEAenNCBm/ivuksclEXRY8pV6xQLFHGOwUwH7JKF
eA7ccVaFBzH4Dz90Njzcwk3JPc0yqOuSPvHr7XAtOHFEM9nM+jlBnodU7eZGdQgsDKL+ItTqJnZn
FtNBm1xXT7nJZ+fwLggeHqoYVxZZbnP8zFkdQBlz5y4vozrzVzi3WN14kVzs0/nSrpjBoTkULmI/
U8q+9q9oTRShjqn3Mk1+fyIM9pWhcdLXrXPK3pHg083dPjbRKIrkEtCVuaddkgWpVLCQ8oQQUgUd
JjF/YthpR9HBREX0Pvo94iNY4vd2E2t58B/1UO3bCLtPXVxD4HFm84nAbT7OnqsJs5Tn3MKd/vOa
o9Pc3LzPvwslx5KrR5z9RPQJKIBWOWXBQTErdSlfgEwM4epr3mo9KsgTBJLfWi1pZJXEKT+RzHxd
MMU+J+b0/oznkE5m1FGK6NVYH1SHAEsZOkLUl3vzJNDBXJS48MRQijUPBLkA1QVjWXzt1Irs7SP/
f8C74hUkcp0fJL5/PWCvyyJ4pzBF04O6hsDkvtwa3S5mJPwgnhCM/BurGz7pl9tuCWHwzv1yyQuM
dYtVdNXOFmg5EJQgV9+WLrXbJaZL6bqcHUqHaePfc+0OsHoeY2jeuhrNGY9GonY5TykTpJL80EwU
lJeS376/AdQz+TWIKxBp4rUU+f4IFJ6OEKBEiT6QOocN3FsSRyRf1XAGdt/UzFjsNZWZUwSEVEEc
RurH3sq2PSh+ezGzncHLl/ZhZKG3Ql5oYyss12vxYLjuQuWN0alP63oEOjR91LlKcDbgq/9Q3gIf
wyEUD8XTSeFHRSbTmXtEv9rcKFdahTagTaAB2WQYQ2M4lMxxEj4vnxrzGGKHE+tRNWrih0tZncMl
mOeYhyVHA+tEY2mrrMm5FvgCZF0pnDtzD6y67dorL1UiJCWWJulwJbrAFmQOk7QtMWiiDMj93XJ+
KF5nyq8t1XREKjdd8ZuHEPAEhEuU5R4Wxxf74ozbAoWux9pRiRn8kNSzCmKNDlYT2I7iInSoDpwR
KUKAxrlt2azIeaYAUacWS9bQdjK9oWb9/RlpOPpu+NomYHM8gbvk1fWu3SNOvIuwmoawv5Pz5ZC1
S1JYE/yh8rM8nMdiIUo4k1gkX/fZbWVlIwTCSqmtDgYOUVhWEbwfbIPfxHZ1Qs7faVusJZTjIMm1
GRN6ZETiIZJ+uH7rUoOJwAl3jJnin6J/FToRms6YrPt8QlSO0u0PMAci3bCP27Itectyro2ov1iB
7kPtTCn1S1xDaFjqaSVAK1fx8SRe7M3a3hLUVFfHkVFwu+W2Alq9SRze9zOJwafL4qjh7mjWW/5j
/71zqIrJqT1cmZnM2G8a0TRyTrv16Z7tI1xrBK8QercLEezcWZXIki9e4rsnmonsVz9+FF5ALzfU
yB+bKWbbSvK//z8LWXDwJNGyyoLdKB7ldr12fGoN2QJYNeWnGYwuUKhEU27c41ICCbJilvC9r4jd
6iX4DUerCgZHqy1nBJbofNpacIgiXd18mQJJBrWygEfav6JtBxYGhiPtfKgZ92KGb4hBFYNtbl8J
YxijakkfrC8/pjMdidUZfH9clTOflP19qQsnaO5CkzYzVM7ex0FHh1mHeMyc8L8OJcBThY8LTIvY
Lr/3ImbWcRJh8oS873SiJpHkolIaxvdbaxN/vUUL1zjG8+HaYDeCIaM8vk0Xcdt6jdYe5x+fX4iN
O1wWprxtGRXB2BB0LyuI9BW5UX6OeZiPcpPGwkPDElPhmt9ZfNNhT2F75FGCZynQdgKsRSNeIKqV
qlV8qdTEe12aEyrdX4c64TIIz6cDFno2+/wRtAyJ3gL8eTH9CfIbs6XMrIshZbgSw6lS04PThkNT
7DFr6Du2TmwcnHcrLtuc/eOZnGZSDZocAF7xsFcx2gatyreuLD2qunV0O/PCfH1mVDjHLbdD9Ix5
KAM27vtCzPwatS9Rl6a/CpOW3TdulFJYl1/AaP5S5UX+6Pj8zQ2nr+uBjExRIR8jnKnfJQkOwrkw
KgT/ODSwA1SXAy9iLZDULEJMZ7CECgvfOShJa5mGeefpLDKHvlz2Q6qWnkR1agoaMWYiOBHxtY0+
8p55A7WO0ERyLFqW6MGI7K2b1kOQ8gUPjXKc+1zf6sWCaTY3wTI27QxAmsLdq9wDH2bCnry2Mftw
YZXqiA3Alg2exhCZ5wXLUFXvRxrDRtEhix4qCUAKO3feUD5tg7y0/IKlJzvPKerAlyJbPze3rzOn
0xu3F3b2qOJRXidzlAGWhGvl19h5+74pC8AvK3Vh8Oi96/mq9CUmQmUzjup7ZP0oLaUoXsKM4BtE
GJD+ALjHIA3mREqL60p9ObvJV0eIRgMOeW4e4FBKEOkyMK7Wuftjf8DshGZR1zv5cz4DPOAEsdtl
AR2XswaoJ/zFfiBGJMtsL+aKwFbRAcJ6XSLpS4K9qv+dJtE7HdtSzrO1k0jV1JlRr/kCMWUrsdJq
a1aMe88dJDvLigGqIwCmdAGI7VN7rFbNcjErSqWNHj4zPt3tboYeiOSZHg+p07zI+eQEB+DRO5Gg
zpe5JjagWFwp2h2+iuAcTUKwRMeEvUPBp4aOfk63gTe/Byd8V+wipFqBZtqJ++lTAKdAy1jJ/g9Q
Zkg+vyKhWjMW78mtAC8e/zPP3GgbaZ7ID/V1vxUjHDXM13iT2QFExjReK9y4OEHk4oU29D0MDXjo
e0Gx5kaybRT0yKbw4dO0CHDPvo+VTxECht7p6qq/Uuk1dg425LWTQ0RFx1uXK9lWpMdF9MxynvDP
CKonxWAJeqBVsE/LvMQaYZfH9j8se2iZCtNIRPFMZtY12pWmnpG5AVbbpjgybkzpwdLdwNqQAXtZ
NkFeHKECBfz8GMJoSudZNG+8KGpORXcqXtAQbOD50CGP8ZMkTwNz0aKVMCr+rqirvO0GPpsJmQhw
kU4mnkto1P35zHodQwthMCabSjOr9KN/T8klKEefZ2ZsGCQa1mP5U81X3FYOS1RZ7xzJzw6wZ5qu
BfpA1bGt/gY5extctT/WJMh/4m7kLJbeu6opqwwg2JsrYa/H6tyI+tC9BP41OmKZrQSTdKHMB5P6
0/ojBUr20QvwJX/1BvnGPE7b0fM3a88FZCsSNQnt1yfOUjnUJ/Di5BJDdLdKLI38LeFI4j0MHKdW
TM8/EXV2r2MITJcRut31/xuSI5trAgZlHuDctk7hP/mz1LVIO0uqmbXfOdOBIKh67QFClLuHjVD8
00zVfc6Gj5A1xYq8k4IciagXC3WglEJtMRjPcLpCP80RbEK/Id0baZ10pC5shNVqFDOQjNpNSGnz
GAIXKqt/J1zleR9veLp7/gwGgyJ6+bgalyJ7YB8zDPsJBlZNw6fJGlXNP19bGWgdlQCD2BOnPxkr
uKggWrMYjEuWTODKCLJYtizGTIkMO6XM7XGCv9cwqKvxNNsf2JZzOue6P8c7KSLJkaz1EwIVcbiW
hoSFerMB9ILFAU18w8jUVMS2uH/H9DOIbp0jarU23Zbsdrhec5N1hTf/LnEeWmDJkVMp+r6ytCjl
BvJ3BoDUBeGiAHuTWs8NtDTJJ3bSzZpXxbxzglBR7xWKXBqM7suZxRYd2Jx+H1XIdMy3v3TJwIQq
T1knwUPk9Sws12bt80JGAy5d15EPo8Bw9rPPFM+odIJvz5CQz1LUJo5njoMsdEFAHnN0173zhQaN
OOSkAya4lKZWyfWVcLZcBTQrZ6wk9k9CMMU2KNq+NWY7iWclOrPGAg3axxCCc4Rn3AOZkgZR/Z5+
rjVT9P6bg/SQIHbG2tMnyDQQxaUmz3coQZAOruGctqSosiSZQi2S5JtJAxqrM6WJjprrulV82EJJ
TswdlWmE3vd/M3ID8nuNAZ0ca1hSV2cwW19FZbjmu5+hxdsyQJWsleUY6hC7xQIJWxfj10mDYoYt
RAUWofxYaKZgq0TpniZvLokq2En/4Tn2QOuVtsrOGDZYyX7G5yZ9KLijebSUEbIE9OUlCmBm4vWy
6usCjIxVaKrK/c5Wry+kU3NRq4k9n2Mvqku2kYkgVNw5Jb8i1UY2ouUu1kd/RAjAfSPDgBYrRr76
/6/IjP/IXIMWrsView3TQUOxBdw15Qg17rwCf+a/92MC3Xl7y0Lib/PVKxzOH/mB0oV/8chk0PF6
lra/E5rgtwuTshVGN84LjZARK5aCRicVF1sGLCBDMTxOmvnUaYz2QQRbvNPtslxhqFARqQRJniIK
b1L/nWlzy2HdtBh6XSJkmyuiF5kqb9TY3iGnlIOL4HmpOgsKBx/N4/ijdPUuJ0VVtpFB8CMmlwOH
+hc43b+ROangoP+zQby26Hs0FIGYj/TkXM9xd6jZIK8hLn5KD9gZ2cZAfnocTcMXbfLdX3QleAYd
vIdXjvomkrsOmubECjvQ81ISOwyzI8Hn741tWAmEaafzNaYE6ss5n9uzqJfe0H2UC4HOQ2fGNSvQ
RhAxjCuvSCNpaxh/2WUS6JJ/mfVHRuppzjUnZSAkCFyhUcUPcmp+cQrz6iG0Q7yhXRXWhWgm+JvJ
Uo023V48Y45BzAZcr5rnSr9NaFVBD9UKhSrOpRpa3F5gzMFOhMVNTxHLZ0FiSCQ6MRSiBvlWrVH1
GWvLQm9/904a/N1y2Ri7QoSYiUcqrp7TWc1Jx5vqXKJCOSiqRuNSXs6x/30wzTP7ZRnUIMZVbD5n
W0YIjQbySzHUHJ+7R7Ik8YiXnSKyBVzFQvKXbL/6ozLmhbsHJh9p4eo0KW0FlKVeBC6on6f4IZuk
iDO87FK/9xte/c3ELqWzm6GrbEuUzvqQ0xYnChhmuC2ZGsys91p4cF5GMElrJTS4P6yUn6C8PnC9
bXslwSPI5yvsP/r2nCPq3Z+dhIiRZdLw35JM7R4hnmgam4PeSs2kkucFCqlcuJJNhsxmTKJthI7V
jxzferFBGSuJ4S0CbWFceuMX+weflwZrk3WVgHQZAFqKB0qD9cMY9TtdQrPasRdZ/EF1FENuLsod
aomWXUMarkA4aKX6MMVIOzCapsgrs2yQEPhU/L5oMVqAnZjKbVEsxFYbUAvOvAPvJ8i/nLt57Jni
RSWuhxh3pkLhFwbpmJv1g8R5KHJa3A6S8r3h2syXSGOOPHKS5HvsbZl0DDtBsbWy2BxV3KSLjsbv
80f/yXIpx5Y4sxjYguRiv/rK3AH9kQOel5HtN87V4Ghj8GvnzJftHH2tbevYy5UyfrDfEy7jnZL3
gymDVy09EPCosq4/P2zeuz0BI+5i/DqWqRM6gwI/0dvKw/t2Rnjqq6k6w4aNHmfTkjzlWH1hrKg7
gFLq9UdEuJPG70k2I/MwQuP89YZkdUBX1uLYVL+OesAGdX1KU4QLmZAcaJ3bE1bEzkPNF/xfNKRH
leRcV7Nt2udq8XibOtWoKZbKYEemTPe8rhY9T6TuKBzYyYGcibEVI21ttTdLSkPQ2CR5ORk8Pbd+
jrfQ93CAbWQYH1NadIllKuqKlk9o8fy419pDvPHazO2mABoEmF2KHmOJsZTIVRA3IJWG6/+UB6YC
jgiziVRAtbyS9JhrfiaI7L/jEodn8BTACnR/QjWoMNrBnmUINJBozpFcOGYTV28A17w8hwb+2/Rf
xxZtMIU91RnwPC1mD67kumcs5Bno5Yrj9cCEDzytSkod33hbm5Vl6lRmD/93KMMmnmIMTziQRNIK
iUgrn0z1/c5wPJEGI/CMw88DgJ70j+HRp4yDGCEeyXL89TmY3QL8O512iTjYsNbFLnDFUMmrCGWS
LAoylG3qMMoTf5CKR48bzxeh6tiLlEsiTHM2bDL2/m6EtHk+RQDxK2CSDBEYhnPRyDrjQdQPY5BW
An58Ah+DktvbBvi146koZKEBOxYWWePWB3s/CDRnb883QdJbDfsd2nhW02gKpl44Oth+q4gyd+w3
LOR3GxpIFhlc7BfVPqbnlKxLFEP+kLBL57HbHYxdDeZr4EBQqpYAqXZV8X661/dIUlyTKR1Iur0b
aQ2Fk/vfpaPpcWcqn8zrFm3kVy2tJAOGowK3MJNtmigDGbfe42HiEMWNn9ahJBl0o6Lff3xYtjvx
6v+BMfgTKRPd+pJn2Tl61ze+ZdOihtIU018i97B37hwvLaGoDVGGGCFyEg/Idlz7NrJRBl+HUK89
8twLQCQZKB6349kulhYyWG6aXSI+GEwJHqnieT7AF1KMJtjl84GeIs/wTLkLuuI2g6PQ+16/3F/u
Qs0x4tkFQHUreGiemsEu8yFljH+Nqa7NWmxXKhA4HuVbW8/yT2U1/wdcSSRze32e4cxek/pBOAtf
Lm0RiFq9bfmLPcpqO5q79kd3JelQqR+23oV4Nj0zgtOqgFzW/UooygCj1Mfdn1fGbDA9sxer/jOY
T8T8mH/YNViI0RlZQSopGDv717v+U2x8Es83OLrRTutsSgASHVUcpAG4dHJInNMmEgQtQhOr8ZRU
7DpfAAUFz4BaDmk95QzA2oDvuGzuIUcvX3fHOpXgmpLeZdok0sFTrU9VuZXHXBrFFxlBnxryS4Jh
o9ljyg8NYj8fAw+h6NppTZW/+xHkpdxvsZhE1MQ/VN44fHk/Qagt/OdebDIFfF8pLRVixnMMyYa9
A658CgWJpBtxaCNaUGKjbsQOn4bMrExj0bJNSPG6eLd3k/xMjdncERkVGg/IXo6k/Ud6D8rEHN15
w3tP1fbXEB7pUNXOOrgohgaueiEEkVrjAAZnsMW68a2tAvjVo7qlmWY75vn+JgZbdyMktQZcWwPS
hsy5B9BNjjb3mBewO6RPs26N7+4W++R7FDjZUpiTmlOi74u5vhBIReJfvPTR5q7Doh9zDVXWWLDU
A2uxSXkHX2NiYoaErIIzXURf6WbHf11zBCNbc2PEnp6S8/gm5szvvRKt8BobTQWEEutBTVBD/WEn
2JcGl3eVz6DfZlaQ1KI43ALs3QNpyiTDhiqiljhH94S9AKtAVI3QkJTHzECvJi2fvxG8r1L1Ghr0
ppy+cChlhwZqph6q/Q7AL41zEzuFnLX+p53sgrrBNl4WDcoSVBjgalNG68O1lURTFuj5bXZ87vdx
LsQ1g+ap+frbnCeFxM4bz4EieAvJ4eOAd1umZd5ZmKYqwEuwYuLnmjVcXcMemQzZRZ0420CD2tCq
ZgHynlgOwcU6DbUofqvWlM1J7rfALJvMbU1mXDsB1d/qIgqMyPHxXx0e3LWey8XWJyDZb7DwnAOX
1zedCtddibCNuYvWRx8OFfTTxElr0c0oW+/SPkqGGOgrIGoJvytzlZt4Sh/YkUELS3U6UM7ZZ8YS
s0o4J09XdXEbkORf4xWXdxtQykGjunHsMXAghkpNT+1hzhAcLfetjAE5/L5/2bZ8iI8WeU5L62xQ
t4mlAiu3UT9vDot7rZETvoW/O+Z+JgVKCEz31V2vCwRPPnejHQvy+8mvD+9c6dw+kLQL6jdqia7j
8lu3jBnghS8XD1JfTfzaG9QbQPX6gzimsOUUIpXzBmet3U50mGMkXyT1h3Hjc9MFxf5mbVMCKC3G
boNP3cXqlP8T2aJ5aemQIboPp6rn5lMhjfcwzVso1HXZwZcn7HqiqknC11YeaKE9BgjWXvGmSCrL
IJwaqjbNWBVGxGoQqRlEVEMF/VDN7Vlc2bnuFjvUbIiRln7Q/GzS73/SJ6P+62BhVx3PjTxqkiHc
/jK/TWr8jIinG5syiNbVg5uXhObY/nw29vGiSMPV9/Vg81+ncbrmpoQy37NkuJospAL7R3RMaFoy
zKqwujq+gU7jw4AIsirnydrQd1+TVmUjtywj309ihImbEDf8kRmA70imtpUxS39cEdPIQx9co5rD
lK7VPqsofLg5NtU+xAXFN4UsPRYKbaFdOZ5yyCC8dACpLnejtSz81DPxzZ7RRJpRlXINzbVQk+La
A6Cu/KVYaplNDjmlXLUHF9FBnLqyqVGzQYjQFelJWwRi5NcIObDOFKCt0x+6N8rw7tFhMLOTvS28
ZnPV+kOUML73hADFjLWRYGexR/g4MLpwMRs/z/YDcshkTUx0gpYpl92Aow3n4odox+BpbhdutgD7
mSiYGr5/9jByqgns8G7GZgKg2b32svZCT/gF0X+QZxg59etOW1fPQjU0p2n/LEtXjYx/ik83A9Y7
mj6AckddQiCO5l7jRjvWIqnMxlLhWzmCC3AJaFCoF4rPJoT1MSIDhjGVOSvfuQ4ox7GVJQ9hX768
aTvliPW+sNirPwEQ6O+A52kwCu5/baHKN3Ke43wIvZ+ZYz7eldhfow2vGJVix1EjodLdniSwoFh4
YIP52gHb0s0i34bOFr+asfuXO253thu11AOGMcIIG0gRQ/7FkFjrnw24AYCuAiAJySmOClOfWOBE
9B9epRMQ0FSoE7WLz6H5CTSWdEymjCm3Jt4czxNn1rpBs1slIXHEr1zo/SYpc1dHau8hmm11zMXj
oEqRocDt5W9UWAC3G9zI6fsIGPgvFFQIDOy7C3jZuSSln7ihphHw7gPAFVd8NTRuCeWaMuKC+x4i
jpHOHgvTb9tjfPYPIaI+T6snK1hnaJL6Zj+h4kOSBWpk87ZECKjbnAG/oyLrCq3Nmhw1ScjaRdnP
Ptvz/V15nkwS6SeX4GSVpmvfUUbaf4lMoATBTMjpmAtSAhckpbkIKAqx5EIa8UKjcQz975zXpAkF
JKzmcIpwVXIc3TOU2qPoBCHEnD2wSBvU38sPY8cq/iS+H9lJZXLL7PzLs0xthDFimDlhmWkiZG5V
svPJcQExNPe5wHZr1dWbWV/lPviL/3h0X9ZD5rDaRf/M2gLXfym8QawCJz6cGyt2PAMVAeXh90+l
EyCkHgGdi+jF+FNZRBjbLh92LwVcuhkGTd9IWd4jWc2SDDgLesyOOb9CytMvcUIYafqm2GJ2X2Rp
T5B87uKorX1wBO4awNUDjBZYgrp8RKZQNLcKS0zbFcLakQBUV1To0NwVGIaXMfvSdLLUa58LFFRy
5jLyqPZgce27xwKc19YbDJ7utO80eUzUjZ5BRBRFEYpAPpoMGftO9dehwmTlJ95357fY1LLEF/S8
H0HsL2Ic2YD2QCQavmXk8hbFG5KdPH6AeDTcWXgXmQKzFT8E9m+TC9Nl6zf9uji2JlUpu0FFc707
dJajwVZa/RneEDtnR2xRzw7z+0h54V6vQiJpnoGvgvoGN9qxhwXIWl0V/iMxqRWvRhj7KysXix6s
Qxl/2z8bJjZ1ZEb1CIRNw5btEseGXJlPpw+mEckMR5zFgPDQixKy/rLpb36/8wFagxwty0ZOWvQT
lpm1+AGJsQip1HzfpkaDktH+UoYdb14J6iKha+SSVuQ5r5TOe/YVYyOdBFXHEdIfiySb9F8z9/Ie
prS2F8038RZJUiSteaVb3w+1hWzySE9UuugiLGdB3Tib1hkqSh0z75kf45rTPiBchVgVW1K7+qrZ
ol9rXHY4PSbGaOEO036N43NKp17LHUyvnzpyXxlgXl2l29Vl0cAxgf3jQXk+4LSQUa90+xXSOuE0
M5dLgJB+oxM6fk4RI1zftjo7Ehxux8+wx+vRnZ7Te8pNbVnB0qMSohjwxWESJxqQDOboHmxEHN88
nDBtC+aCe9/hLYoKYlFi3cQdf7mkNn/ExjVqkV5wSF+Oq6DwsKShE+xxfMrEz7bXPOsh3yL3gLFR
BAcqWQxKfYZPJJLhmgEXfthAVnWqD0jZ5lylUhqHwgBShKj46Yxjt5qR+XqJsiIZSWzM/HPgLLq0
vwMfxUS7cfPnzPGulu3c1GR4iTKLNgZ8mvSQgjI6GQZFGGLIX+pxerCB4ikg09JUyKqKgJqJbL05
yb7nWr6qjgA2dKgycTqnJThrodw6V/xgxPK5jmrjBddATNcJO8U57I1Oaxw39zZ7iBxB9hEpu9ce
5w3/iwZzuWB6/xaHco1JZ6MD0nKpXiGKeuoI0Rul/vY77DAVczcF9sioD6BEj8K0c1hK+yXTFlUH
X0V7zLp6osC+A5XmiBCi3zOuhMnCjrMjmUOc3kMPL5OYPJKDxClAGRmXHMtcPiL1Um+qPjlYMuRp
LJxESHVf38nAW1l61ZpqXNw4TuwlaUy6N3PDgoultgHmek3F0ZkKx/7hzXrbP7SQVcm5iMEmLnpu
RvVxwTSMUF1qLStQTeaoIDMLT7PyRtfPrDHHETP7p1RS5u/uyvaTIVBmYo3c8NUMGy3eO2Iqy2hy
ASqBOOHRNg2449SZMXLBUaL43GAqy9WyytZLgj9i6IcNM4d1hEaxoUaZe6kt7hfNYgVVOW5BPVQJ
cLwDdNKcDfSfsD+BaBuhBGqB6SUjsSkK5ZkKh03NmB17B/MM5crgAv8xTYwVD+KE7IPlU3JMTBnQ
nuliSajm3GmSnluZm9dZOw7k4srtvzx0deofGbXopOMD6ABQbEu2tRyg1jHjhXVED1b2iIPhYoCM
VUSaYwcVXZcWXMfv24u1d3dlkZGnuMPh/frZQJTErQOthgj9g+WgNLhKy8f3NXIfOlQRzGscYQEw
GrqKi4ZTPx4JzLxVl+e9aj3usL2M+N42gcihskw0Z0UiPLMzjVoEn1BpKO+UWYPF57flP9z3DWBU
5ssm1McvY1DTKS8tBs4iyEtFdo7Uj2U98ZjP5ltJmoW+onyMYbDWF6Zbsri742VA6jVQ4w/JPSbc
R1PiRJfyBGeW6JH0jhtMK3tYP0GSdP/lX7LpZu+nge9MUkkbGfshakmQz9o1vNJRCvL6soLUMFuC
lr7lKe+ru2G35p3XoMCBBi3Smbu+edF35uOxcm+6ct0lnhGKNiw9Ui7ySMFnN9TSKWYdRPsbCk3g
fRlLC/HGOsWr0O9oUUZME5Im+mkvO8yz6H41lJcUrh9Og8xPkcARx36bNsMe7xmEmzOr7njJaF9e
DveTNg/MdHYdUl3XeyF9+rVdPTSqT9K6hYtOhzi6iOitVYf86Wlcs5VBmOLfHCFP0WK267Aw+IA+
lbU+U4AomffH06nWaMGT37HGiSe0eH1EfLPzN/3NZkDMKY4ZWMYDrsQw/Is2TLcQ6KlavAvodasD
G80QDL9IPFgxcA4Vm08bUtLoy19QN7mssYRGgX9WvESxszDSukUR8DweFJrMxysDw0z4v/yeyyHQ
+fCBkyyhU4AUP7HBVl1ec6ghfS6TicXpb5mhtavt9CzEj0OfRHrPW8WY6gLpryGkL35zPGxBQrgR
uXxZfdFqA4Q8Rx0nI51HkO6gi/5h0p1exjQDX0wux6qfClYjClRYB4SKI9PRhZ1eBSxQAQyTHQ2h
3klGkMMdKuk4I9DtX7bu7SVW7+urt7vkSvXG9NdOBZ6A2W78bsJ6S/Bv6nMr1FUpbTcH5prMwcnO
vswk87sZCaD6+lTxauu30B0ntG+OKX+dryY5dbjE82HyCoi4gR0x8nIZ91NllF33zu1Tfq20Y9d/
DD07tT+qb20kVHoBSJ24/vZhsBmQmqBcBYl+oQP6AsC2wjO4ZX3XKMGuIza4bybqKWPueDHphEJF
bWJ1m1SQTlCd5mfQk/JDKb9LYJ6xmjOUuCOVsP1p7yROXrmoRJqgMDdWlIJHxHyHnmWEQkjY5J4F
0ENmyn6fHQCTZ6WpaFIFkVqnYm5lrXtAls8jR4V9Wxm+CosdTvfylJny6ys82VuEJeqaQPyRpWsq
yTTztyjdT3IzQ8BGnZWNlOGDnPPfOWksTsXR+R6BBRu06okw6s9aqGF8FA8IH99wpO8tTiZirAfM
Uj7AT8FocP8pzHtE5ljVJUyWlsN0QRE78VdveY4bvVuy/SuJ191vBmjd6hBG6QU9I/tM45iOXw+j
d8/UjtDQbQwkWP4EhN2qDPDN42AkInjQmoQv9VfNypxYUCAmV59oYr60CYeSGWvCohtyQaBpDzNw
+eAISQnXpDat9ESklx1UdqVdRLFuOOOgQwbf2Cj+Sc9zXhvcjmmu43gV4s0QYkTMPcrUeyuNxPKX
S29C14v0oUtz5DT5jiXMKINOfMfYs8z3KmXnRHs97V19odHpVKL/JCNbtr+dHtsX4xCYudooMLSr
xJMETOnjp+teGup9/THKFx1ZU3MH6dLY3i9q0/4061JxRdTeY/qDMvSZKlWRRvIb+AKTiGfSjru2
DB8mVR3J/ZrU+qwOBpFYVg71DAlEEwQSt1jmEi8EsTET8q3l9BANaF1PwSfbCMbvXWNty6GAG33J
UW/3tciMNPZ744B9D0EVpLgdPdGzfcAQhYmNqG+98AdlFiqTlGYjguSwKez9lLiLA415xCMe1Ty7
gXR0gZq/F9VfEDoqkzyNUu6puO37+xT6yNnSuNaEVpBIhZnSpgFlFUHPNSGWxoUJ44HAGVpV+1Ey
BtNicBm3+JFzQUkiZwhMVxtFevV39xTwjLThprbF9l8/4SoegHWdSJedWJskWDcn9Qt0jO+lITSE
2c9n8ntrYuXj69EZkkem9gRMW0cARzaSsWLiU2lI4BInaDpfCyKrT35cyiqH73gEOxHVNaEA6lLx
78kbh1Mz4jHoM/UDvFu1dnrtWltqjB0lwzRitqxwfNL4V3QydSFvBa8RWar3Zp/uWXKwcre1KCdf
dFecpWjixIc3fRBwjub2klDqAiUu9UjZPUsYgcf8Ocs9DDT3mS83IDxVMv293S+wadjR8B/Wiyxf
tR93uXe8BCv/4PUBQnTyPiJuwLbndGejNbWCjo6fvTAc7iJnqyXaybbJmbxaPEASTOkTB4+H5GZw
FCijl35N8bjHPu6QJtEPvoNn58N5hARorrbQRgmr5lgqmqgxFUj/P1oBA6ptTctPBQRZKXYI5iJk
IS74YBA/El4u2b+3HYS7L/GrH7QP5JWVRyDhEWNeT628dwGmenevmh+SAPPr3S9iN1fHHkGmeaUh
b9CfDsf9Wh0BWd8O3RQfnsRqe2rG6PlENZ+gSNi64R/9j99imhPSI21wRIxZHHSc4JFXy0iK0kaB
GKJiOgrK3F/o7flQDTcQQswl/4kMri0TdKAqtaVhP6vbDQC3pTbpLZrIgg5cv0V31WIQVje3xNpA
6irQUK+2fQngRnUVCToxPgr+6AiM2q3WfofvK0f0t+ROaqWcrnd1E0Hrji8Z2ITpRzVwqHY0TOQX
r1AVT/DBwdI0A7X9ga5mvDefHdMiELIxNmq/lXramDIxEu+ABZ/H+8NaHhnxFcye2KbKv+86eGN4
dOBc6mDA0ddRzEu5EcpNRWnsMgPMXm/1DN6Y/ee1vbSULA4vpHfPnnF9nxvyR3u/UDrSy9Jt3GsH
cdTkwi3JrCbm1W9dCDyjKs1YCG0PaqQrtKiUJH7P//ph+x2mJMzXPejFJy8uclxrUgfCUfLwLeaV
A5ZEyuFCZeLY+a/Dash3guI4bpX1AuETCh5lakRR+EivgacHCPhCL4pejGhnXLaXq6i09uoxrQSe
Jqvud1J0WDZa3yyh7UXEnQCA31mr9rs/mHtvouuHXASQArpv58+qsqRbRicjouy7GPtdOwL1NVXk
HyPXGsry2ekvXCPXTbhPJrgqRrTiT80+ivt1P95cvSYmEzM3WmlJJTHQS7bUgxE5B+dJpH8T3LTN
mmq4pWh/pONFvappO37HclpRne0WxmPN+1OkS9pOBcVf9vy6IrHhtYDiK1aXxSswvwPStdmOcvK8
kOXbIVO3j65oLuKZxLHUxmDJX1ZQRTVAfZth0GPt1c/ARyZj0qgCIfRNjirIzeOSclPFPGLIAijj
8Eo8CP267vljD9h/TnfA59UrNrB2oFPQszK3w8fZ2kb+tTANaCtj/Zx47rldD+hJUSU1zuMQa66H
ThsKjxNh9x8t+dxqGo+misYG9wjQbmb4o6HQfbublWpnnsMkQDFaot/Gi1E54PUIXZhQ1BhvLLWS
EGUgKO6DdBV945p/p5ae/oKpcBfAjFamXXFSXVtsqroaHXzR8Akei+H2akTz8ho/toe70NXsgcxQ
+BLRHP9vqNX/EU4nHKFzVbuk7FVWtE08hMjzXQO3SFik0GsQyU4eF5anfuLlpuE66OP36qnuQwRs
OrtY5cu9L6pXGje/6HPH3sYzti2UNBdPsFb4QSvQs711/T041f8tgtiVAt1LHDZaN7CV40TPg+nI
saDMAZ6Cnk2hKN5Ed7EVJpYqFTsDB9ARA8gQrlmT0u68BxRoWAozeV2MBPrB8TBBDYzOgfK63Nri
jWVkJyH6MeNphB3uMK1T4XkewGIZ1dyqVT+iAHAferZkWR3cp3YOUPu1ApJaalEWvQ7MGwwnR0q5
wCMSx51BO5GiHjQC9E7kv6osIdp6Yf1VqftN0YWt+BdNX2Fs2UrqZQ0AGkQyRo1kVAUUPedd0C11
hPqQnGmXUAjGahlKhUdztBqL1hhJlArwCoPDufshU38/BhO9eATAmMvZKBjZxv65i819adSf2OQ1
cX42aAbtEgDqsfSXc2mKLdvGvC106eBblef1PQVJdul8kzrsKzwKyE9PgGTnxELnU7ASbt0FrYyI
eqErzC0YFUd+K9aU3MVE2uXolyCSywjDpq2IYshXntg5vazPGdnugtsev4q28pDhkSrY9hfHaWNd
T1ba5uChMazHECpKl64+yWKEp4hSOcZkA1qE5aw81OHP/wj2LnwqlBMYpdxAESuHkN8HbYuqFnUk
OAxJ5s2Y+cHavtTVMo9GIUUd1sINfON4NMvm7mpnSl64+Vrp3ziCx229QbqF++INHLkB4FDvpvcK
Z1ulK57/totTGziWTFPV/5G6J7aoM7ScBAhIPcPiMDw/rzJ6uKoDU+5LyqCMr1Y3NvArPS9dTMny
OU9M46WrL3dN3+ol/Xe2K+n/YBwriFDBxeg/in3eB8EDbKI2CGheDbQHjss8xFlgvFGGdyrG6aFZ
Q6L6hXXbO6Zo2jmR+ztxOccbbEshTD/5EEW0LsDeYKyGid+GABoHbcgFB6IegXQXmk5I2Ir+zwia
NPqXusXwJ7NA3LjOqw9Bqs4QOS+eQQPVXOxsvcq5/4oNTLyS5AtpSjhJhTqI3n0EG7QeteDZkA4w
LiCC8toAHOUPaiYzdKGla9PF4z0eEtr2UNmp6LzUGM+75kDsj49fOXlf3uLOCZUWvsDbJqJEqGot
gQPHPNpgOTqXCf9dzwyE81qv6RiK9d622XYxDklgdWmMak0fESfOzP4efNHkLkryiBSSf0ngVBhs
4FCWpzH7XkgcSVY5aNJ2Viig0RTeP3x1Phhqx/w3JBnAC+g/FDed4M7ASfNicoUF9Jx9+imcc/24
TNR9+DpM7wZVyZ3ox0LJncSGCMTEil4gjr60oL/wb/YKYSdfT2D+tU5DaN2wMCmvCDVMhS4NZ39E
iu1IexChyEVttygD4KSSmYTg1+C93rJKaVlqTiXgAwCgkFHLs911lO9rDMnlJz8p4m2QoRERVByJ
4HHjODGTT1OAGu00CdOG7F67dd651dqCuGD/RiB0iloa/eBWcywQqXHdSydin6beVkCN1qpUSJDD
sWbBrKjJu9KP2/1lPFST0X0nmMu+/ReA6ZuzKYBdzXw4XIX/KN+JeOJ03N3oGH3ScMK4X4whqnQw
W5uHSvzN+8daEd15Xkil+Uj0YMkCzUNGPOEctQ4Fhn8E03E4V/KzdwyccYhZ/nmT8c05bvn5WSPY
LCO6NyQaJ9uWmDUQrS9Z6dRfFa7j9ZvffDR8fFHmxf5jFt3W+vyf7gCWeTWW3gFR6aLV8EcrpqBE
b7RYONMllmhq1uRXqm9sStXtOzO+/NvQgBpa0DnhaOnReuML2+Sy3vFBeWtnSaxXSI9rNImB/u2C
+b0ZtqFSgiPkloqUqX8HB9WXB4IsxtjK5tpzcKHk1sYTf5mGufh0r6Dtwl2gxj0S9TkZR8hJ+8E8
nsw6wo+5hwqaI6Be3qARZR/zqODPDN6WyAmf/t5zuF0ptyr8aZAbbOH06N+tH+ViRMdOyMO/iyhp
fHJFhXt0GrScdoYygW0kJIiSDrHi4fdnDB4eo2lx8wEp6ilfIC+LIEv/ICMYdDVyfrg8iKxyQ3Jj
9Z1mm76KM3cXrxhNUAlOoFPTke6XejzPMm9d/lNcRaTir1ZDQ1Tpxz4GyDK+TLHl3ng+ZRWHhOc4
vyTOnKaXqxfasQMv9eXQ1m9n1FbtQEblXU4oNGJ0TmuDn2Kvhf/Bhyk38PatapsZ9M5U2rpbaeh+
OXAGkrCkDWAtcVpCsQLrsPTWP+6FyuzySn6TOEVG1Fck9yWp+/5Q3ZgRVi+KW0SA6tWuTDO/CuPq
86Uh6jxh097rQVcHxindFkbjdxEMB/GAWFrT14B4CaxrI7K5VfmfF0CbJJ6Y0IIPeiDp0wsmaUFJ
FfPuwUuKiQN8OWqG/fC+sDMMPY7AxJEX9JFxiz5kIQpPqiRUoiv2hOzhabYJWkX/UrqrTpexcUmW
pN37VX2KsprdL6aMDGZ1qp6GqMjxDK200A/eNVjPhFjlYSXRPlGuVflQhoc4ZEJcLsbSGE68RvJ4
wCHiO1jI05oTXHpA4MBIooFlPYC+1RuWHDjuB0PmLx60KxAIXqAwABTg7GigcoCTBCFA3f8GKI7S
o0GH0wAP88X7bLHhFL670Wk78JPi4TkzERxE1QBwdw/VEJ+O1jOEB2/RV5As1ObOqVPaF0YiL36a
n3XUxR+jLR8V0ibykRg3mQvrh5cWRS6Kzon22OpXbPQboGKuc8Ex1P23KmYWaYypVGe921WED4Ip
l4iOJvHBijeokkFeT/FtYx2BM8Keh1wjUuEDWakhZvqQACnSHualAaA1Fe6dCOtGv8VIh4UssEyk
rLi1+CLcDT2r3fYr8kJgHRZGp1nKl11RJM52YV4IBrNilWhubH6RIBjC6xsBLTHUl6T1t19Ng3O7
9Q5bRDZwOFPtaJICIP5+NU44jsU6FFOhxz/g4oac1u3kadOFWn9MB6vg8fI9dmfF8H5ByldoQYwt
wS+RhP9ASgrk4kQYOsViq8q1fwAP/6Ij7Z0hhv/r7nt9plOKiZEZPRRKEEOYEi5abpzZq2vE4qic
codUUNNYX1rrH8EYLnUDEh2MDku8QuCtnQ4tCCgrO0QfEWE2INfR2bi53ZVa0NwJIG7KQ3nEyS/u
wf1lyi/KP4yZOJdyac6KqYM4putrmE0o5dumhbDD7VJVW41tVejpXrP+6kEtMz3O2wGDKwA0atqZ
12wHrNulvjva8JrgY1LtgFI944B1ktcDHs5qg31M0YPtR3Plm5N16FHReo+GtAFkHlt9wrvrrQ41
zeHgVXzjS1KC2LRe9fTW9jI4fQcWdQtB7UGNGL7QgQExDv9uLBpMfMBHbArLz+ySteHhHbc+QB4G
hpQvYpA0VUhFRwMjcxmNkd+0xCa2DnIq/QrdyGNzMHkXC5Ftoxh33TE2hTfZ1OQXzf3c+Lcufx0B
Gg1RDETHyTyIgijloyycVEvTdhDAZWTBZ6fEVBmHpL5PIdZ/geatMTmINLuixn+s5jI+PMAJWgEz
lFz+lRBCZGHYmSHsyqy1BGntfVnwgHgYQtfTp+RGYcf7Q4iy+lseVgu1od6giWgHW8EejAYxn63l
ZqcCKXy3xS+qBKfJw/px73oagbQzk0vfYTDooh830h23sipWIwUJu92rKFhzOzz7MWEDgxNpxWpm
rKUj9uhisfTU2wnsgJnoIcfxn0CZ/uDzTvbxuAcEaPF0wCHW0NuVQ1TNZbj+hzLm6OenuQZPLvoL
SC30rGB3GiOuD1ttzhx0nyZ3oRCSF4Lr3xFB/1IvzX+AwdGqdWGVrNSIk4zbm6kqvRRQp51p6rIH
WlKO/6meIj1GBCJ1u+OOU8jie/ZfRrr7TtIGITX3NPwiN16mWoq46PbEoTdIY7h1guhMKYpRYhwR
1aHDYvkIvIw/LjtOEFR9xoEzrF6Q9/WxW/9y/Ahhow/36luQn921X7Xg6wMHfroKeP85Amh7m8EE
prYkzcqakJqK503NqiNUTHhrB74vJPVQ4RYRT6r0KmbeO8ZOMzMvaavfvD+TYJAWNigrq0GQYLxX
mZ6gDqab+Ipbs8ap0peMl0m9BXd/MkgPxPTp0x4/UHaO+8yjZjjZGQFZ1+zUuu8LGd+zMfN0OAft
Da0zAxwzj3y2ut20JNjXygnBl2rdca8dSAuVuldvphJnCaTfHYicI6qcX9QNTYHcQ7ZxxMauFAvF
9QPDmHRXiiAXlc2SmUZ1THlQfEc8O//GqTG5cRdH9LH17f/N0tEO4i7UmgF9p1pamtowm5zVz6af
t5L0ss1yUHUvu6j78K3QKRESBaCa1A6MZldT8/5i7EmzKA57VHKDlNOKr5xPI33LtDg0qdhZUUAN
uSG1ZBUgXpbCYQrdPt9azfdx67i7tGtTN4fNfz1/ca9fhkCkhzfmey7Yuqjn8lmaiDMQpFSYaHff
dVq8TM/elz4EUuNRxY8n21aCtNEIwKqsNBOChE26MDCASvpUaDMQxdzPreLvs35d0uuYfSIgE9gj
3tnQr79hF8oN1J0zfokK8/s8rfVCX8CeRyNI7v2lArXH2JJ+ecnlCCn0l6P2qOD8bR883XXE48ei
kNJsfuX337/A4rqJDvc0dUDMtQOBQ8mNVPNXQWc7Hwz+LZbG7ZEzt4IUOoC+mP268IwDJ/ujdnjB
xh4riVTpRiGFgTEf0ogxOVoqJVQH9RikjhdxBSDeXnG+Wx65Bow9b1iRkFy8WKWcrDCelnBUMu6R
5XYYTCuefMTia0E/ZFrS3WgdaVRH3Vui3cIUXSxMbh/K6TGoSbiZYR3xMSrX1ZC0WXwx5/gfzfZv
8iJF1XnTwb47sSjtIkEU5pEnDtVkN+/x0a1zt01oQLV5FoGtMOjNPnWLCoSkdMJMkj8YKy+enzT1
iVX1QP/hP1WQ01H9L817vhd20A/MZvtg2d5xYgT0dijau+tBDRTAJEc/Y2mTn2UlVnrDjvIPBayf
HF7JAKhvNpJvF3+G3FOkyEL78HIy0q8eki1uEO/Ei4zOgVrgRcS5Np9XJY2lydLEAcafVLQy4lZ6
VQdhbVpzufLYFk0P+tzNK1j5e7xxxovl0zGoqU+fxW5UvYIDjz9k4fgHwxu3jJNoc23mLxGYs0lP
ML/Fs2in9QV19rFv+91JVmx1vOD/KWySZJfMwflq4BkXTEE/oQ8QCaphmZUFLSSMXjaB+JrGdzy9
xmjvXtzzR/t1Q0nxk7cgtGABH+0zYbcbTXuCijgE+o4V8xBUxB4hWAx4FMtSvkZ8jkD7fyjgDjAt
rUQ4nCV8MRxJeHPviOi+5on6JuLIn7r5dCvfOLRAXvmBUyKS5L5tVXveWHS4Jatg4KrUCmQvPdPv
btPRd1lNf41aEuoBDy0Yw6LdSzC6DhIfqgxwTn2u022r7GmJQrLTJ26LpNMVNqNRb3Tydcc0dhVx
sEeEykcDVNgWFZV3c5TMzljpjvL7ZiuQ/x+NZrdF2Fxo6D0fNR35JuqtL+dkSlZQxwYiYzVwlrpc
BVQr2sMP48hoqBFLTLXy1V+ox9gPVZwe7OulOV6XYMWd8V7UCYWptah8WMNVj/rKvwe/rYM2n/ez
SIIERKPNpW8FlfLoBYQtqspvHcpglUIqnqpaOPihTURyeJjx74PE0LHw3px/n1iBq4TP6vQLoZdB
TVMD0kiVW/7bWbzBQBymb8vvk1Heb4JlgWkuUlQ9ZxDv8r3aBh9hrwNU1s83EAFAIr7F9E51PL/r
2vlWZP+ERPbJ8TmWos+3Jvs6xJEE9oFr6fIlHQmJO6RN6gbteui2eI7/EOaabHEw+ePTf9NHHPAE
9NaTji+nHEy5/vgPbWfuPFXvlR4JAIsf80+IlDpvoRT/mAnBMisaeRSNcKGToBV3Lp/ObazPemNy
b7Hgx0EdZXaVg6YWCUPPuHrEMS3qIE++HYHaetokeL24Vl0n8Ri7DFiZfuN9JKuogenjXc9KaKm5
ODwvn6MIP+9Cpb579kdm9skY1ouxUkqH/bOmM6N7qPfyQQlGU3hJZ7VN21vd1/w40PL5b0fw8ZU9
gl96HsvCaGlHp7QQPA06p+jcvjVwwkWN0FZSDdk+RWVuccZdjX0JWqyZ9sAms5SM7KrqMMyuQyK8
jTpiguDpc61jGSFnFvreE5p/gVUtPxRjnoBlGj54RffPOI+0OfKkeMs/cjoupOViNMLz1cLhHQ4Z
Bpr5ROUrq6eIYufU1CZKZ8HNeKJlgVxQD6K5Rs9KvivmOFFhuUj/eswQTC7QRD1pVGCJkDNxV9NR
0FU104/R6G0HVBmjCAwnPel9HPyZO71Vvk6dghxx/bWQIqkyxU2M5P8kTPehZ2Gx2dqeXeYdcR8Y
DcQ5hnoROXlVWRf0TJghEctHI70iDBaQwwGZyoY03rFr57w8xhAwNCN3w6nNj4yh29YDiP17Hs1r
obAhOaNOl24u0O+fkaG+X1iLAM5WxAGpMfG0axlo0q5ZZZBmCUhWRk7GJF5xWPZgYwPb2ye16vLK
yV8Buh24Fs4w/fT9veLIuIZ0uUeUSyui5qx94h5I6AgkwRHv6FPAch2ngio614xFHxGun3HlAjyR
RAc40DuMo5U4ra1hYlVz+lxt10U3vUQtwTwnVEnk4VJ1nPl/BcW4Qx0VUx9cP3r7j5TTbfBPKfq0
5cIJVGKajF4p7d3PTSOwcXEVMC6Z9m3ezvHn5sOtklHR3xbqh/9xXCwpG6PVEFVy3+PN5BE4fTEu
MyBGQHBOVcxwQoj8l9LJifmnTApoy3JvxtK3Zyjky+isg06vv++BX8pF3mDOQvXPOyJ320+eHGo2
BDrtf92ae5WnAIo5BTAaNR4d2hcihbPOS3pHTYL+7BiFiDvCmrQQ5VIqO0HT/l0043FyeGtYONyn
C83cVPU7yFZWdh/ux4Le8A1mLE/yfhpzWnr4vGKV8IzKm4gOmb4/sWr+dZT+5lV3vHjyxHT5hc69
y6uzJ12u5zKdtTLvkcWCvuBjtHfMXgU2vx+dImtLO/RBYhQLnZUlxZ4WqtSapYuE/l08UNe2jz3q
aKVRtNW3GI3GAcUAXRnJEvBcl9ZEoUD/DHTy9qzgo7YkM4G1fZXZy1t99V+QfRwn1ExLXT+raz0C
IaUzJiTyjyeoazID6/Ox+0C0u30wpSAy1MEy6LjG9L2uB+KFEFueL/f23f2fmBdjZmrSlxhlHFSs
OWlhHiKRG2FbrUJ4rF/N6aNiyK37yhF76mkMDI6nkOMiMGvADLo3Udjz2NWHFKFa+PVCf8L31ox5
Ye0qATHNixkkJ0DqLYyiYt18VtKe2Zd7wWlt0qk8vfvkd0mbBrtwxbU7Eu/W1uAYPvEFNjLMd79v
RWojl/94XuqMB1EOk6qNG0rnessPRvU1m2NiHui9BN1hxJpKNaoQ+EcUz35InkN6RkJ6TuX1rugs
rdDBDmrtOzop1n5JJ8EjPrWLVr8glROQ3x+Dd6vRxHMRYxIuVXwRpAOQx4gwYPfWk4jVBCKbHUJX
XN9ygRU1C5AAj6ubUlP84mdTZgw0L/NV+UuvQu3tZocTUto6l+dQMRyWPxttNBCf9BDDLQ3vudOb
hqyCxnFpEm1ZLqCqG0DUwuV7BJtIJY45ot0loyLKW3ecmAdlD+g1VDK+KCwXCujdOQenxHtSG6Zc
mf1Zg8DFN0JRdDBMBt37F4YDXALAwIctBWovqtuy4dDReGo5KcDZpM+jmDfphowyNVNjY+0uxaQY
8BpOh6aco/Ww1ncVxasQKgGf+oCb0svlIur0oTzvm7eZbn9s1oUyBhFoD516PxxUq28aX1FRC36u
ynfqxeB9gqzss0l3oMlUylh5C8M1dMuc0bxnhd8e+j5MrzyN8Ov7X0xSCj+pRETb+nklt0LgtSiH
fE24s603VeM9eeJY57UnFod7Om/KQ7ZZ5BJzHD32/gtUIATl0AJ2o1AKOeuDk02vz4SBsNNc2OUt
7vEZHCHx7ua4jivYeIuNdUSlxJNAd66yhzER+femO5mQLuBfu88ivgGmoagKBkV4/kkcqKlvt408
It7ZnYmuA00kz5T6XW4fg0zOHLt9h0rEwGd7q/lt5QtfZOjC4XcVqIi+BWnV1Za1EfPCDDnwxT0w
4yffl/XSxqV5A/difxJwK1i/XxeQcHGKfITkZdaNHxl+YkZr/5cQY9UpJ8d2B3Lcd+IJ9gfpkMny
d/R9BQvdAZo1PFB3uLvVHM0t5sxWCqIpIxitob4jaoFTg8NE+3Rojl40ijB9OSbeZNrYoysiTSNi
YrKGi5UZ5/nWcfZKqqcOsjWuPkRmvyw3Gs3xnAfaPNb6oZ/tFVxrdhAhFy+HMd2C4UBrPsVG3Mq7
OGf4IpqpEuWFUHm8w7lSYsSxV5enHVscp7EfsCcrH9nW2rQZrZz4mbvTTQgPrgC8Jzk+qd/nQBqg
83qBN6wEn7J87qBpqQ7BEAIVcY6ubmizMJBzaQHDqYuJYC8u55dj9n/HxjOD3DQf6sIGZGVyycwJ
rUpZkChkGtrYKWQAnoAuaFFj1uXcxvqAL2WZ3Zi50fiZFUkjuluAF+wkXTxQCIuZzmx+Ca5Bpx23
hqnr8MPkymT1tJE8XWEoETJIRA8bvDXj/TmTayXnfXpNpX4Tgz+08Bq5ZAKHCIH/rkqzaw3wv4p3
po0d1BngCOH5Dhv9CN9i6Qcbyi0LaOEzjdxx57LEegBfqOX/tDKfUfZ3ZCuY970GOVsVqqmb8ISU
/O7+N+skarnZxE4HDx2GLqwbrpeAwogLQuMJOf3iK/NvoNxL7EjN37XtPvTXz0KlZ+6R0ZMpcWNj
m4qnPOu25BXbfHc3qEC4T8C3xE7XMrehgKbuAq4OYXoEEdRYWiV+Bc7CNVrMbEVXzPV0kgHlq+k5
roEImPTnpVuV9J9uGBMKWX2/FDUGSWdwHCnxow6anWzZ98KPa2jixZUlPemR/cJw9vE8fr2/+aVF
TMQ/ed58zC9FFM8CrdDb3xIaH6W22qcwVpdXpso/umbc/wnnHl9a5ZxY5GhSp0p6BiM6w3j7rT61
3rE9aRaFrt4di86Cm5j2ka8WApFElUII1NTdWutudxqCQh1Cij+7Q/uVLS957XW9smTOPwW8TjHI
RhXaklUaNwMoK6Dzo2xtKcfmoyGDJ5rkampuCpsY7Ay6/mHyiMhg3ZVSAFIPkpIb5kvtgDfMVR3/
uGP/SK9Lwwe0rxCBgpDUMACjeVkRn+ArzldKEcf0gnhqODIoDOu3GLUVPudeCTcG8JsRym9SnNYr
eI48GqzSfv6Yxtd+w2xH46CKMl+VW6SNQ6Us436IU3zRb4CeMyrc22lXFQiO1HSwZe7AV7N1LHLs
uAQq2vpSvdfchbsM5f0zPYqkoaQtLgnBLtL2mOCqH5YvaMy+7OhnoB3x6GKtBEdSV/9M+D/z3he1
+IIMP2PRTJnq2aeviyWsnpBZkhCUa/r/tj8cn1hyQDaaWGNTNoE5bOidHwyMV1/ZK59aIcC0R7is
KHPUaMGepdstsjAf59AevsR9blG75J5TyRj1qawICWiq/nVrkH78S9FkEcz20zQDz1LcUpJJbjCp
a27gHDcd1enuxMcnQXbmixH4NeXsiiw8abOj6upwKCzhgZ8P3d/wunpBhnLHKcp9DvXwouUsxkXB
Fn7LndU0tq9v1E1hzQb+UNKxhOMrSrYwnmahM79tSsttGBIYvydK2dTU4jgW7of+DWSo7KaDCGbk
F+X+05SIqxXV5LbHDAtNxQge53bv+LEv57kbCqgBC7o7gTaUAG/fsG4ozLmjFSepN4HZriLbDo+f
KqurYUa19lJpRJ0Jqhgi3EJBKKTbmxTdZu04s4PorxGAy3WaQQ3RaLtoTU/+TR7rHMoBOBegxmlm
qb1PLh6yVBXUAOLhDXUnu1xNk8aoHA+zEN5EgZqLY2oJz9wow+r8qbdijq5vb9F/kyrwg9BIY9fG
RKeQ2pX3ApBaYky+CrTo5JyLV9kLYhOiESxykr0MJ9MEtz9GtG0m2tlnYR5q8XEeIxWtiagFp91L
JcTwwqy535xhEx45T2EP46NDKbhJddnrY//uuginQ0MldcWMCfOS146WZGjO+szAWSRaewURTmK8
gbY/HzuEM6rHcuxprZNrhoYsEq6Mx0cMkrtljd2Gss8ndXuC4mQIbyMDqKpxZTU/r5zAFkzprZN+
bTY+Y4A/z+hKnyKTR9P+x/X2dmewJK83FwFU+4VtPz8HwOgAIqQKjVcyFKlFJxNSL6cw1p15pm3/
z8wSmxsSWdEjct640vvW4+aKV26WidmqaiYBtz+R7VzxYliXIusc+l9b9HkfANgv0CqapTR/mVNi
aGFcqyoS1rPXImR1bTWtBrkhvX9DorBeYJyY8EY+Md1Hs4gRmUY4RZvugoC4C1Vmio60L04u3WO0
aS6UhIZvIKzgzluUn/yJgrqo4KM6y8PIUY7rJUfzLfC7TNiD8sDNNl1BUl/NEy9HB8HwmNia3r20
5dbgC3Y0sO67gMFzZBVdLWWlSv0s/GooENgcz9INyjeGRoh4j2Gjh44uJaMMWxmri00KHzqOcf25
715Wb1HzNEpQqr2K4Z63qTcQJTXahp4ne3FphLXKlox9NYQQZNTM5h29LF2Z1OMXJpsG6K1BMsNI
DH+EoG9XC0FORRzqHxbF/l71CG7bUxYrisDgOMleo2U2wAZvcI5zjp1aaE5UN+JbVeqOeNTdnMB2
YOW2tPIIcdFWgEMd2oJrgKu2SdN05BUApCPskX+h44/7Z22Wz8ofk5gGartMBHY/k+XXIyN8H/sI
2s/nahLfR37NQEh4uM/tFH1bprWcmIWNjK8qgGdIjeczlerlbfD0sBXzHlAFsG/GEeLnEviGn1uO
16Yc34TEsz8n0YhRnp3eBDOE3PBue6/XTWqfcHpoGO+GMNHjqKbY7f4UFGRBUyxvGHdcSK9oXroA
L7Y7/NdYdUYHber8JboywruAodAPVYspeUiroLcjiUSvUcPe7QLOZ+3bMha3ckgSd9Osbprya5Ut
g8UpPZbsnGwHcTxT7SHTk4+nEZk/J8l3FgA/HLvpRzvDh99mMAP1Cv8Iq58nir1hlmq8NhjyrWPw
4uafW1ol8sES4w7IWvuIAPf9VYNahOPW+aBwgSk//IGCmbT6NrwCNwMp99xT8uV2Z1gz/g6O1XEm
QvgoQjkDQgYypycUvM8vLtzunL4tI9FXnLwG3UxBPvrrcFz42EavxLh15vH5mV8Tkt4YCxegfcjj
69FT8cHenAnXlnsIKvnM5xzXmK5WXihCllu6PB/ZiJYQ2t1Kj8yBwmShGasSTkUM37ND1SlAL1+R
WBMoVRVidtSmdlnJxw7vA77Ye+Lfyi84o+C02m4NFy+YZf9uOrSbsr2xYdsqqu2KmqN7yz/6kf1w
eM6Y9qadNOp22ouY+sl8Y8nYPsgiXeEbVrohXqWI8Pw2HWq/9hESFqbQylva7GxnLOzuqy7XWSYZ
Rh/sbMs6L2HtqtoLTPKPXy0hgekWbMh3GKM7mp19so9tOMr46F8ClDe8S8bMYbArga7fr7MmD08F
ttUF8NzKsjvR30Py1CSIv6n97nKCq/q1j+dPVJdRq4+JFqCCAEgruqOrWugA1SSWf5GYooa10KEi
/EPNe33hZS+fLG2q7F0gTQ0FVDxVhgEhzvJlt21AVWckp6bhJ8jN8emSCCH4mchziZjHMK2Eim4k
bIarY8A6WOesVEY/D8nVw319sJVwYf9n9g/h9DkiOz+X8uo/HGxfqUjPgdzR2i7sfkbMX/tXWMew
+9CPr7AUmK90IFXf6Ebe49OXXmrzTnbY6ICN/r0pykkNgQbQyAY0/jM8fiqxYrhESAAKHSDaH1Un
zJ5JEawvmUVmn7YC3tr2U3yBQBOsUAZDvIS2yf2h5v4YH8axcgTu+H4regb67UbQMfolrRWA7SS6
Qx7ewKkQDxVvkYxIvz3QEtHKEXSD0Z+ESf7i5+6YwrtuH96hjZixsosnFTo0bpG6k9Txv98qjjAw
SD+vaDC2tW4TYvvp6NqcLOc2BXU9dFm/mzGRJ0OicPZM9/g2pikxgZvz131ig7W0eU0v+ewL/wRo
02bTX34y+leEhf5ifW6iaTPD5O7pAB90Ze9AnnwObQcRrQRlQMLMWzfoVuxSwvZ9KtcMTqjWA/0b
WBICaU50r8KH+3Dw8mG0jZiD38BXvzWqHfLuPzWopuDV8mjhxwPI38c7MqIZo+no1755ClvxukZl
mC2+BGR/0WPKJmFhBqMLJnULTG9v8Csv/laHqTt9ICvjQCc5d9EIE/U2gxj+Mu48Ry0JLbQFjdBG
4uGsu5ERMefl2Ryo+CT/n8JwHQ2mcjHyfgV7r9KlicKG5pno0Tl0W3kknWOSVmPpeuCIECttcBrR
mJXLEbjtkoTHoiBFuX0kbu4+bJpdXeqsZcg+LK8z67cEtSISAn3d/FvvVAqoxU8IKjIx0fzcHQvO
UHKBVHEKQlQUJp7KfczfS/ZrsNo5pXIqn7mcAgtcsWsiU5/tVa6AystCIQhjqgUBskekH2cgw7KP
deDo8jH2Rxsg8bG+jYCrzGbRW/URYpSelzg1iDc1Uz6BksA2JDryai8T0+H1enb7Yr4sMRZUTWId
YKEVGt9pONLX1WYtJnosgLS6g5wu6yvVshde6ruSaBr03I4Tjxx74q5Y2qT7PkZhCMsetT624Ppb
4U+x1rp3AnApPdl48FHVV0hnM5nnddGK+A99RZWRrr/6MxNX/e+OYx1bxVI0NxpPUJulMHGjtSKV
fvZ2Bsu+0BFtjdbpppGM09ijRkxmANEv5MXeXkXttfRp0af5kdu2C+lDxX1+i1ZKlyiEzaU/aGN/
tzUdMQfXNvcKp3LnNOejIRUPXfO4Z7rCF7s4z9JyzXRqNTFOr8t0RJ6jI7QgFL4UWjliZmojhrjk
DXum5BplG31tn6OXtrqtuMfP7cVYt3ylJsniJVMJ8/3aVHNmp7MOM9dUrd6kSStWkF0MH8IP3rnp
u7KkA1gP0f6t2fQz8fZEiyKpvBX/zFABteCRkGzFxPifOsTgMjKUKvH9Z/bLP7PZSGm9rVvZVcEV
UEmUc3/d7ULyePLIi68Q32sB2DArbWtGEGXySr1m9gDw1NZILpfDyLDHqM5NH6/Z08rSKZh16/rO
GmgR9jA5CrrZ9nJouP6o6Ny0Iv1fBXHrElDvHZ37VhT9wViH00cnt4ho8E9tdOkOqvt+UqEEdI4L
arLXUR6Bjhg5hdn37+PfTK++xCf9XJ/io9I5BzCLn31OIG1V5X3K8JKdOrj+oJkQBqECjw9/AYBg
ArqVxEwiLJj4mlMjEfbpYb6/QXn8H3xMsuZNx5DxLrIdv/gua//lhQtWOlUnByBBA5JVgqLQpdD4
bmbk4KmYJozhxeaynbkvWcisL+YQDS1S8FKhuc7ln9IMwFEDltCvFF4Z873ZYTsKKBM1FNwAnJvv
NoCQ4uOp/LEOK6geUJtH0oQn8d2l+040dY89VSc4/1UjIBHDj7eCcLKnh43nfUsyK3FtVoAHF6dK
QHdmrkezZXnh1r948AHpBYx8BGythEXHi8l2qtxnmhf/kzqg4g5YwrPX5kS7bVFVmv6vh0jyFs0p
mqx3AP+T7xCzF9AhIh6OKo0AVacTIWZMBZvl1FB9MfuyLQmJL7IvgRlp8ISXnxHeaxjkM+tVHY3V
QDeuB7/cGx8IBvi5FKzAS9xpoV2wEmPxD4nVhB8Y7+zNMAN50EJkk5sGnB/JAwkkrh5o8IAcUdwv
rI0Jsz3y0hOLeAIrhjqBX2h50Ar1HDK+htZaDZdEuDpSJdC7zKATEArv2D5VKiqfYwWhw745ydP3
BtlP1Fds1VnLJSt2WXS7ZiiPNoE02OWh6UR/hXw2/eCJcuRshLHsrcTCHRcZbBIGJKHmoa0vI7Y8
/A35Kuid+iklha/ymArGH6RARd/LGzgqSmQwbbVfWw5OImsfVzSE0juL0CKxdzZWNn4yIg+tK2h8
FZjlKtSaxOsXikGQg6ErkIxEGoBHDmK0dtl9YWwJbfI4C7qAPi4FtH8aNQmCPAcEUm9Q/t8vlYLj
QmXuzPGo+ZGuJCBMGSmTJaX29oH0vW6k0NoeUpN2oM64rMSuGHBWEzCML7D8xUIBzDeoWLaMr3dL
CeubdUxohoOFePhY49dXYSYCayqJtVf9+4kuhL7soDOJF/yACzlcOhMKqUbHEuRFzVkQqTIm1x0g
WHO7V+MqpNknhxujHKxjUQX3Qau+2Z7PPZsWhtjWUNt+TkiR/UNp/IHy2mM7BIW7noeB78DwE2xS
9LP5JiS1ShzVhdfI6rC/fU3m6qFO4Sj7a7hXRPu920OQUA47M+nHI4qmpmgYviBSc2SeiJIc/l1h
LdrENbHONtYgfAKz/H7btrMpOTQ7BuWJNgeLDEbQr35wI7nkD9XzM+PXpaxAhVMnwwVtDISjPepy
7dL6710binpEXUmqn+RULr6sLYUDGyf3fpQL1hieViU9zW6rOC/z4NMnjsuT2GCkI8c70Xkm5lxV
135RPai9KWl2SRQNcDXLKVTqC/8tMma+jFV6ouK6EdaCeyQQba0Q4ClGqV8NUPX7tEikbjBsmf2t
0y9mVgakvhizjbQrBHsl/NgbOVw4k+kq2RsYb7Cl17EyAYNRZ7PPfXFq3Hv2qP0FrrJ2B7W1gMx1
GPp/rp2To9tckwGLf2WjLNI/QeU45sQixeH52xlnxauwBH6ekS1ksiaid/jRHSYC5TaOguJooN7m
xeIaRrQfl20lJdIQAtQTCRUOmaIxqy3FRseyZS8IiJ/s+xVk1Sb/DUi0aGgR+CDzj7jug1WIuQNJ
C6hxSIT47Hncbv3WWnVdLOwBX9+BnTwHZRzaq6JUMNWPM2LaKiVYZAhMCdg0UHFTZT+UZEJrNnfn
aqk94kbuk23u4rkcI+MRCXIgYjWBmkCtfYHjCd/DNEHEDWPLaoYsigCfs+e/in1jvzJ7KBKY094p
Iknf2KHEkIKUDJiLCxlF3UZipTd3+j24SZFerQykBs9Akcf+sZLjWNavF2xCHgFxxTIDbodRWiwn
T4h+bAp8+TOoUukaY4k+zEJGDi+jqX6otwljLpf33hPPaoJ0j9J3XfBdbBk4ogAihtdia6/Ew7Y+
MJBzkDQIgBb0+gMQfimlL2HXm7iREmcsIeKHpe7r30UqVcKjRudrD48RHIh7zcoKRitsiLCylS9O
0Co44ip/66qzDd9G4CYlKwSfEhKRprhOvQye6hpXlJmjSrGcM71W6Ov7yr4krjoBw3czWe2F9aKr
HrznQ9P6xkRjo1dUWZpKtY8k4/yGq4BGMCZjizLqqrVOoQqGpNmlyJdO9qDinFjdqHk23OeVZt5s
6+Ohvejy4coYJeWbTVfv4sODIMjjvFoJqwSW/38o4hHcyETarOl2XMmCXaejHduDawHyr3gBQhzt
8lo8/rBG4q0UUD429pj2/5fcAw5/zF+A4UAQJMILsGZP/enfhGqBG+39sVPNCM6i0ai8EflMgsWw
OR22hZMrxGluo9+vZsKt5ijrnpcoxPuiOVWfgNUBDV0/UILAWwhGyAeBtw0WBSG3DCxWPXmlLYFR
cuhOTKX5HgTvT7elDdsaihCT8mMNjz/9gEnOO29Yh5OG4uBGcBlN+vprdA2J19LV0717TtIJRBiu
Q87iLW6a1cTGYoLnt36ZwwLd27XyCe9NggKruHTa2OOXv7C+9CwEEF2dvJHnXnALwEvroqfnv/2x
pa1z7wUaWNmU2bzl6Tde1yHf4DfKrwfm40Ob9jUU+vPZCNHc+nVzeMNYKI3YTeucJAiz7+gq/Rrv
+HoZ8jXsrgaE0Bb8tpOVcAsLfZa0ZFYMLYq+OB4RRqwBEJtRr+Slk63VtXO1Q54E0bd5XN01VIna
6TtNDM3anFvH0JuUlsVoz5Wxnd5TULvXQnFBYCic5Z4XibcldC80bQHZnfqahP07Tek87rb9m8R0
YJQQLI6suuirHihw7+JcITWENgb4sCpoaVL1GZH6silxeeYXqYI8kimoAU263MWQGVMefLstV9UQ
X4SCyShBE4sK9JbepqA6wVGsHeJZM4qpTzVJXqTCA8ze9knC1yUDfnJsnk0Darg4ay/NekLXcQVL
4Ggp3w+Yaj7NpUGrmpipMdu7O6ffDQkCV8REwZtrwqwgUd+gvjlDKNkAHzxDne4JBVfQ1A0menwj
N/pqD2QBSUVx1mUTSb5fwP/l8UWM+KKzEDWTjC8glJDhnmnwiwGterVJoXHHGyXza63cSwKjFOHS
TEZQAgNzJobBMUEbBvupjKrAJIX3bz2ovkAMXWpFTUU3DnzzsVIhLib5S0GjZeRaIDHwa9kdiIOw
djlGmtLq1WXyhqQMNtCpB8Vzc6UxSpFIBKDhgLyxOPPcwUpL/+sADsCgCrM0tWoMez3jXbw8vRBV
zlBNuZDlifmAYf3s8QjH7gKruw/8z76pRRJtZKC1RAZ4ww0FnOeYy0GVhGLHZAzjZhweyi+fJ9GF
b9jyKx6Azwy5JVFa/4grrYCJ5w0nVKEp3Ztq58QG6vrraujZ10WtChuyNWsh+nS1aZ8ULG6RVLBM
ivsK+hlmKz/AfeRcbcLDBD+Hucc8qblS5WifoXt7lx+u5TMTiEGCoMowhNpJY4mixJp1pkqZpvK1
xOSA76MoAxp6F54utChoJ7OfuXddCNdNJ0YBwkhNjbuDyHPZ9u2SJYHQfMstXb3GZfYGmbRSEFRi
rb7CB6BBkTcVTH9w149He5G0bNLqIDT4H8mIYtWrfq7AClyFbN47uenafYS6/zzDkDUTzgPJrvzv
h3ul3nanwCO4Gt15MiWVMv1zABC1mPi3UPcE7sV2eGJI5k/V8XzJ34W+9sMtnRvpfzr1j5lyuJqr
QOoKJ20X5m9kRUGb9vjI6aF+c2TRxNVyHohr1hcH1k2GrGO5f9b1iPBjl26HtoC3BYfXfHJ/ZqLN
nnkhQfun+5TOCJ42IXLc3OqzyZVyg5N2Qgyq63n9lnTgwXEMHERsZjRhUXSSL7fgG7vzJ2GTjQMC
Kxd8wJbO04lTTc7HU/qC3cth7SxltgDCa8cLkxg+OUEHLaVBUBhHqw1iIDH+0FilgsSbzOtrpF8t
XBWdlBTzEUSLGCQbx0DYSYR0/AeqlmV0Naf6faxQRmSrO5LpZVxga7A3Zhr2+dYptnyxiUZ48EEm
oTPl4TgCsza5bi4Gu1L71+AzC5OMJ2BsU/ynzAmieuaPPqyj2ElclGQ6sbr6ojRCbu8umBdebK8b
dNLkpw4uLSjKlM4vbxjD9gNn8LAQJJ7wn2o9hoaCZGKmYtiePNMqdxKSDgL4+Jts/fwHHTXcO6IG
vScmVkhwY+19a0EyaalAOJiX+qzqCg+cejHWW5zk2f3HolKz0FAObXDfM/NJGYE7LgJns0DWblPb
QJXrphdH/X+ELE3coop3mbjG7XZaGhVBEeuFKmo6WXK8Y087oEU7b2ZnBesVeFHyYMTtjxZbVSTo
s+4MD+/oZQM+uxnvZS098VlKTydRfcxMXybHY1cYWdw02ksASaK9lTv7LrXvAJHAL8nu/0dyItI5
XtFWOC4Q+NQFvPRelBtaYIhiHUVycNIhEydb/ufP/FdjS/MHdCdFu6d9Hq0vQY5//jke+l6RxEyT
HmBPQjZccwIgXlAyXc8ymImtysiepjBipdxw9I3z8JNHiVbxOkk5xGNGcRrp+n1QZ6dUh3gLl1wj
R50HKwTEvhUFNMucIfgJZKbXsBppeWPkGKCFkfHoU7v4PqBmI1qL/AU84mw7LfYcvkH6Hj+2kPqB
6J428r+ILBkgY3J9UIYKbk7//bSmfFkh5UPj/bHFfNX5bfMqcMCZBWgtIuS4iJhryDzFDthZ8FO4
AjAIpiUd9tDi8lHNuzq9KP/qds1HuSCKy4zG1OgA1SY7izKyH0kUISLO9/UNvWnR3oOSMpIHKRV7
ckM85jbjKGU4QyTH2AxVi/IfiUhD6ydJAZ8GvV/i6MtseROXTfBZR2q8kLC7Z+picoimWs3xBHmD
fL69+2RApHNg26AzXm1g0DkJlKkV5pAbZvv/npHxFVKftjj5EtuDZYPc2panmgY47eAfnQ1nGNxY
6mD6FBDCTvQ8PBoSThwCXt8J/hVCKrtc+4biJNHyXd1HvB5MvCEcos5+qlZjKut+uXH72Fw4+DCH
afhs2dzL/qyScBEL9BltbrlgM0QluVDImjMgX4JoQc8Bo/tJXOirncE4kOaeSnCDkenn4UtV471K
HQpRHJWY/1zay0zeVlFPitIAlq3Fu9okXMrdceo+YO/S+peeOE3+nvxs5E2LBJsjX5vtdCspCIAF
HaLkMq1Mjj51z10Mg75b2eNkKHmrV9sXLr5+9tP74pWINfe73O532csXv1ml6Krz2aljPtUPu6GO
Rs+JuBn5K8eSazTTyNJqWJZ6YklnWpGZjgMb///DEhb4lYgaR/0B5pej1ebWytKRT6crN0Hjp22W
kFQVgIQk65EsuEbQ3sL/97Ilv7AxbkmDNeJNqlfzagaiWZ1JC7pa+X0btsqy1odUW17jpcRDk5jo
Pr6cJ17CGb1RlrQrvxTJE2DmUk/fjwpVZaj9gKUO9Pg+r1rG4SfKup1svadgL2DymdyZV8/Pibhj
TGExW0fcFGAAJRTLf6LbXVrx4A862eJ+mZLo1SubmizSiC662BsivW6X5D4qIfkTkVQbfteVHtT6
Rn56ZoxdJ6dw4es89QM2JnEuHRLfRX33ell/uHmVVmpBLd6XDsqhiNZau2sSTjvMnw2f4CCxFfYj
4MFezCe8QtDyXGidRD5d3w4dSSM55YmdOouDxmCblQ4ycu3PRVK1DgsJupo+T9PqCtNcIZa3kV/2
QDW53PqNg5Qg3qfcS65P3+7NbtoB0G9JERa4cOjOxx8kg1huHH0q9Xj4EhljGYUck3+ABtVOO3ve
bZUXJlU5acrDa5hRRQtPpK3HTOavkgsTbAUGqeJi+R/UMiaBqlXhkjpx5vuJdMQteqbuomQVX49L
lVmqffcN9PXrUZ3yrC5yflk1zie0fBvv3u3DR9CKqI7iz858Xz3kRAWUjD5hYjbLfIftWOi69NMH
eK8j1QpccJUTCE0hGcHVnSuJpui2EWj6vAIelQimfKQz/HXvDclPVZVwyW4KwVm/RvDq1TWp+Ec2
ttO0LseWiZoMMEiv4+v/cAwjCyUm6Ybmepi74iekyXxQ4rhK4bPKlQ2eyzEFpiAJYTQwq96sfFIc
8JOCJNAAIrJ42PvqU4noSxv80ki0YYbm7eIfIx7dNstmyGzqpp6irpjBdpRmqm4iELqg1rxn96OL
38rX8lM4meD6elHK+gSIPsqumbImvZYuglUo6aht40cy2PO/pOq6+2v7+9lN7qhkV+YQmKGjThTn
tuWMPiRIm5H2I7xVtAIjqYEUeHwSImio5o9wSS7rSeFdd5R4SYtRCHemI71+Nj14nOywyYuTeuB+
clFR/uJbsH0TLTmoZW87Zd8qKDRyC3e57Ttb/bf/gY+y9bY5GJdaHte0ejz6UkH+/NEf5+fLPw5Q
uCa9TcqPFKWQWB2dKB3c8LOf3ejv1b4+eJeOieu1CXKLICXiJkto1NnlPWRv17uiV1UbROQ10qm0
kmwwBVEK5ReQUdI+BovGOOi87dhiDisRnawCplbQvF2HrbXteL9VzsW7Zus16pwfBrftOGdwewPk
uHqALqBOxfEcQ0rzN0amq/CzmaFDpxpQoZK/s/HL76fks4lXH36UtL7fLHB5TUZC+972RQA1tnma
3FUFR3qTD6bgvE5/fiuun6j6taPv7DO+j5s9e8IWIx/oKzOuONHnfRzSz2sbhkL1vFcbDW0yydKy
if1XWn5OlBdSja5RYTybWjZDLTLIT2ldKDpSKyJGMnMl3cWfvMTgm3wIjUMA4GL5mHq0QbDNOEA4
ALURZxenLpCHWgvPsa3WDz+jk80Gp+Tam6OaIf2AnFUVPwqDkswTP9kbCxEwRCpldDQyBFCiOaSd
TiTOUjyLkauqCmH+hZgqAwkf7RTlKh79CGZYIjhjKvO/40JeTcI/KcMiqEe3PCZOaPfPVtqZaxkZ
uAc4iVFkeMfvHRVg/002DOcsBEBrgHRz/xrYXz1aNxKH+tl5mHmRRxLwyKqqG+FEoAOq0DaJ7rZK
zuGWEvEkJpym+SnSHrcj2NjRcUvfoxpLj4f5L5QORbuxtDThRt1xDrRhBWA+n/Vy36JAsoaiJldE
jcgpnjVsTr/vHOBbKGEZEhMGaHkOl8KS3GMnhgrjtqBRZbz5Ot1Xu+shM3vMZGMg6YRtRvJ/gSou
Dau+6vmANEs4C2kCrPyIOdgGJeVr8CR17yJuJGhIFbjWoJ7f2qJq5z9COQDKDVtuTKAzwyvZJSdW
TxJxTUzLODnAFzpNkFDn+ilicnqJY9L3To71WwoZ7v7XSalHDJm9cxN6LJH9GSD+GvV8pDUL+pr/
3NUyAeWAsj7y859p6CKGhdnHTeYAqhVA9ai4OaJly1pCp2gYg0dc+YpzdXwfwte98ZlfjeKZuizg
YucA9eTbojHxH4y2wEphE/hzcZoABK4B+OjfA9uiguQJgAc1ZFprfZtqKQxF7w7BcUMaiNeOV0gq
EYnqaKXyBDMznm+D2I3Y6mWkuBpqksba/HcsznfwFG1YLHiwqHVe9wwfLYGXCXhoQHAktAOkqmTw
Jqlt9pGSsPQglfrfwNdOhL/xqBUV5oMm0JFQdt7uAyfJACDpixHDUpWCkrkONZTbgOL6PdrxqYiw
hKXUDAcfUoSJlQLWbfzHhG/YFV5+ygg6yUrrkxZPhztJKlXoyZGLjJugfdQZ7erF9Bo70AY9LFEj
SD4ksocFeGNQbND+pr7tvjhoiil9Z647bvopQzcY11zrebqPI3UF39EYsfvS0SySKS4RAJmfoaAJ
v1bP0+wpMWQ3CmTGSCJ4JR+ss9EpWLq464BlLmBk7Rh7iEf5W9VU5eHuC6qjoU0L+zJCUe0dASHH
IlfTBEkIHR7SY4cVfrFlVlAfBV3TmQnuQG3IuUKneYskKF/tABuUQUgEc/C0sL6xoNWnLFYBHqdJ
fSlsBOIN7h1BmiTMLmagorZhw9tYjw+xzJcQaJrPT1ak7Axh7y7vX0yqjWuU7rPcr43chkeuhl+R
0uoRtqITJc9kNngMVCmZqUPoxNPboXZceoN3oWS2NZKIBHA2BM+bHPRkCDJr0LIzJXcfmvSWI/o0
e2U9lHsuoJFEYtrUCuoeXQnrtqHco/3n/j2ZZEsXjvSomT8YdjVUDvs90zSo9SBGqEkS/ocyiK/5
drwHeXI/RuYt+b5wXRu/ZmT5RpyazYxiD7hLUM8nq5ldFXoQGA+b4zMeYC8GZ6XniJJ5k12X7oDR
4nlpD6570dhYD9ryCbxnrljyZSqyBDmWYhc+Dq6MdpuIMXI5QZai9+uzl/9uimrkBfz672yrDYgq
I8tyzuOcrmRGYF6bZBk+d/QMNUqIjU4r8xWSqpV3hkx+vwjzeBOfNQgSAQ0c1bAIx3LNcz4A30UJ
XSk+Rcc7V+zVjEENhTZSOrR/osk77CvTLVstKy9GGJ963hrUG3XvbYb0eL7N6ZZG4yNg3Alv14TK
+l44JnyZnZ3xF7PHXvIWGqsFbrj9gfmwaeBD+cmvg0k4ql61wDYRpAErju9kSAkRdtkzkC0cBuWu
79zPPMSdbLju/Y9Wj2Xg4Wo6Vb1Bn3b8NW5zi/xmnIE8ZTzrQYMNuFVNfvDMUvNkT0i1KHBRhJrK
MKbDk5i8j7vjA1gHWd7TINLUrcFyNXkc9ckNBbqmq361mgMCIPjV4uAGE2Eflrz6MLavKh1ffOQs
5TnLOMYX7OzwjC4plT8WRp2IrJrNAlO3/vCvLqPxjFjyPqtTYwG5BNCN36OgeoAeLNUqztqOr+aZ
SYKG9J6DfOtkABAhXxXqLfveMpM0ZCqGecIkBoGm8/KbPr1aWlQvyAfLRveeJLDckLm573dVatoS
JDhTjI3ZAHFZLhYNa8/NSfm9jzsNdJ7ZRmPfYrDfZfD/IxyxDKogizQh8bwTM4dVy9El2+XDPRms
dpQ+tGyF9ttcoVUhtBwK2mlwTTMgV00IVIn8Yxk+Sdge+vJIH2IDuvJ+hVAjvD+gF/A4j4w4GWO0
nKJWx38K6owigZg1D11O6f7GqtB1PBGS9pDQb8u4ksPUnZ6U8j4YWsbKB9KNaJOu0cYq2jH5ExoO
GGBr8XSewnitscwGCgRautlfZ30z9N/n20hcO7hfna3MnzwVwPLN/Mz4TQ1VsSpbd7LtalZoHe1G
Hj0xx7bkNYdMXdP42lFeqrd8gKyDeqXMdJO0HVBhU2MwAhSvIHbEkuaiTmUOuuMAwPp87YF2ZjEo
qL3X1qMeAx3gxTC18HgaGkLPosZE3HfOkgo4+AWFQ8F6O8WxX/MoiiUZdJXjyVmcrfKYkGoHc2jA
OQB2bjmeT5oDWJZb59MD5DwGPHYigN4MAO3z9l89+VR6nijGDGOc2QG1xGSlQGWWa/XVd6UmDupl
oog5KLEGejh1jv0zmrYFuKAppn0wgmUQrV8TwgfSLZvWCOL9w+ael63jnftWSOAT/qthB5ufHpFV
/j9DACacWyFZQCqQnP0CI/0jw0pDv0bz7vr6PovKidzzEQ0tJOhfAfbJCTDJwM2WYzdyg52RcORi
ZFFJidMNCz1gNOCfLmBnslElRYyYClI86EWuQIC8GbV28KixN3ganMUn3HZSuh30WlPQFZgk/5X1
Y5i9EnMbv2nHFCi1Kk/U+fJuOGNZrsVuQyXHCFySyxtbliYneK2RIinRat1hxGGYlb2456YuKe04
qVqI4y96rl1sYfGVc90gWrArOuLOtYjuZ4sEVg/I1cxHFzVoGxhajViOYTMjQs+65n1mL7akyHKv
N30ZPRMgPA7QqAueapQow1CjohKzBv5D5VUwoUHZuKFmN6aqxiYHK6mpsVhht/Fio9aK7z/1HXaK
Rbqa90Db9+e7StIr1Q3Bd8K4Y8ULPoxE1j/Jtziy5UE8zmqCMBt2W9GFFzN/PHAss+Geqa6ed6j/
VcZpUIeC6s4SC2Bo+52uWgAwXIlIidSkVWSinoRMDOgmyjWM807JyzV1V6M2yIIDmiFvO2STiGPN
ilpyibqh+LzqrSscob6NnjrlvnybTLLUF6YRNYYWsw0jPfj0T4F0TkM2Nr5p3KHAswsx0M5MOLzS
VKVEUE7n17tIW4ew5VVx+SgQxSjsFrwHDJqKPyKzUKVuZTj6vfUZLBuOXHH5ToTQSjRjrYuvahEu
Xif58FFZcU+0a7+Ag1Lk4XkZpAjpe8vv9VfEIcjm/19nYj3imqYVud+78Uss/en7nKMSrpWnGbdR
kXceMicC92BD3dxw5hlcVNN5nzjdn4SD/Nci/viltxBeXfTxR7oB9Y4Fwbg4efUGP/dQv04o3L7Q
2HF+yoZnMBtH7HHWn0IUBUKpcrqZY1t+1eN12HHjE2Leo6AsWVXcJpl6LcMeaQ48DFG1qXeAcY4O
s8aBDexRnwD6v48rU11z141MzvsZV+5X/IDF/myZFiig9HNToYY1bcjNpOGuLQ9/f9YvxjpvRnLP
PJSRHGnRRMlLS4HmiE0zIhG2iJeouqXDgMBd3wPUK9YFHGLBxwBR9yVEfK2kOqQg7xVq+0ledZCN
8RTDEFm0RMMpZNvp6OwzixYAHXlC4qfj2pFYWrTRpJai5bw82mc8McmyrYq/K4DxYxvzJOcwS2Ro
+Z+N6qnfE1XU5LqDT0jmv0I0FCXXPdcw/rByK9e+I1odpol8hs1wqVp+v1lWA7P/BNTSTiAYkPK+
p3KmKZ331tw7ahDQB20tFiTp7PSFwOCPqduXTsHUzbrkwMBCh6kh7Qy0399MdTy+TdAlat2pTE/3
WHa9ukIzP3ISUTZfPtjbpfs4aVEq9CSlyNXqseTFm5eQ2/xBTQpjZRaNLj1yOgeB86F8AQZVaVCq
cnGaLBPkeoW/34/qq+Cj1txYHw0juj42Dz4vagovF/PeBiWhcwbELaqaDys+rxRefIKF2FBkuQ+W
URh2PCnkbhaBJDjigL0E5sr1BhrZKXKUF5vBoWTPdv1jYslTOyNC1cpY4ogYerjOrLvMsvZwzVkP
vfAGgpBJX3ofN9pay5cwjRRI04KWx1CFmPwVCmM0lN0MVNi4ojxUsOJGfqj5KN/yvoNz79Wd24P1
C4UDxf1IAEYDGiKCqmDpOpjVsKDlKgNnml1s2llY1ijukXvjQewrXaFmtOMbPFC6ZQGmFd10gEJD
S8llpe8qlTuONsFirRJLFDkMHTmylF59S5UUtbtRUr68+rDhBoQr3suheD/YgSu2snb4PUYf8bW8
q3VsT6buqBpIZW3kF2E6B2E5u+WELpjEJPEnx7QOy3YODoiC+FVvjP91C95SPHs0gCDwKyJDR0uV
vVxvwvLfsRAUUbH1/nHa4kE0L14FlMHIbKdBurImdHWuiw6pO987kbvtBJGjb+u6neg2AVCJ/tl6
/gmbxZeWer+tQ77/0IuNsb3C7vVjai3OeS5WoMqxWV6TmuEE+n366Z5fzdOtjAqVw3xDUH+B9R3q
Pm6l1dOmvQlNKakt+cWaIUSNcFkuhpl95yjL34H+XU0Se6hamQJK9kaZZXykVC1mFjDs/APNbMjB
s2CNNMr7E8w0kXVqcSbOFM5lOWsX7FfgIhzEePsXDl7nqgY196923XyW787Z7VUezG/8riG2tT5n
aUZdDNBtOa04fF3LFA8nG/ceQLk30EvYu41111TXt/47cWe7fs7rwjUjGUJxOk+EIQl3fvQGimYT
OP6aF3kiRU0w00cg61ICe2TLwW72xLh4vzhXL0mFwE0Dvj4Lppi2VvkggO/ZiBFkClX71QfZNAFy
3CDRJgDHLGldX2HnY7SAeMhUqHIlrUEhzs2eaCAEmdGuKqiopezk5IixpG5x5ACpOMq9I0H8PAAa
98YfYHwwmW5x6CKTZpExhjXeqF59pHH15/8RNiueYbVNszUzQfSyic86zuWSzRYm3ouXyM6SPe19
5C//crpPcaYVAHtP+KAw14x39tzVD/ikZEsF2Fw7h2xrsPcW9+E5BrWSwe8YHNTlgZXChidgDOrL
dgp4eJhzAU7Tzn79Df11bOs0buR4W5lJwtstRP2EV15M/g/clRuiMGbFKRix7JUdnbTAg8lGPorT
bXvm4hT3hMDBWwiqh/GfuIglR8BJn7nYIcBVdFL/LELAp8QQqMNMWtt7WAVbotaJww0GEY6R6kCb
/coVQ3FKLp0uy6VJ8OwzgL6v4Lu9Xj9JVUyiiQZB4N9/iY0aTyT6nOefZqD7FTLL4hydTGAcN04e
T9XFP0lviuebhqSNudCDzTnVnAK04PnKDFp6469NMudZCM14H3tKnwPnFZ9yvWAC6FznWIx1LL1S
h/YESRTB1WBYorT9H6Y0IuJd23LJ8SsjQXWqNsFUqCr5m2eK1IfC6NAgnC1DAB4Q5z3dzYrlypZ/
zlSvSfaQycwXWwNiwNPcVu3eux1L1dqfCMTsHR15HzQzwCDtralNKiDm+6EAfFsgp1twipL6m2J+
Q+QFt8j7R0r6xFALZyMpd7nVkvorgUcr8iJZcEgWPxyUZMTpw+4L0feMO3HIQqnk3tVnS4UvYf+y
CBNJzwDwTRdMGy36/CIanBAY1FCwCSJTJsM6VNZtOH/BWAwj2ZulIwwi0lMaReSDukNnhiRT2o2o
yWgJggh64bS9FSKfsfj8EaBYENbZ4t1geR1FYwCvpVEeGtT43c/T7t1bSaiZAgm+2VIef6TAHLb8
sc0nUYm5i4uNwe0fc8pgrMh2k4nA8gqcXFRu/GpL7/hRSYAwaYonyOFF9493Iy7a1slDXWqCQEQg
UFaf8zBzX7gaeSeetRMaGaj43pCkMeUl1cPe8VsDsnx14l09HlWxTAUQJMYX9BrokIa74x04/bXd
zSOxNXYvmmzFZKktuWCr4QZ7s48jfNvTJl/qg4o48mABN5KjNY1TaHq4oxCMDhtyvZ+OtMmb1Ur6
5D335vq95pLquuOs06mbGt208X+Hy6JDxqhmafohYF9wDdio/GAbu+FtDKHgBePHWVk4pMJv6w88
fWTKF0FOc1G7lTx5w8XoJW+L4rKTZ1aPRmwMHec693JyBoCqeDSPJkUTFLERvXpg3Mu4GMdsWyU0
WcB5QxE8FMt/hFRyLXjHO1YjlvNadi+ys80hv8maLMqJ95Nv5bmmfOkLfr9sH0hb+mo7j745Cefk
q4hpmlVnyJTNBmgI6bw2XkDgKc8uPpSm83HHEDbnwlrt5obdhajBV7qNwXVxSDTdkJ8eP4K51KHm
zGJxkMxBjO6WppRGJY3/d1bd8oV5cRHv3xUwlJ8yWiBMYQYfkrQI0P4p9c50AbQNB0MkhNsCvO8m
m3slbiFJC+ZkiB/fhbQ0jT8NS1GoCoZ6uohUpQTDMwsN9iKy/3AcBKEk5kGYwa7l5DzowiOGMhWM
bE6HWWkN8ScTSK6bladKHCeLsAGErsug8G3qcPbxi7WY32PjvFJ87OPfk/ThBJqs8DM3s21NI0U3
DfMVQg5Hs0ylUJccN1Ozb/IyVVDXlV9TQvVgxs20m7cQjE/2tEvpeunEfYiWiCXB+bX4rtr3P92x
KY27MeYkY5ynOShVrqceNXUTpAS/Ogoskiv2i4lDvjjKMRkL/S/AA8UF16y//v/owphPrhVNHX8M
MINPm38E2ZkjkMumgdiugYYMgvRPT9DYLlijEd2IA8UDVn9GyCaCS6VUTVWvKsrkwlwqtVbcI3+D
rb3XS4RPojaADRXxhyLE+GakZDyhN2bXoZyFNwvJKqeKsi7w1Td04N1xphpjl+NPTn9VCOOH8WzE
eTGqUN7hF684ITRPZauKs6pEP3u2c9KlMaAj2V2iqxxiIngLv94B9a/ASyiEPvv08IkKyGAL6VLb
UXxQTMSeeNyFE63OEsQ1APZv/0eNdskdG4gnz+Nph6ti+GZzCJ/Z5olf+mT7B/7pWqw/F8Lz01Sw
Y6Y8rNrRBlKresobZVPHyPS4nLCuy27fjEOGd3zI+qjE+4m7qximk3MIcPwYgeQwPpgBC9mahpPD
y37BEwWOgH2pGiQTlaAj3zSxQjLVlFCS+I37qcoIYMevOWXQr8xbdskVmTOEw7PwCPjB+sLRWNLO
4RBHgeqhi+4arITowlYmDK2YnaN5ikjVZ9cdIDWwDtuemuDDQ+tC04OAH4wRIul5OB3e24QvxZtW
TPrL3pqNyuivSjXW44zPuKBZOnhZpmSK6vy4ebiAQIROXbt6bMEzxRNL0k4nme3H0ztv39Ml2yq8
/wlJ4NAV2IlHv1JVvD8xAlhPRf9wZlPbB/yy9A1BCcAx9SXaoEcHkNIE3yGOlfjVqg3DM+HaGeB0
iyo3Fwv2vVbx94e9vp6snUaQ10EfdnUTwFVO/1rf0vWo9xIebfmrsv5NAhMoyz9pvegrQDHOs+T0
R41J3UhJvcfsoB0HlnFIGfHaFPlh25UJMFCMJhiMMPjP2VaeUJ8HY1PsTfyrRIJ83kVRTZI0EEkL
cGg5E06gRgnuOHRafbERDS6VWCkwbEt6zCu5+p6ZTHoWjzEFVKjI6adj1KkjK/mV/V/o4Aup873C
uzNn7u+wOsmSVg3GRahAwGpJBpxRFtjpLCVLq1jfOhItM1s7nj2T5XtyhmqR//DLCPpP6rxfEy88
viNGcjllZr+HMhsqI/jLW35tNQcoD6+nF3WBNzijqGOVhp08TwBmyeJRG29fGyFQhShhEppplna4
1NBRQxh1KabK5qpPqW4CIZLsowyqKM7o/TChFDNcQSvUXCERe6ABc285rW1IpRDNvBysoMb/16oZ
TveRqJ0iR9s61pJyAQfGwVs5AQruy3i/NaENy9qypb8XoT+fDWfTNAepVEATV5mZNwbSeL4h57X8
ykd6TXjxrljsPoU/+ze+MUAIa881oOzFvTEl3FYsNs71rsi/zt95COZ/e6Bz0DYIBQnXdRbpAAwz
1fmwhRCUOztYR5ATIHFF32tFMhv4jFr1tAjmb1piMoDOSM7YwTh1BVylTZMj55l1ykC7eEvu5r+h
sJ4+Q78WtITttCMQvZXkVb5vH0R4Z10cycZy75q6JHw6eNM6Jzhbzj0cBvi8JqWIBnuDsRlC0QZ2
aOFim/ItUpGbaDEgKdysRZDpxNHkWAK4pdZRatQgYWl44OJ0oTAciXZaPWu1TQo5egmFCix2Gn5w
cv//CxjlaFLrP1gtM1dLD3hrp14iB1xehTM7W7ld/RYk6455oNsqBDywTO5sNva2V2KPV+aHR0W5
qz/Z81tN19ynczc13pO5MrQnb+wzFyag0aD0f1NpzRoWJwZPHUH8iB/Sl8Qxuu+TzW6AJuPsHbjR
RKnldpITlMaCs+TCpqbWaEtjmCF29APJstNXGg/XwsQknRk3C86DIjIITys1iWW9bGwZNj72knbP
vKih8+tbwy7+sKuwg1pi0MaGPCB+OQDbhCmuEEkssMuYYBbpCXMoUL1FgnJaeOjHoFxlwW7dbLj1
T63OKA6tas6abb9YXe3GVdKZgXp0tw5ItORH/4ugzDDsZtQMYv9PPyfnGvZdPmKH+l6Qtlm7+NHl
9AdYScWjwZIdRe/tHhEenlBdUUtKQceJ8MBnbm8XLU7Bihz7CLr7+aeuj+klG/bn9PQ6HMpnP3MK
+SHdPiKQtBefdrVgvJPV04c47+NmngOwK1goB436oOwb2TET+efsA2+WWkocuABUurQk32Gh7lmz
uZc231K0EVVm9MPgqLoIO7VYYYPw+Yb4IU366Pbz6XX2g5cF04Xj0FHzFLxKS52mKJ0s+Vhu/a0P
UcpRTRqQ5dUIMVRDUBJ6hWNKjXxl0ZEBGCauNmPixJ7tu2TzQA6grkZUMwiI7+H9JZ9L5K7wVZXs
1SCQwR67OA5nuhUlDxlbd5JAC/UouuxVD1nAURMzzfzeX6NeYUrEVHq+8ptF7fvh8G+K+VvqZBsu
qUHL1TNPYXyRtJS/Wq0oAfCA4Tmbk+rNXqgUOJSCuMxhd4O1MGIkOA7gNl0yfptb37xsjm6rOBQq
RvyKfDbXv69syuHB0HnPvqVUeCcIYTa/S6rykQyZnYaogX8cLfKPV51KMgzQL1Yd6oCGEsKKEc9t
MlM85uLV7r3DROqsSjAnhfQjnTSCds7GZisoVdqIC2vvo3igWsyJAFno8Ocnuc9D8qHD1yyuI5Ai
Yto9d6wwlSbDpmN0U5p0PeBiaNjT1DhFoj877knvrV2H8Qv6fBeNBiFbxGLfLPhl2gzj3CGeOG+r
NvcRI2RoM/GvebfyCacHw9zWobHmHOAg1HaZ9r/Evsx+oNkWA1/mQaG2MIVfEGiHtsIbGKJsRWnf
+/yXKpWea1QiK5zUfTMLbowWt8vGCYrhAQpmoDZEsy+BafwvmLffmiH+mGk50qCxZ0uE0W3Unr22
uwaCzBOfq+8c5a8C/MoR3MZYjqMXA+40mAV68d0HLgpSJiO1Pj3yqdbjLGN4X15hNdl9sPYao6Xi
uMna2qNwZRmzgJyO30CVeT6cORvPcRgCG40sjLgUPOCRDhykeUr2coXxxK8kebwtZSm3UBKqZ0yg
QO3Lx2Y9EvTHOvtQkV+7ZmI1bL36V6e7pCoroq9qjK2RmM0wq78syjK/YEl54+F3+M9ZDsAQjJFy
4j2xQlUW7U8zv3QLC0J0gWdyrV7uj6rVipHOwZZS/GDk2SS+nGISSgCymKfasWNKnumlm5PpGRp9
Pyt8LEhhtndcp0ABWxhG681eJSDROtmKJewzjVoZDbLGGHAMEFCNkuxSC2fLoCafMxSuobygVy8X
dfRIH+/hyiargGmt6gscpq4jloqrIVzooAt2/RTPjCqZplyEfCBsrdsxxNK54NfpokL8cZslr/aJ
0d/yqsDi2e2vCwBzkyuYSKA5j3AJoWgryBV0wtImzSbl9KQanrAmfg0Lnojd3zLDKcJVoQn5piPM
h1KYJCXhdthWaQhj3xteyZ4yCfuhxSrWWpNJgh8m1DSVvbzExjUB4VBXVOGblqPnRTZIC/cXM2hx
bM0yWUrePYYG4krtBt/u840JsgGqpswNG0nNlyEja2Bkhpu3o9Z8kO2273D3qTb+h5cFhfPl3eE1
HFTzBbF+Lxim91kgccenxA7+Hc2TmwqgWnXVLR4FSDS9nam48TzVWPsCTxsXRIqZh2i7SWXFNaoB
lQarRYewqHbmt0WMDHt0yCn+/LQ51rm8eR8XzDmk1vsELoeRvHMDGr1yrGVRI/SpuUrkNH3AzR/U
KoRJ9AVbLLG6KlGLNk1OhwhM7i7zzf3/iRrmrNP/W/xWWtCPPg9OKzqyMmaActbKyc8n+Lk2FJ+k
tMPmcyRFcc7h6NrsgZHbbMFCFMh6Kx/GSHvUmlCZSNKHyZ3i8A6Bcwq9dQUOTFvLCstXa1ClYxzy
nJ+XDBYHMOnejMZtl4Petzvtis4N4NXUDMv0xCSoik2B19x4PkN/7/oo1Uvwv6IztVK4Yi09KSXj
W+UM7iQUGNrmSL9Q0YLCu9gpK6o45JiIM4lgRlYdaLhg3fvhRm7+TEIbwKbGY8+5hz9PQzvFmpBr
NWuPClRaodc6c0Jan3W6hMTq+7G9PEVL/nrZbSysE8J7ksC3FAayRdwwL4RT9xrzZqtGOKzZEzQ/
FU6F+Z+q5tMCrWWys2/MEQz1ooGYUNtpYuWWk2k0ChFExdhiHZXN4eDcdRATobMRCAvQ660AsUzn
5oCxp1+2pp9lYnL5AqFqXg/6oOqDgDcKEVLBSv196Br3yztZY/XySMvagc+2dnM6Q4kb9cZQ3ErN
5y1HzDyQ4xWv6asL09HBFwLJD9yBXrr/cPNVOjhKwobgvRvfip44o0R6HrK4NBR6hEfNHbDimOCi
lWdAwL7icRtWo8udzNcOviCb4YQm6aY7rfLmXaEyYf9AFu122xekqA0P45O8bmW46nwcwYETuOdJ
FGLECX8WkqI/29uOgwiBWAtbnNBOF/1zmravPmJ4UN4xPsiwcKYKQWOglpz3ppKW6oPHhDqkLhsr
bCixctGN4xw+VjkJiwoUIdUjKvwqgt1AWjhkVPpqfIFAS+wkDVfkzfs67Ts0YXF7YFof02ryekp4
1ecTRdFn73ij1sf0/c43rVwBHuy5SMkq4cWAoT5Hgcyseb53PYf/ecF0HbBOXx7ioBHTRoMTXZee
h/31qYWBIOjTsssdnyVPDvwka1gPYJYLchFPOqVpah2eCt/pLFA3YMlk3jdTXyFq9HDEpmkgZHNt
K4X1ZsmxHZQjByT5U1zibtUiTwbkf+AEBHKuiaZA9tMizsBxD05OIHW+V9NAcn+hqJCpSuwaNvDS
ZXwVc56Qw38gpOUa52NIZpHqOvH0eH8yl2JaFb2Vrq2zOL3hZ0PayWW3XBH8/v+AHMVmDLG3ERux
fIdR3/enlDtRnglRVWo2nLK83yLcvsyom6cxBILEOdx+FE/dvqFwZOjz/0FXlEeZxTsh3dkaJiil
a+Z8aBxJikqVHfsOq5hyZDq5bRH0Vyn8zjSikLb4NGUJON1kQhE2b0BLBDriQwAbPIIwY4dJz7+n
NUrBZ46JP98jr9oVA8EjBWPoAZ0ztABNOw0DFglIwENJzsBuCv0mBMy6LBhwJHjX5urG2m1iDVYX
yJVbQjzj8IyOgXaOjpKYlmibsWRWIX5mWl/31e1TnjKROpYhbCArJmfrhnu0Ij0aSnYaEwULp3dJ
rrU96q6Jukymh5gMfNP39iYmVAIlk/hE/VvTomXIZ6DC8zYIqjlN2PQe8KANtp44HJpm4zfdi5ty
Z5RXzePWz5ixVKuEgYcClurjVSZas3CEzaIRYtT8oil2WvPMVUEeBi+68nF6buTVlL8ZalsuQsT5
CpEryhPc+2DWzscPBjClUEYqCXq7Rl3mIk4ClcV5jn+MECB2UZW57kYYwv+8xX7j/fHwIHx262Wh
FzQa/E5Ag18l6BR1K1b1SCF3sZCSLuEWX1pxXTy+5KrVgLH+C8tYBsd1Ob1DHs3xI+MEGF0eC/k1
PmU1MP03/HbAhKX5fIp9KGWrgpRslX9WnQ/HIW8ufA2HVpoTN5QXecp50g57u5kUP+qD+8/6X1Gi
IFS9Q9w7dR0ymeH1aOpuvVWxMJi2t9b9yExjIEqy2rDazGzrZ3EAu5eAKYbWueKiPQmEuUwYP1+9
+BLoHuN7ZWGT/Dr7jH5QmF0nvXU4ztAvedLkWHrOnF78VkF+15o3/dFejpyTUb5qVZcMapi21Zyn
X+CuOzKgDXXIaQm/PafYvkwxfo8L7nNOmKmtCrPXSGRKNwsy5M0rjuZVH1gyuqP+Tae/e9zVO+gv
M4ZLSLSnEVtfcMZMCk/a+bi5P0f6xw+quG7C0lyw+BEbI/ls/UmDk3uNoyN4x1tZffxN21uxaJyh
nhU2xGo6sfhzQ5uSxcrd8yDREi5QbDJDcmxUcxXXNDmMfdxErBRl73WjZRZg++r5IqaHNqfWlFkg
sQAwfecIuF2XTYIcHkKvoCA7u9Fjd7RvyUc0dQzuGPfDmoKoymiRcJ6Di1NlYIZvnyD52qhNUDPQ
P2mj8crVY026PSr0Brs+77vNPurw3ZI4Dymo7oDAJdZjHplcVarl12dCHPrX7eyh4td9QjjQoduS
oDoTb6E345MhOwBFLkvW0JYIoAhiOcVm0PssB2gCAscRXTD74g4UErYyKh6da6wm2eAVM09Ibjv2
ISX9n2/EOBJ3CtLKIqRZ99h9qtWWNJJ2Ncail6Zra8RpcJyubgYNCMsrq4qXksAiczYCrWm1ZNz7
cEL/CQvDk/1QxemUiDdM0db9PBc1/EdSycXVJVLINiNc/wuoJDMFvvTLQg6pAaHxa92YhbrREpht
YtmOQBMcvRVj6wr5/kyy9eLKqXBvr3yK8MP9e9ocU4RtzzGIwy0LYaGyHCn8VOBjkLsC0eYCyJku
q+C51iqdeAB5af35M5ZjWZ1bH2dXx0LvUkFq9I2Wx+qeblANUUmNaUqk4P3oWeNeEcW/XzTYRrs5
ORQ54v0r6JVJiBgXx9drryNnVkGPCH230mt8Anqrs8d0NzU8m0x0JqIc0TEgsqJU5fFkDrKZs6M7
ZiX/mIWknJjnj9OW7gbzOIWTxC+f7LWJfBe8PX7qYu+dYYLTwsEcocsUBwlUxUw7AcTcvn0evLkq
Z0AtSkUD2LjPmXPEjqgjq3NB7zBXy5lV9dBGm1jZthyQfGHZBuc6IGvlkN06KCLy8xTkaMwa2XdA
HEdB3SvUfx5fNLPvhnPBc4iOagpTf0okuFLcE9GbqCTWW4JgSPB9f/ZETSSrFy2s3TnG2sU5Yk2y
FC+SZxFYXD9UIcURmqW6kIm5WJ/Wifcxk+BPADN98Vcan4C59ItLWlBWtjiNzAo7YJlkUxYAXbCs
L920X1jR8TXrrbaI5NMolBquaTMdoYGWkRYmajO+sCY7+qtaW+/ASf1TpycGY22y+Frwe8v3SSKE
xgLQSSmbXhlQIa2eJTQ4xxGbDXx8RuKF3YPdJ+KgCqCiN/O1Ylh8tw7PBy8f7eElnRs6aOZT/jCW
zQp177W8jXJI4G0dktXsqb8fcOgL4DzdW1XwylEMJqCMxS0jp6T9fqH3P88eOUiTlkBhbHvbCLGo
mOSD2OrnxSKybsHIYQL4Hb84eXLZvJaCFRt87ADJVRnssBN3X6vUaCEGpks2PeeFywL/Ns8TXxze
+lz1diokXfbIRO2ouQyz3UDKGig1d6Z6g1P/gECJNRHPz7oqkbEC/3zWmZ/3ZrXX7VfyBIJkhESI
0u7RPs8Xtr5w2CiXGcPuwtL+VB8GrDEGb9SrfwlKuE79EJcHrzV9tY7tD9wmrEJ/xe2/3hd6s8wD
2NePPnAWdo8B5p4nfUmkCjmPMydizVYA6U6Bki2ecyxQijuQq3cbid71KOtkJbDjjNzVenBO1BlO
PU3Wh/4jyKFdOYJOQjN1GROtAp9ujfM+544MwnEIwav92oK53Q756nHKXmkz8Xcixg1mvEfwYZSW
Mv+dd3nK8tNWvCtHvk4mLipHog4IPtD4EEydxAW1/DqHal6DH2Ro+DZnVBg9rGnYEqKPVNamW9PC
uKvM1DBkwbLpwonglE5tz0MczJmnsyU3NhqeKf0ct137ScEWTVynlyuAEP0yagZdckd7ikwJ++54
e7QyExbqVrLPh7DLG+C/haCM37bAN9YCKuhm7ZhLp9uRrDdWTs2qiObpHHVwAPdIFj9Kge7EIKpx
u+xnEDqJNOI1adh3XrxXpEmJyeK+14htDxK6oBrlq3la16QWD8lEPYDl7Jp0HWiKkcD8W925SRG7
OWoBxLFAqrGNQHvM5JHQl/e4Sqk9SKEyra57JA9F4hkGjjxF4Z+Q/5Dno9Uuou6Ky/90OQZwBO+X
DhMnY+0Xqi6RYOUKQrIphja0JBcxYfwQYqghfZPLFSRltASkjv6RKgI4XRQAHes1qZaIPo7USda1
MmNLXWzgpMbeAoet87ZcCDhlq0OJkFXHLV+Npy6yuHBPgT+3Z6SCGgk9my5BnYxzA3STDQOZfhE5
QHET8gEUlcX2Unt5UjTL+vCvnX+/k8/9EPo5vU3+mAgefEvTtY7g9g6Y3pAZrncbYMX17mTIdwZl
QqE5zSWu2xiEwzK4r1GPCvX3/M+i/tZNb4DrLzZ+vCqiR12/62bbVEvEWIiaQOEV/SvQvmT+h5yE
2WHYvYTh33n8zEfhGFN5Rz8sy8sJQSrKekQod+nHbqs8yvmZ8sVc+R6wH0v7pjap0R9A8tMAxNo/
o6Tys0DmRg/UoEmBZGzfCOb/NtpeNLaAw27DVZ3slBa0P6ti/AsgHBsU7uKZ78JsdivMkVnDSDmB
73zExqS7NWmolMUO8jFBqC2Bu6WM5U18l7HVM7YPwScfm90f2+hpARx+MMIfyUsGP2CAqVXgoMmN
zWJhQ7fBM+K/3ymz46OhFosTCWMHcY5XkOslRbx75dwYp8Rwn7lk30kkf+xHbgC9K4Xfw38s1EZB
NbUsURecT7pMObf1dZJ91aL/13/hplZVsbtTZSKL3POAYOWayJ2lAWoUN0farC4w4GDJ9REtbfw/
bgqIftER+V8D1EIYZAND7ZKCtIY2GpIKdb8LyxeusRVxjf9QB0Wd3/0I5SR6af9x+xG4rx+SW4qw
69yxeSKGDUyR8KLlxpH7oWO0XRocd3RWB+V8EnooDdE7B5gmmaxuHuCd0fqCJAJNuzIxrt9kk1bS
aHwPr64zJVKYwWIzAYqiAb4ViRK4vjehyQwf4Hnn/ymU2MSmSgV+qCfxAC0qB9cP4AKY/ctxNjbc
eXQ3Qr1mcHYqRyQU3qODDf7+w23gD2gJVJY1gIkv/m3lv2QQoNXXeh7DDer/G4cMumvlFal1SKn/
6625pnI7DqjfjRd7gUTxBuBCY1EFn4ov61UbKy5EcHFWLGy5Ccyzt2ndQ9HRG0j7EH/WoZEokYgP
RI3AcuQnc4RZ0w1O1YlFnPT6UocU0+XA9/gUyo1GPbDxKX/Glai7zfd+VPN438PJPREvUgQiGkkG
knwXm/Ol0ZbvhTnGrSvLvbtm22zqa2Wqz5lzlHAs8KimcvzMrpUHLFSVV/5gFDggrdxUPYfCbILR
Wc7/MpAyh5x96h6vdHKC3eI8AqRRqb63/h/lDN9yW/xTUkVRFIlhY9ANUPZnUn1Cmn4uhiAsLeHT
aitL0BUWbI4lAEy9ef5I94f6Kq/AYcwMvl28PTxtVNsgrHZUdqs1dUo80EeDJsZIbb9BUU1SFq6j
2pqvlA4wy1u1K7cz2EyVUfeCBbNO8C7Bty6cPSO4CkiILr1BEAdB09PVAOOYZLqpXrdmTOm8KszG
SHsInR+YvZ34qQcNt6oyI0dp6tMmIxXBKxySBhk3CX6I4sRUNFRm3FnSMI7BuW9PntkoOY7CkeCM
kOWlV4WV6RPcF9pKq/njbFKjU5+b02EYD+v+cu6vPlspRnVxc/n39GgjZ+v0DkULX+28NfoYfiPm
fEoewNO6viCnotF1fK2mCzpkDnrOKjmESpmfJWDn4TtQkTUpaif6eSl8Qqxh8y0XiS7hg6s2L72/
vGjRQruUsKWrG8zMuxQd4a4G9WhdM5Jor9g4JeaJ9gN+mOcZO3HVhKI2J0H2d1xRPYXOFSpQv5QX
AJpvKE6J4/iXoBMVzDvLZUa7E2V5KdlKwt+upG3wTwlzD5TlMoz1tyNgJ7NJhVYL4iYPnCTwqnPy
wo1gzHXr+SsFcaiYupO9FfchdcuC8IMCcA+HdGIOc8xl0hjO7ICyUD9ijj7n5ntGZw3Tj+toBoUP
xk4/lqpRkRma5csclavBZgHKfYEkrhaAUmf13l+fmSbPnvWrRSVjB1YLIwnMaMB70cUuBkHbbwkM
TWsqFQIRU/y7F7PNLDsGkkWE55cxjhTDqMYG4Gaxsh7eVANlSy3wJn/IB1ZGJlxPqqgHJlzpUyFX
xYFMRfGIvuWwJ8is3ivYeh9X81R3raago7YTa5jv4+cJ2PyQbHpJt1f0MBv0dIEsEGwD8WAiMBPz
N9EkuVJM2QtfTbzl1myH8rtVKkiIE05PvEGY73vlAJTfUBs+NWZ+vXCAw1LgBwQgUFo/bS/afFjB
juMKA+7fE5+yU24D1CqefyrjgJthQYbs+qqtz49lzrtlcz9NMDkCZHV38pbISpj61iQcmXlRqeiL
bFNJnGhaRVsrD0QHGn8F2Zz/maX/4ei8GRpPxurDubhbzhECpGRBx4REmWko/mgoG/f9k//yUP+J
ClBLn3rwyGmqqe7CmWt2tdetm6DR6vooMSQqReB2xVmGqjpc+ExUZB1XzE/AkxXLqBnGgiHIguAW
JQLm1eIqYxJkhMBYcZ6bZR5w7mHWIv+RsUNqsc1UEvSWeeRugdKuGe1x4FtWkR/GJbB/dU09rjOc
PKrI6IngAlkzsnXVsIL7Gf5KcjYvu+8mUR2BFwrXkRJVBvDwf1xqASJcMUa/2Z77CqzfmUHpVd6D
nHUBj4ksvGrRVqPiWMH16XJ2m43fHKU/GN2L7OxB6t9bpQ4ZGznCj+DU6wk23uU6LLvvMXwk6Nqs
RaFSi7vX6so9/CNu3wtWfL+lp9WifuWB0VGCrKO5Y5QYz/OY3ZCRmVqqjD4dh9ScQCtZEge0GtFO
tN69ASU7IbMlNsI3/7EIaRduXWD0VsE9SxjOSomsI5XinmRqAEys4pPxVHVfiRWSb5MMJuvIyWlm
hKhVQznKUj9Ji45aj1uoA3p70zN/wq/mdXea1uuyE0/23slP6l8UncuVwrCBluOC/Ez9JqU1vieA
XMpYH0Gy92fz/kZv8lDOrBqxss6SMq4gy3ARvTWF8FMuH3HVJziV9r/FzwJjVI2YgTi4/Vivcg9Q
jAlNqlloIDUIGdHd6yt41MiN1tUcUUohGI7kGegec07M6FS6fYYSY0Ui+rwvDPovxP1xl4/j6+wa
je884FbSSDDYX3bUFTDdLH9e7Zkn7bQvgV2JbJ+jQ759miLLyC1A8+j277iQ40S3BOPuQEEcJ+L3
ghLuO/iyr9k26Xl+fbL5dd4vs72b5xbqmmW1DzvCcX6LepLzqYX1dR77SgMlOBFdbSJqRDor8qKd
3mdOJ5bN0fuLY5QHo6T+RWoZ7QRy6U7QEisZVP8PfXgkTcn86Mz7nn7zg9yAftIOl4f2XiB19TIP
y+cpmzkWUh+Cv78tKK1ZdC8TEHMUXVwUFm29L1uO5QFF4p2wsk1wEzf8MEMMjSp2vFqGcuglNhA2
C1J1c5/yIP/+nTHzOJEuFqKLRVBoHDTS9WFYmA5oqGmDQ6TLc/8+6uMtrW/7uDhzJ9Gb+1Z/itUN
ZYunDf5ph+rt3+q8Mk128Jd8Zy337z3dhdszP06v6pmv2qfrS9A5ZysF36z5+86dz6u2ZzUITeNF
W7Tq8YpoEwp8q1jZgcN2xcGmTnL1I850Ju0yB4UPvjqbAZd82tH88WhDrpRd0C+gGCJGr/Q6gn3t
bN1wqD6iq+1rLSWdOdMTFIi9EzqmHkhokDHwZXGTuHdeqiDbFp043Qc+ieywAMc+pdIaJkUG3nXw
0WkLTtdwDmWiYRcU/DOUnZfMbi2TAdLKN1g1S0Tt0FEia5Q4jtkbYyQI6LY9HXGFK2GEv8x5tCNo
hNOaAD0XnVChpy4xLhvs1Ajavpuz9I587FjJMnRSlO5gTjbMMbOxBzpLnD+KBQPi7vWWGcpT2VVw
P2DLeiBxO+q4hhg1Y/CIyLIcoqZhjI58FPBVWHe7vfdzsa+SYLR37kbNdtoTVGvItu877bcHr2L4
gGaF+j0ZaYFWFGOhgwdn4BioYCM+nd69efvilunHTtK2d+ohq2wdTxNJS6Xscx1ABmhYiHNg02Dd
P7k2W1/GPZtl+somW0m1n73mxflAjeKni0GKOLwFx+ikLk0uSqpo37Ssyk022eCUZp1lTxdTu7GO
90z9G7rJd8G91eryVDnp8bTbtNmBFZ7YHpycY25Sb6LEGF9Lc5DU5SXbOn8crgmFflzC8lGwz8Zs
QSBu15lZy/hiDWp7uQjzUsMPSPWavYWTYrZ0Egk+/55S7zEdT65jRNlgPWReTO1cmnBW7qz9v/xT
UqKRWuC1MHQsnbql0TvZat69ED8pA2mOE/96n63hJwr2hw3y0i0gmcuw2gcDw2JfrJnIOPP4ijV8
560f8s4SSrMEvrEWMCCs3/NxlUYbzAOHylKRYmhMKqi3ooeL4zNdD5sVx5gUJkjXHwF6M50wsLku
CjTpL+S27xXeIXOnHsucKDrgOUsO1iEhtKjw2EW55oqnsjUUwi7MXka1MUtmS1oLNzx210Bkjcxq
Pm6XdUCU9saBng4oQMnUUmaM6gx0UBaBZokQ8iMDmO5v0FNhzwixZR3oESS+ytdEs6isUEcyoieJ
wnHErdbBOSSlIUEiCQmoqp89scL5Dqeh3+Kk/aELrLDl6WcfSrLqDG7f4g7/FxiB2U/3rrJBtV6t
D97ijma21Viw/2q6ePmRnlxZWmVN+C5fyuO/ZHEVUnI6Lf6VA6i4uEKLkTJnmmpK1Jh/qIk48Qn7
h+N4aKfnwiF1XQ6gTLodWHUvnk/EuwYEgyIlUqCf/AoFjsh87OrjLFP7L3+8TsevJFEbrjRZmymJ
KOKGhLvxgTYssTtE8iHlNU/y3BFXVnXGobQ3HG0FhfRk92KFUmNywuyU1s6YvUpdA+wojXR5ND93
cVvCVH1CEktJmQ2EcJqo5RuZKnjADjKHKg2fDqSLk9Bfi3IrnEpRAv8aIusuUzRxq54QC4XKPZfV
7U6DMDjVMhmUMWbbdJTi6ckkLIvpNGNKDTOWyuLL/lVMAOayTDpi2kKOnAXDPOeZNSpsAcyVf4DW
c8d1/ocEmz7C60k7aTsTKvrLmURmsLEarf0Jy6mTDCxXV3oPaLevZVjLNjS4sNPrhWhb7jPcqX8q
TSNYTjYORbHZHFnqLsA1DI58It3xQCO775a0hXEanqB2W/hh7WfwBAu5igDfhDt4Xh4Jeghu4p7e
prgaGAvaGLY30lqtUZjnwjIhI1NHLs1UiU5HNCiz8GQev/Usf5rkKwJ2bguDCU2CboBqYoRU/gGI
YFEw+xddC2zx88oX4GtlOXJat289TqGRSQODqkHcBsWBc93V+QwCv4vlzfb9TRQg9yw8HGFspBZ4
bBRjnwNvuGbk8XAcoB8/rz7rgYtE13wSicybKRhdWL3/KfNxCrRqa7z/O/JiOpd/wYLtiOQ8LNfB
rR0+PQRVeTzKlnxmrwCTYVx1DOjCK7d9b6Ei8xSHZkmOpFIxrHuzvF+g7i5RmRUNoKW7mZZfqvxo
IqqPuusMl4NGdo1ewldKdou+l9/Vns1jc8wasHJg4BHHdwOkFxHobxLnOsHWdLLFqo5nDVvCqBXz
aLw0OcapRuFefohnK8/POASAvQWq6uspRg0kDE3IEO+lQbmO2IYSHbj+kTNA1TkBFStzl/cjzR72
yJ8zrlZPJ6Er5lxOBh4CrWNQMeT1Pb2r1w5c5nOOAXzlNTN27SJr7SWP+G78kxeDdYvlO2Djs0ex
qAoZXetv9Yj/RBBkTdkrhHcAaGcDVUt2lAMgNkKzWfoCYEXpVIKaDTbO4sPja8ErGt//q8K5SVvo
C4VTnZplN2D5srSn8kpguCad48/3T3FcYBhoIw8e9RtPBa2VlpEgg/FRUBQLc7eSF0x/TcAiSyI1
18LUCHUt6NpdSzzQ/xJvHQJvX/h1zNYdtLUez4dDCbGGuzahWKp3XELvnDt69BfMTX+HqDQgORam
xj6xUKEQ3BCqlaNJf0uyXMCvs/7qpX4uAhJeW0RPtjxNyMuRwGKeglfK7K7FdOnrX6cJxhjf44a4
llpCSdtkXzxbFElGtdShjhVKUJ0wr8O9Cmd4xofF3Zb51XgTdJl7xASU+Tz4+l7E1VmwXd80yvyL
L7B8aX+Ab+ba00V3VEuaJAuCKAQwfG72EkudaziVlWRfaLclPVhChHAN+mpV/mfS0C4LEdOZyxEC
XeWpFyWVw4ltuUYQJ3dG23EeAEUqFeftgIT1u2CXrwfvAy5POAH9nl4qzhmy2eUVLBhX8ikZV7YV
A0Tjos4zE2y0EUxSf0nr0S756o76zFJyRCgf/y2L8qV5XgpEtu+tnQdaDT7mVnNKuztBHzAiYBR4
+NV9Vvshp/OfsW9Voxz1aVb1CZUrQAM6OXJX6Eft7qep1VzokG8V+XNeSGDAHXLkLNcO3jjGRPUz
2jPr2gLndkvAcJdqoC5fTPyIoDBvz5NW24imUgShiMNjKSjItab/oPXQSR0fcEELUrvf5jpFRVGP
tjzF3jaiiUwITfywUqG0E6zy+rhWyvw+Vangu0fTCthnDN1QlfE/XiyBBsomIVZof7wF46VdCAUl
22DwgaaQH1SVbkiJqvnnZbEh8/c28cswuhJfb3oJHE+FZwZ4JF60DCdGQLm1m6k5W9nDaiyHphix
rqmJYBfTZPWMnRA30ub48jaLU6y1tgEUZK3PtaFbZWDHFjVtvS0UaPUTOJ7qoqUqGpAAH2r7oKRc
WEptohqpqsBqEfFh4ddF9IU9VVaDkz3hB4QGHsNb22p2Nad+DZd7MdOWu8fl+whwUTp5AiGrgCib
K4pl5e52GQc0vKx0dINqcZ5zmXgDQzTcIbxh9lcTUPtlZLtd7oEi+LO4oTGPzGQsyQVXUM32xt8c
ZWOImyiyvVSdSGmRLzCtNji50xmrrNcvbUYJdZLBSKeGHdp2ygRacnaOjU554Bdjq5pEBXAhsHfH
8m8EkbhSV6fgYsNVOUZcGt7DqEPq+3AxsZvUiOG9FPTZuREsUeWotwYRTkpsCqJQp202e3P9WDT7
rJ5h7tiuk6lHqoGGKzAjqmzunHbNMOyd2NKqS/vchsJyJmGM6mcEPs0wjWnnTi5NYaRvQ2iYguxa
vlXY4ugeccxeGpXmKic8U99Y5HSPGVOFPje5Sp+62JVWN/BQjc5mq00UDbMXerfWcA6Yrrhl84ly
1MyoCCzzEBdrcS5oSePdVjrbD92Yk1QnxT1NW6HH4rNarfqCg5CTliUPoP/VoSNGKc454Q67/HrY
57i0cCzb1oCPZ9OtmzcAzMFx6yUwQk15r8e+qk1Yx61IxFv1kVUj7Qse2xbK37nKLjhnMfLcL2lU
wTIK8BSWj3cU8RCOTw59IhyxprZy8iwC0VY+aUrXpcR0QFIYYC4otaMIWMWEcdB269u5kXCu2P1G
RHtgcm/X5UJYcM9VrOUGbwJWv7bha9B60D8o+1McJ3/VfZpkuUokGup6Oq7/a5HAfhgURBz/UeUW
MZxPSQ8ue1k5laTbLG8URWSFA6Kinx+58xY6lbDmOGWJcopx1kpy484jyfVoqCUt7BSf3mhjn5Vx
KrlLitCQU7T6670xPUDVTxgdyp79gGxOiGXhZ/pRVvZvEuZBefpAQqs+Gw7LvtNCpYs0yuenWzW2
qoymjVUHoH24glzgxdFdF5JHfnZO6Tw3u253LyLK0jRHyIMN752Znh1Yry4E1xQ1ABbPSeJPgAPG
6EKkK6xxj7B1BF0J+ZoEGRzakr3JMruMjP+wr183L/HMtgQCPl4Csfam7+j/ZkXfEpwGS0ucbINt
xIWIERoHFawUVbfMYO+3Hra3/HHr6SGwq7Z2Kwcx/5O25n04ahIyt792FS0PURrRhII3Eg8CV0HZ
wMtbPjHEjAbirSguX4IS5m5slGm1ZWeAltlpHYpN86SAu9vsEHtZXACH5HPLhOGeqTahJ2v77wlq
CkYmys4iAxEpqALuoVix+iB+QswyT9trnka6I2CQBH2e4V72Yij4ebtliSYfqhMSC7/4rMQTCNQg
TFD/7GMnp3Mbyq+1GG2M2sFENOVweurYm48jzEmWdWSDSvQf2R4Kzkaz2UhSqRrhgWuIBYJgoivr
neAkC3eEvJW1OAh02+7Ia9zV5kvZGfKqA3fqkrfmxU3xEu9vKDmibru5LxXeLpb6EXGOpZyBGgcn
kq0JQeP5qn5k+sxXfesupPBCeveefZvG7epyV1K2tb9ZD/K+oiRHEC1MMIvlio30ozcVAKSjaxUi
n7QYaeFo/V2FL+wkHXarsfhfWKjExbeG4JkRajZjIZP9vreYGj4Pcr2TJ0IPMDpNRIPN7WX8ASpz
usS90RFi/7zEPq8oLgoBs6oJLc+ugllj/CRMgrGpX+KRq6KYit2MfP0neTi7km2Fs4ev/UTZq8u0
HBU8fsQwfkqLSuBMQiK4SXNu8BfGG8yLwZcwS1H5WtGpkQrbJqchQD1dMcvgO9GJwsPIkMkRM8OV
K4oGSA2IY24nWqZNiINDCjpWzJSfSuHPKKxqZG4v4Ut6kdGecKVbtyzHGIHARL1OrWmvdNoCVPlq
WZLzaZaDl+QZWIj+x0t1bAs2+KAMsLVsJ0fvXZZUxbSnw29kFGEmrID4cfiptyp0M/VbSB0J2WTn
AwDD4MuzaJQL/TFdUyPUIt+QEGoL/GPNfMR5Ej9rLjt/xPuCpltXi45Szz+SObF5+/fvWT59+/wu
yY+9lxhQleE/wKL49rULdnPuOlxbuNNaK9JlcEcf+j6tfj6/9O3e9K3v2inQmo9rphP2NX/4IBZ7
soprifw88FXoa+QJD6X1LHXcrbEBMGzBfyw0bD2N1E13HRs/LKv8LWDBPuIu0rwPA84NuUxzQvAP
i7bk56RNSubLJwXRZUI8XEuGGL7mZN1GHiOn9FZ3H1XEx7x48nGofuuDYDPf7nnYmlH654Cse7Qf
kNeYHfeff+wvw+YQ7O03JsMUNrnE0oxVfPCEAJAKJ0jhJjjSBXjGtVcA00+hmmNoDFR08iGWx0Hg
+kQ2ioRvQYtEd8VhMjs0KSWxldSdGNrdImQhU48S0f0xL7oqNC5gNwFdNhsBdiARqSrUuGJYhXGO
lXlMvMx0gl6UbCgq1wMPjnLR1QjR+iEJj0RpZ1mskE9OfPhRMtRY2cLNneKYVfhZMUZS8yVf4H11
I2qLo+VHKbPRwBzmwgFAuwoj4HRV8oVE1y5KsAIB/ZQvAJGv//QYyj2wQwE1wftlz4l8+Cmd997H
/oGfmhqJ9bG8rR2OfD2GG9kgSfK73v2TGefQ4sITbaXXl/PMyXIF5WTKd9zm25IaEOTsHNzewTj0
/AqpcRC+OlbQrHx5EFKTnobp/rn2imnPSvqHvFYWYJU/Ye3G87qMc24YYnyjtTNmx6RH1lRy3OyV
GjN4DYMPXLKhH8JfJvTdfTdogpSBwvTt/xrUgViMVocMcq5oOSo9jlE87VYJ68stuXrSxfd55YFz
Bv9z4qDcwOdg3u3Z8ht2siqrVGZzV/H6O5rsHud5NrXWLC6C+tgFokOzTi+W/6apbA6llXzVyClB
mU/Edld0gZKaokjaBeO6bFxH18Jc1nKW0GG91AtCIxrOMc7lTKHajLoUdvCNaZeBYM5tncQkLGzV
mNw4CJxdtq+6kFfEBED2scNh6BpZPbcjcFs8XHnTG7AasBDIZu0WoVxcalltK4dfEs1LrL46wKrL
l4Aut+KNRlPmF9vTLRvmd51yudyaLUyG1rKFzQiGrY2q/yrAaPt4rTZ8dm+Fft16zHGrmtZ5nV57
BD3ZM0Ay9vw7u1alCTzeROEueQSaXL84P3NULiOZFRGmuMCOEEORyf62GdcNYqq2jeR5HDA6vFeG
cz/v87bQR5109/PQ8Q8/E2qutjVCieP5+2lPTuW4TWCJhBMTcicrlgrmtD/OfVa8plyoyIfu0c0m
H6IGkMk/xtaQeYnC6HiwVBPA1xgagsD9L9JOGRRz2L2wNCk6Z/0umgDYBAxTeTe72nRFroCjG78I
Q9jG1v3MFuL7K5u2UwOC4Ogb0OukgVegbPci+LnFcLouIZEJdM0XT2QKXC+/JEnTl8eumb6KEJhH
OeaUoPcgDVsbkSM0EtgPZ7xwYkBUeUm6kmOC+eV77CpbgAETmjpIyOzp0o6fOZanJwdnaQX12DRF
+guE75I3yuoY6xvnCEA/G9lMIS2shoHuqjLJs/45Ghony6eLsA0gMNXYhFuM1AipbYSCLfWlplmT
OmCJucQt3oTTyQLplMhMJHTORknkNXiyko/Ugwp/Kt+6rxydl+MeM7YcmnPtqGnf0YI+ET/3Ei02
THJwC7ZRcMpD064gwI/2W4xKU0wkthfupQ6SIcWTHZQrPs3+Kcni/zdaZup8FfiifgPeM0RRzjzs
P/iHOAP4E3Dj2hXAbo8H5wx66Jw5TkAKu3aInCnk2lok7DWv15lI3firsBYyuaXo3JEVXpWXO5At
W+4RsYJ6wbOsBMczxXuv6FlF/5kBFK5+rnyri8EoJKrPbOyrMLIb2jgwiinJ/4/pX6jUuTrmdj6c
VqSSRXGPigK2HccBpzHM6+Buy1weSXwxFxaQeO3RdP5GHROfkoysx9geqNMbYPr/Milkg2dLNk7Q
tm4q2xhGKbzL7KH6LXK8UrPXlnjxodAf46X30nvyDxl+lRhEKbfsCpNmBZPXZ3he8zeVntXAQwz9
IpF48J9Py4jQFKVZ3ZmMojrsctbf0PAZAAZt0dF7txu/iQcZKlqrvMZcx29s1elJACPtr71RyjM8
LkRpNXB1xPJNx0yZZ117TrJ9kej8bSG4ZkVHU4jQrnJf9nNtv4UPU+esIV3zC85TfseJCPa1JYBZ
50s4v3E8boIscJvK9ibIjr+b0LKzJe/CrJLWt7B06AZSLIxGTS+LPn0r4rHcHDa2fnnZy9O6DKUB
TpxwDjDPS7ozSGvr+zbb369PZQGDJLTDFhIt6XDV0hcmTg9D+2ExyZwZyHBogbI9UTU9xqteKXWh
4g3NwPRSyq72zbLFw6qtlTf3y5vIw96Jdy/abgMP0eMOz53wHrU/pUNf1wLBIS3+KXM9Umo3v8he
RqVljwKBPPzGhe21dpMsPfFKd3Dm+1KjaK2cCV6+L5oTmuDcCDu8JB8cDVFk+skfsDYP+g/xqvU0
jfhwxkLvj4KBSE/Ctak2ZEMtqev+rJF9d84qSI1tzkbpMDcfcR3CJXKOmenBzaNQKvCZMXZchvqV
boPSPHtW/OmtFws9+XBNwTt2zaEg4mkYZqNEoAkhe3DH+uyIGz3ec/YdAs+zLX6SnGgTr0OEBoQV
FvpnawKyw70dv+rDFXAB7yGCgU7qZufoiuqtVu3UqABaLBDnHDEUZ2yyF0a7FKBtf5Hvz/xv6fQH
OZbcaCcyQ4jiyLoh/U5zOXehnToQTIM5mToBPOGFS/1u83vxJlQVERFC7/tusD4S5vK8EHZ6ILgM
Kf1UY41pdP+2NFzF+XRWe3GDzyCLo9jGWnT+HOnI/qmGKfFhW3Q1+hEmN0O0JYed6GZdF78JVNpk
gjcJsqvWulXnJZ0MD/zYHt4IRDMfXHAjDArUzKYyHtmKNoPsDODXRn+dadbxBj45cHfKOkipmgVR
1iRG9Il1L53zl6/5jGWs1bjqEqYwIBTR09DYak7hMlm0OFzc4gJKug2E9GKR4CHzJfn2FdjNFofL
EjRuz9c4bEOtN9SZTVIipW2yEQ05LsdAIeCxyspZchz0XIJzhgFWsef9JSk+wsqgZ1QBqZl2rJzG
36z6v8+r1Q3PDtSakpPQqArvtJgJlo2LoDV+hut0IlawxCYvVwpv9EWjSN2Pw0zbq8nTzESjEzwD
OmbHs0Fc+WTk7yZVjbGkrLguB6KrY20H6PYGq8XXgQMiSVRTkf9uUplncxIl9HOdftPZNXXpA/hl
Xd7jBw6clVMDjTc4FCxq4VYKrxKlATGQncPmY//yVFamm9Bz0PEhXHMvWDmoSCcF3AUowb3ymik5
gP4OQO/PL40GawyydyVsWZk0b9AuzWqYjwdwdaon2Os97I7/ki5ihBG+BHjzTxQcSpHyTo5h3Cc+
KdXHUmaFswSg/0cxGnMRugUOnj1YzMsixOGSRQ/l+zNn6Pw92HxZ63dM55uqSGbeT/IRPpPtOJw0
TUZirOkqpE4E+yWPsXtfdSz7Ic+Uyr4XFlAo33emmxX6Yj+NL7U+XYI6hCOqNahnUfrXLPZ2La86
+HMgYFalbZgZZ+o+hAHvyZAIA51UxC3rzRYj/XPrZuQNGLe63s89+2D/r4pdSOvUVjxM6R24PkUG
V9dRiMGwfg1MfGSSrqeYLon7vQfdELkn54b/8ozztECecckELrWFPXCv5qVuY1nZDqReVRVwuPR8
AD5p6OrPUPJmNXgXfGzyEcwwe4R6uDZs7L4hKlOIwSxFX6PmzH/JgqT8XoSMxv3HL3iYOeOL3xay
cJMn3mPAgsM5PxBUQ5L1e9HGYNb8K+NaU8Hx3cJnZ448NEl66hBnbYmI32o+RXuNVoFdR/EP5hrs
s78DtwxXeU3HKxznvINjBquBlAUDSKY1pAdyA5VQFwGuX8Oi51of1ILKLI3ZSN+SlldxjmQSZeCI
uUjYt8Ep/35aN8139tZJ/p4a+iUSZkbw9JZ9TzYC/gwCXRAg9ZcBt4/n1530ajmV8+Nm6txcCisq
XJWtnxKYHCXLHQlpcoOI8nxZ8Yaa4WA4VyinDNnAPebt2Ydw9375A98V5XYWOldJIsNeRoZmsWCg
snlK+vYnsmav0wjRngu46d8aF67tq+usffkdf9gXTAMc4NrqFf8Oo5ktzp5NdABQuQfrAx3OItI4
jb9Awm2v8rhM/RmK7evXUYxJwsTsfaLFgxug1HjdTf5OqAmKMz3WDsRd6IObt1wM0ecZqlJJo+3G
ibGV7vGHm8qTvzAzRHdEZVgg4F3BcDokHh4V3aQ/yT6KWQuRj1mD4h6Kl27Pg/qD8U+9ED26L0SE
p8nZn2VxgRep3tuDlUeS5YH2URBtjDUAyixKkPwrsRLltIvqubKq8jEDpej3gZFMSVYADf47/Ckr
0vsXtA1VTcwCprFbnU/jepaSPUkgHrfIY/DfyliQNbMDK21y/go/rzyN/te++TBhMxT4xLZPBZwh
bO67C8wFupA5HAY/U3RcpkgTFnYQw4BNBf9vyCtTLQzCTlHxPM5Fu2SGtk2iQXTRsOuw96WhuXbE
wG3aR92MZrci9BLX+ZsySADyFSer5jZ/fotXuOkCi37UVN1d8WzlPuyJ8JsDvY56jtU5Qrx4YSpO
ImXpcOetpegJC/jSS3eAdAeOw2AaqutS4Xl0x34G2geZaa05ADwMenng8h4K/DU02vcGxroHXcTK
+Fckcnw00PWId3WwyQx8VyF7pRWFEdOjBStiJvx9xYTIG2/QinicjDF1MRnBRbjgcogS3kUe4u5V
7i29poPum2+9k94GMucOmrv0f03jnGXdHHtgqpQhIjTJ2+uJTeVYfkwEQ/Hguz/BPp/c3HUhd15Y
bgrpeDjluEILjJfhFGstayDepxNXnoFZmU4MS//Bebg9y17ghswssH5dIeZrzlGnwjz2qgOUs17x
rM9T0SmQj9pM7MDIrRyse0B9lbEtEEqS8fO8707D4O65iSHcfHTQTlJIKlWrH/7wQaQqhjbkevJj
OtwUYFAZkaUhz2u6O9nnXrrs4OgSwJbeNBVS1bN+kJqbtBrNQVMplN1yb6Hyu4ZxES5pKnaqjxR2
Hn1zT9LbNqLy1aLhR0IB5l1vDXEwduGQFzi+Q9Fcl4PxE+n5rm8ZIZUkhPyk4m7Vunx7Rf2ZzTQQ
LqNWqfgHcgX99Zh47d83DyW6YtOXJLEHuIIebGUiZgeFGJJwDgp1L7Y97IdoYfPmCDlddSUWhSnZ
b2U2g5/NKqfnCtj2w06x2dTUX4hnKzObgiX8rB7jPZ2Eso54ReUV4I8eqFS+69ux38TIwxDw9pr4
AcWwAhxh0CG9eAA46kTIWYP7LG4oXQ8kN4XQIAngtL0rZgEOHf0qt1JfPsi+Sdk1TyD8BtVzmBoj
ZSGd1HcFF3QLkpqiqizNVscYRE7uRaYiyhnQnLDO5r2Fdl8KuCRprrTIGgEVVq2TnvpaNrliKLoq
r40mqqh8oBDQWIdBZo+PSJ805o5r37uN/mWX5X1IsaQx9BcyxcpfsvCto1PCuARG5HByStsRMdIU
fXEopZS2fKPcMh4+BUwnvchCwugqlXatCAV3EcKJh0QiYt1VnTDQr58WgkDIFGV0g91t11rneNEo
eEhvALd1DxTNgk/CI0KM7g68rxw82Gc/A1GJNzydER2p1JVjVZINRnfWTNxSWlyeBnKGm6fL7n9b
4SQHSsH457cDROXqDudQLS3G6ZWOvYqWVlc5gsPDpASt5dyICOLW4xClD/P6m3B/6JYUYlR0rvIr
nn4QyS5jmEhhi5LUVIO1INlhB7FKAvSyX4/CrUsVzvkH0OoIxLkMpun6ZK8xrLPPWOB1qDSVzW6v
XJLxxj7elRDDrGK2o+XkDDuwG9d4KWycohHumKSm4dh5qJcAyhcrsggFhr6+cfkS+JvFeduAoEB9
Hzh4xnceFl5JpW5jlqKD02IlQ+aeP5CF26WPmeVnqFrsSva561WZBWCyfT39LzP2+fDYbLguGCGy
FQo/mCu6zeHv+tMl7Ls9lFXd2LE1HHz+f+kKopn2kSRVOxcvtOi2Ycs5AX9FqD8QugVENHlafJM/
cLsFbitlKzLg2vUsdPsaWQvxxvMqL8BWte0xKE4YNlPJ60ZQXPClSi47J5biMzzBiYFjt9sSKt9T
+DQad+7bU86CWVkb7tZp5X757axRsMp0KDj8GIZxY8s5JBi1CZ5lj78zcZBRYrL6C6jVhTGnFbul
1r3tFDr/QbAp4veXlZ0xI/eS9SfFVmhWhyLPL1/sr8tQmnLQ9Ihh7aJOSKMjHTj8d9MK1bfWo1gg
exXG1/94wqz77dT4UrMNUhHlnlP6GiYnqQC26GgMIe1Ip0TpVrivBQ6Vc1ezEPRFve8oliJptKSo
2p1yzhxfv3giJuFxuLB240x2e0BU2lESopk0nXCcmtapqwMcsVZblmAlsk3L1Ehr4C+S8yJtbPra
azkbL3vho5/JoC0eP4ddj3qNmPQ1dgy388OzsLyAbQ4BKyR02BglN3XQ0ZGILBDrM6zm5ftxCckD
lzDQbde9uRxMQoUkcdQR2UUDgIa9/Io4OTQQOSBbSJCtPg5isYISdMDEnWXKCrxHLZZ1FDD+llim
u3gLGL3k9UmUmjZk74xUmUJd7XP4LPAO/FAjqyxYmAD2cWWPWav3bT2ezyUjeePb/HtwubidW3DE
T4M2yVOQTpDytIkIGAv/Br/FnMamu27iIIuRsgWAlzG+1m8dgm5p/21WxXf6YIfB4UoWQHUlPmJP
hmwrBduvpHCiewUR5jSL/iY7jg9jQpCiWP8WI/z4q/2yH+/jbOsbzq90LYkKWvFY/J9DF7umLySt
3hEn+me1ph2EzinOP4CLh5kiSiRNTU5HSZwdipVOob5H7WzbN88TWe2T9Ql+Jnn0dWwOWw3DctjG
33qPWzexery+/NtobenVR5axRMHn1RZ4yI70XZThfP+Zh6a25tD/pOCyjfW3yyY8lPq9vl2dtEr4
aDkDdH1Wm2bKeGfXvZ0YGZadaanYScOZAHkcHbpZaT4QfqHSvccTTgbW0CnbWs5ZO4s34RaQ2ufS
TGeCASYV8bcbXKsg/10eLnHewaV/7S/5VhO6tA36Ky71yRSpxHUJjNrAtNgSBacvtqK9vxaWpGtu
dP7AR5LWbZAtf+XJMWdGibD2fK9C13yILkuezaN4du2HB55QPh3+DlRh8DS+vr8zLeML9ivaw50O
h/8N27tgQ1GLjA6+2Thm6FjWJENswTg1VnX2JfglHnPd76huNfZyi6kMe1Q5zezlnIbCKA3LBxd6
ACzPgzgH1kNfdjMAJqn+S7+F8RarSDEKCQdRCngVQ7lFHxrHEMLYbbCYOQGpmsHS4vX1oH9FxBcO
L5zFEY1UmCB8JGQxX/shzy/9zMblQ6z/ABnSiXhVYASfi4uWXVJYuRHZ4jPfzcFS6K1euSgXIW/k
eD35VL/tyUpqAb0oHNhlG83CN1BowSVuz727fEN5fjvZ7m9eCq2JDV82P92en8X9HqGYuFKqA1bM
q3xKRNjN+Et3pSIXp+ORrxKQC55oAD0/EB7Sb9DMHBo/ClsqcDvIOBPkSafzeOrqp3OrefP9yUoD
KwqRo1JAOa7BVRVoo2aTKmjWsXySnew11ksFcywqGDvS5cZVPdRl6FJxUr8dJS9RDevrnJGyl9sS
4fuOw11+Bv3AioeaBDHoXfpsd9bIkqetLWtYZCXMd7Pe4UxiZufxAupJm1lR95sK8QgWFHaMf0Hb
9kYu66DOIKRU/JYaBqkxXGVmph709eYfib9nYkLzPwB6R3BSy3PqgdDMRR2McChCO7pXRALhlDar
yUeAGQH63iFAfkgmDHlb5onlVuzTWGdEk/pH6N7WcJ//ozPTuqLN0XE8StGrbZdUbbhdNh7PCK7B
8MD4BqvhBuIwyhq3HpzeJ/gfYvfSJOlvTkpf7FAy0NmGW2jhPAE0MrpdZFbMDF8ZXmPxlvESiCn9
QmwQauDaF0iPDlTariFTJPqGmuKfTf+9/2u5NNBiQBbX6UclQgJr4+n7wo6l94E83Dch7oGHko7+
y9c02Oui27uIWoLvKJAE2WHkl/VbRDjUGgAyAqOKkoWZzsVXRi/+oqh9bHCE42WndkIf0XfoK6Ro
8L9qFOJbWDHI1/eLjMU0YrhUDiy/zoBT9uCKLS7O2txMHLq7sdXfURIhKW3U+af6VHbwL5ZVUGl9
VIKlrPVImslMoE/UcTvo52sXoyHD5BYIxMh1AeaWcmymn3ooQFO71WmzHlmlBlMyeHLEt35b5lQy
TimUA20D3VV/WSf9Epl1l8RDRyLfjX4oM5fab1fma00A6gef78lSh5uClyxWPwGorDaoNNNtNfXm
SZlEGVPlfF3Ncpv6yn1HbM2CZeItF55qofqeNDrOQ7rVkbAbqZ/74yt9gbmka5bV6zHb7qtPLrh2
z1gcm1DcuKjwN0VYIWkB+W5kJ7YUYTHakRVAPylqwP3eOSoFbCLE8uwqJrhXMEWbWhUAjhAZZvaE
IqbnVoRixPG/XwVMv7TDN8SCifGEc2abmqAQ9IxVDkC8D8tym7FxZfurwY/hnkZ1N7Fyv8zdxT1N
ZzO2fqkHrxQvDqqlGa22H1XgWOtWvC87P6WbSPzhS/EGx/ne1dFHUeXjlmih6lkbksfcG73L1Bja
bqaWYwp7Ig7tHsvMTyd8foE/70SuFZaWoeev6Jm80sA+EIFleuff9qs6nHs2AJX4lKL17KiddRHF
28+KRQ/UoiUStVGdW9ZhtL9Z6CXekZeBxibionqv4EfY3SYgUTK8ESZdfkOGh90ZydovevwEWT4n
RrtF/0fnEJPCeiPB9gbQCB4m+M8cbSgJ8WHykY483uN/LWiNmmgJH+rSfkYAP1rf7AQ0t2FrdpZ2
ykMg5nq54juAbG4aX1Ze2mdy8zsXOJdoL9v+unW/RNdoPJirNRKCMZhmf6WTXfWMRcqIjqNib95z
K+YhlrR7xYcrGhO+IUCwfZJFIhgzn/RjjEiFgEV7F5rL+uC1MXfwyW2ixNM/Vce+vOhwmDsYjSp2
pJtAW9iUiuisaZRqTSd0AM7QtnlzlNR55iGlvIP/5MS4Jb/JK763BFkXsa4bq0Jtj2Pms7yi/UnQ
hvtOXdNwyBS0OgAcuApDNOpET8FCIOq/arC6EAOggLU6XnwzHkmif8eNbAiTOG96u3q/ZV6Xde/C
1JGZEdQB759ZYApxG8w0S3abrKoYwOEbp0lFG2FMAPNsjKx36e0WXAhKm8vji55LwMr354WaeUB0
KObduCTZjDqkcgdcjYFyDTi1+2sD7+G1vXwYrtQWg9oJsdKDs4L1uuoZoKB2Iw2SH83Z5pQFW/Ez
pY7k2m2VPuCGCvPyw52aJYXDCq9MobGBfpZJ4+ReXFOpoNs3sdRF9c/tCT5b7GWgKpLyftNllLYB
yUOPiPWPTEqiROivGfh8SPGUIoKoELsKHeD/y+K7JLB+nHov3koTKF7eWSZ5bzso5MUExfz6O4hI
4DPIf/NaA0yrdzMJAl9TrCCBlPqoPzGFy/kb5VXhrsmoWdEaAsIma1fbKZyeQTc9sxxfUTJcrKiq
Csdd5hmZFpZePrhX/w2f/b/BJxYikRoeOFNNwtNCblJo3CJnBM74L+c3/cIk5waS0R03xIAnAqwV
31ksXW6Yqclv4bVK6PLHiLvlDMAydcsKLhmsTSeh4UUp4T/jZgGqMaQX98meF95Gx9C9GCneyB5i
f9dO3BZdazzAf/KmlDYx38EowKM4rOvM8TNnbkTnd3DkrO4w4pv7/dISRL9qjCquJ3ly5baqbDu6
Go4hDi4GcZ025Oqnt8wNuKHwsH91A6PB5tWWtdQ0hSeQwaL9f901gH9Xsnp0b4a904N9di+WQMME
98x8gz3Vg/RJm6Wu7SUROQ+OxqCJoKd82t1mVkXx2ta6HhvmNtcBNTFJlViegKkOHXuKhlCVycI+
/yj2TI47yMcH5YlmwrX+Xow5gsnLy/Xy6azziF0kKivGxtxcrDWPHUznj+PqR68w0L/4iqdHTqXO
mBq94F+Gaxay0OXsCUfyBKZQswf1hPZ561FodW2lFEQQU5dqGLGZips+yzZwYSYYsVBjDuPfmc15
52CUTJuvu8cMQ1HyzJA16G2FRyoZWtRTqKHG8jFINAOtQBbex1TKFSeFt4n84dk0KpknrFD713H3
5Za/hyVfrwYuCfm++7pFHkQdeT5j7jVygfglstrNvTQK26p4Uz9kIaQM0DH3QjEWdbo13CfZOSI/
xfEypkYyzUtgTdhqEB0fJ2u78pgROX/nJNEs5/JKl4czYC7q/+9CV8xW8x3HmAAM+HaB4kzEj3uW
dBBfZ/+WVsfg7KwXnr18WxWz71wDDfzimtnqS5st8L2oJcccFjujVpIeJvdxem6+TCmsjBDWiodf
CZKxMlLTVt8Gs/tljc966/sd99sXCDZLgaJkq4e+JUBfTs7woQSTccZng9X8j3fDSiDtT4wcysjS
HhPSbB2OD2egroyVoZtyI0SDEkJsligv9Z209xJA6nYMKg4vRhzDkXINYhFqOexZ+QWN0q5lCD2L
y58b7pR0iocVygIfCLgngGlT+ZQtEU6VVPB6DzvpS1WO9wt6w0xem1P0ArwFsj+PYR5BAWUMoTQC
ZkmLgFNZ9TgF2hH6bHvky2qxt3WnHG8hUIb26cXRXdkM2KPMSssmnLMogPDljrSEq9vY02Q64SKZ
tnNvzN+h/6Axz7NLmxB75LCO3zTcBT3ORFInehQAFHzKkIEt82z00oCOhl75E33aDLfDuYWnagMd
4B3bRQIYvXgjr5NoZDcdqS2JgNIrk0YeItmyTnF1j5MgQTn/1qzHhuq+jQgZReKAC6r9CujcS1Fw
Fwurmbs/j0hoW4K/Fg/qwTrgQfKmqoRsVH7kaZAKhyzGkyJdIsJwKlVS7dg3Ws5C+0txs4r/3Y0b
wiJc+z3d2i5pqnA2/+eWxZeg+X1yvuisnOgpgf10CYbq6GANXtLD21O/J+2dkJ+OH/qLHkSBjSQG
fLxQLYJA8xOPu492DymOkgWqaasNGeVBSzwLHFaLnFcYRg+E8X9suxjUfo0C7jYGvJ4biBk/D52C
QFd4gJJ+lbJDtfP4iqzb1YnLREbtwZLP1dAWxm6iV5DuB+TZWl1Q6oQ50Cr6SOm3Aran1qb3+rPY
6m0dOV4e21Iuuaoa/+o/ctLAnbzqnmnVJaS+iROHMUEwF66EwMSxxI5onysuTESal4TYhgofnYIX
RgJATPZq/b8lG3qtIRxHduWvnzzWY2WJURIr0JBqyIviKJEo6iuBF1ZV4tNFwGDwSkKzmxNtA+Pw
kMhlpQVErrRJ+0C4AOaXzZehCqBbtPcyheyQ7zxq0BnWqvaaerFGPCUHR5uzfPFvVZvitkyM7Riz
JWNjCDU1Z+cOXhC1ErU6UhllzdpRA4d0TxVGiaAXEyWkUr8I2CTD0PFs4KzopoqqpCB37NLCWbX6
pdegEUSwZHsFTinp5vCO2ohBCnYMSRXfExZOhLto1SyDI9XGpoFBWOKadWNYVLfrVfSMycsYjSd6
foAcWDNYxrZ7oaUujRK1dIfMgRdEn+4fU6CBNCEmSiNhxNVv/Ti1poDuNYdavoehqwy3lGOCyiW4
kt/FmfhVK0ncnnKxLCFw9/KDOV4u/IDYUPCw/G9dpEZ93KQCv5pseOvXO/k8+TTYifgDzv5GXgf4
ZqWKGn35OxN5Veo54iOo3g22lKLav1PCHgSGT3OVpMX0G/oXV6r9SxggSU9sdDRzj8ugEb4tqFUh
oRI3MpOatkSztlbHdn01o+A3089xu+KWHpWDfUWrh1k2I1a1c7S7oubmULnoBOjZZ1pgTXniXIaS
s48mFJUhKuPrNqiylc0tYzWz5flFAMGAzmn0mkS4PaDOMtj1+2ycjEPdpTW2mPwApJGp7WN7FuRZ
zBN3/Fef39CcgvRwRNKZya1rCoNllL8moNMaQj+4Kr/kTh5gkt/ri4z2XMqIyo15iHLHU0jWDj9K
wVUtcl+PDcROriHUFy4Tc57Ph4eycsh/5Qczuc0PUwuYTARB4CtEp4O+5n524JDmMAbchWvi0jRs
45IU4IIt/kXuBhmvtnSvKLBiSdwrJ5+ApUeyNGpsnN9pVtILFYo38wyfEkXmb49GJo/0FqGkjDyE
nbCx3KudZKGWzYZFqw580DVc24d4BGxDMK/mjpIe+uNFV1/Zxlnlu8NkOnDpHiGN6y+Fyjnc/Z38
BVleECHLyQowbR2dp3FJP8/6SQGiKJemvYcxUdftoi4SRyaLOoyR/+FmXCLCCxAZ2HmE0AwSviTk
d2doaG4TYrBNJMLmuUMgUegKjNVpx2kcPYRRkTABUgiicXYPhKzMeq+j9NZP1sYsGS4koHcItttV
+Xfxo5xdy5Trs0cN+h8+Q6Sropiq5PVylvaB50LqHwM75quRKC0p5x0oApzxFHYfkB0qBrbADvcM
WExcJsUeH9eoYb/idm7SU/dM98SA51a+E+1kL7RYpPX4su0CsXi8mNXLBETEH1TubYutX4cH8Luu
LK6nxJlGxEjN7AE8kpJ1WZ9YGgZiBRC2unks4PEbE9KSMqNwMmRR3epemx04WkW0xsP0O0yH+Ins
lrDNuI4d5D1f3+s5pqFj2zmg7SoJMZ7BFMZ2MV36d5mv1pu9JwiRQvNmOWIZPa02/+NsfebWRadt
dYwGim+STLYQXTgm2arKiHOJXXzZFKtpe1XaTWWosS1uRwL3W7T7hOIs+1TXpreuIutV+3pz8gQN
upPxQga3pF1ccfCMWv5I/4+pj1E4+mHQ3we4bPSqh8Fy+T8R5zZFT/zfFLiEjkriTPyScCW8SMGs
5e6pSSfh00WdLnFWo8m4qCSjnHLIiuKSYzIPkc6ydRZFU5uiSlgXCpPEQOhAMryoCHqjwq7Jf6tl
6pyfJCnpDG4xMImaAy7PgAKPOrCR7tZqOYkI8QLU/Y8PTgdz7mASRvOovUBaYrLGbl2fPuNaxIc4
NC7Rqg5Pdy7t62/4BPHYdg69UOQMkuG0EIX5ZQuPh8KIzmlx/85H7+I9tfY7YnwObqk5VtKWMDRV
S3l8cA4cfweIEd8JNoJOTmMkf1Xl+IJhwtLkYqBhNAFDpTYwDQME3GsLVxjhpUGj/P9ztQDUCHJ+
P5YVLJavE8DLEBU5NwjyZZN/KKMBUcnZcMTcbii50pSA4Db6KibtXZLsKUURqtINHMUHesitFvGo
CsheKEyA17Ydc7wrcC28yWs+aF11oecslx5PXhS7hlXSNmVBpKfYyCk8oRDkVe7UPc1NJoOIZHlA
tOrpoFX/n/nDx1+6xA5g4pjisJv6isadAZ8nLetcoVf7+sbwjsOQCA9g14sK8oNXASTwZ9PALnkE
XzHb24FLaWh1ytCwWcKXeBcKh8LRvCSaHGsmG4mYl1rTI92VFROFGa5gH/PaDdunb3LX8Fx89Z7z
HwedID7aZ5xKDA07kftoCcCtZsumyCsDwY1ywS0ApXS4qTI0Vi1+J08oi+xfqN4IDa8ksuCd4m9/
3QOq5c7OcRPFywH/nly3OhU5Ks17yiOYxmqXM7IyeuRJtktGFdHY38Mg5lPMMUMOBY8P41zCouRV
MyO+oOAji4BGdPcN2Bc3dxbkrHp8krsgp2xcbp5m2fF35vPe6eU4LxtEEKY+Oud5c5ugyBsPYy9p
R6WIv7FZt4Uyn4wKnfVaKcxAVb2+OY2xWdG/XGC/2+C3cp54gGYjLMPjpwzqV9iGhJQLdC6B0sU6
nU35Fan2zXA6sfY5+ctAf2jtEdZASky/iEI6V2hWwb2Ehuj1Ptms6nzAQkPOrNw8oOOjBS7B0xxi
ApHVa3eQWStr2nQclAOIgQmUv7ve6RhHeefuA2nzOEtJUDbtN4XgnXDiSeaypeof7PyBJIfBWrwx
JE3QR2dHMzm6XHTwzjB8J/h1xFCyUda4uAozY8XsVASeFT3VmL4zDW7pQ1qtPJk/Q20pS07lys9g
UNvKekPNLhogGsrdHFLkRQ8U7rEyS+kJ6ApJMQ0S/dbAnzLVBZ26D0cYDtXzP9KmCRQcbEoMm7Xs
sw+p9Q+QwLV3MxPoN4CniDQtpOW2FA9sl5OIm3aiI7p94UX6xGgeLbYeGSb/Fe5iydTP1fmekSf4
U+wG7WvdsMLHFKOxwvWZiB9EZzCVCdVm+ocvstw65/ZQZXNhMGfSdx3G+cgPDJceb2HBqoaoXKQJ
/1RxKt/Sz+aFczLp8Bp8tRyeunFXGsAke5l/0QJ5/PFrZXNCLd0ZfnHdZpDGfxYd7T2pWQ6ushpI
uu24C37pXPzwvt34YuNeBgm7a9tGnk+NEabQzvPvM8fK5iJrHgt35i4WS+oWxTjjB+hmGWns2TE/
cEXq3UGyrshH9WGhE/m4YQenO+jqA+hEKGjMjmhLc3BOkzTKk7iHradGIfAxokpHauXWvxWvBVdX
MYeEZtf37LPt9JVNZBm60H0vk96fax9v36c09JDobmgJR3paYSB/OuBJQxJDS7V4x+c2wjba0qSu
yzqB3oLw6QToWsO2X2VnNDpwWyUyL1uhcAa+GHQLlgCjbmctdHaCqi4BdoZACX7eea8FNuXFZMHO
0EDeHA7GY1M8loh5FdigVYACuBaYklaq3WvZ5gjS4CrBkRhXoEkZAq0g3VmPH0lIYdHf4SZwkyJy
uDfDZrnWcl43aE0EGRS4G/fMRqecO08PRPCgmsyfntfERVyQr7N4Bg0QtFMJ/Z774b6GSHbwvERM
dLa14VCYFjkdgO5aa5vO5KFM3mzipts4TeY1sqrnn6FoamR3cG8ayt6Nm6FZatfZUg9rlxPfVriA
Mrtbvy7dIl4LlcOdnwk7zZokVB9piTA6a2BOwdlsdB+TahuAzZr4upjtF3tZsGNU1dgaRMclDz2x
qjhXDMWDa51aPzIHIDyLc2K7TPrcqazZL98dme6T6ZfBlVfhIrpPD+j2O1gVAWdosFcIsXaN9krB
TgNxm/r1jT2BpZiNP5Va4uQ91pvZcGofj6FIGSfie8zhI6HK9TA7RUvRgQBHIrE0b4dr3KKgBp1L
SqT+vcbVOo9DUqmiC78yFetV3kBArREZ2ytjGstBha7qx1Jn4FVid2Pat+SUJk99nR+M53Ju+Ax7
HyjjQfN3SJZPZMXjmv4G5SGvsyXEghxFiOzYH2r3WsTuvfz8TKT1mlzqqESrVQT96hRcvtSd7oN+
ZO7LKraToFnEZej4VnzAS+Rej16/7sbigMQeTQ6qmDNRMleAh5ME8ObIk3NrDXyT3sTITCsoov80
KJ6gcxBb+0Bxug6s5y3qxesVShy0kwOAaSFC0azmXukQ5NXZAGDUgbV11bWxt1nA+Dl2k5M4wfvm
7mHk9JpUMW4rb5YI3eGM2hskjYM3Aon6ZbuRcx3mmO2elGNWLVZe9ScDQUEIaR3l54SZcUeA30rA
fQ6CbnY1QrzemnleB8dTvF5CRe8nX2C/xvY3JyPUeoH9MGrwOeIl61mQdgWMPJeQtqVFPTpptaTC
nJ5J7Eca7AFEhVBXVw07BXSzsiICUADvWfwnZ98Mgffhhw/wgSZzxaKFMpWXoWKsG/nbz6ZLhQhI
R/VET160Z7YcyeFXn2mxclWLDKXmcrxCNlG3lbrjHFmP3Lghe3myeVP+FXOZymIvatu+p1w48JQd
/r+66EqB5Ko/hZAHI0tFMIFEJaWCQv/t1V4aTB0hHemewPUlMHuuEbVFmukTqkjC/FZuDo84iviA
Ly5nVrGpfyT8H+jSAK8I3A0TPAmw0Ao5RDC9vSsobSjQqetIzE41/iSlH5SWPs+PZE/FGUNnP0jR
sLTBHVqWcFq7PJ1/BDcd82pBqYSIro7rYuwMu/RPGstfchywfpwa4seuPIa3oiEyTJ8GW4idBUYb
gSQzBBDpj/LqEisR2vWkExpy++Xv+2KcDJf7/4aeFnbP8vqcUQZRRK4AAsPCtiMDG0GdIk/pE6OV
57Kw54pBpLvNqJMkneKFrRloU6sU+d9cvSYRLWc1s0fBy681Zg6lf5Do2zsmRn0lhsXt/cYs0zTD
5fqxYyogPbQYWi9mJkRHXpFi+6WZGkmYzwRlQPgEXdZZhyNsBAjjSaogL+Gq+uCQAUwj8I9C+FIo
jPDvw2rnjyMo2g3+BWQujQXPCGF3BteId4A3drNYf1xtBuXtq5sBqnx4EPfQu3DGwbAwoNaKBtnM
FctqM4WTm1D2zWDntFsy7cjb/iSd59lqPKf/XuCH2emB3W5pqbEx89EqAsSaqUKpWTqzgo9cZXGr
Qrnnk9Rzoqf9GoVqsO51/IQEGNMN6FiTbgP7x7/j+Me4MVx5ODY6bLpz7QH3+nIxS3XPJgripILA
wZuYMg80wu/+HnNezvfkzGs+wRJsbA5Fi+vnUmS27XLYyQW7LYssBqwbQLNOo37VwcDVdpTl4zYL
y38pMTWVxV/6kijKM61w7sR1mVi2tokQBrbR0K8eIAZ1OxGnEEhMWjgArH5y/+wott5wjsrbfZWV
CWuKz2Z1j20VVNyShbquULfIHIYdiLtjbsVavQ4dka2DVeisFu6v+bNSwXkeantG6JrH3pl1Ux2z
P8hIfpKvDejpOywFbiGDKn0mzP28A9HOYzVnxrM5qV/VrEfIxgXWGEHmqx2Ac2pq1ER6sjHV08Ga
B8RulHhMfVOgDwv5bb1K4uYkOSOelupYHUZx9oH6hfquKP/mqk0/k9NIeRnX0rGBVqh57+4TTARq
WmagvhNAif1/lLymyQiRtsNhAkaYz+lZMAF3q8Vb8gN7elv/SYqL2fv+ecWYcJ+mxtymok4fKT6P
0UXgjRtyd4GAeK4+eh2dU77KqT8Rk+h4oWtTENmbgC6AVW9WPGYDWWNzVQ53bQdzMwAr8SVK5lIF
F3I/aIp2f5hRx0ZraIeQIKSxKlhQq6kOYr61yz4vq1Dxu68AWKiSCYArpTbumkePADQ98Y1ihB4/
A4rDgj/yXw4Rtj/FPkte95IjgpVXXcya/cLGwP+yqpKXIOBa7/XXtEUCgij0gt3g69kMPIQo3Qat
jLx0n+IZPyyQzvlIk0XqQ+iiOwcLJEQFxgIkHZ/JrXlJiUoTz9hZvBreYGkEOTlTypP8/kBiLRn/
ZajgN1Q2T/59ixuzB78ESWFVtTaUU0RG5L6tMyW4cJ+nUKwaLzzI1zCwr7g0FEiEd6akYlg//MFx
yShTRW1CgoSH2lsQej/cmhPrl1I0ekvJZtjRdsAB6hKItRbW12khcvNGGFJRo5U5pR55C3OjVpMf
JRtw1rTNutHGDeVRTCIaIQ3WeWkXE24Bf5dTy07sRlLDJ5mg1Ofwy/08Rd4ZXP/h8cQ0FsnpG2tu
gaScxqLi/QOwnfmuOL653WdFAv+CbK5Nq+eJxPUXRmczqcQZjORoWfyAPObuLgSx6Q32BPi/h97P
Q/5upAJH8zuYc4b9qhPiOJD3LhdMEtqKEHWRgnI8hovdTXE+X4JpHQyYtQxr1uiuNCNfooYb6gP1
fpAfCX46KQWB0F7kOTbIvW67modEHqbk8zs8ch7YHs5zM9sBmPTu9H9SgEmKtyEqnNebpgxGjWyw
uTyri/sp1qneBMDazMRFnWN0z5h0WfZjRJNIauJ4MG0Hfkfu3arCAayJxpS4Tz0Y3IE60uayZQXK
v6YYOBCi1dsbwAjYQaY6sfMKVGRD4psDTsxB4S+NZk/Cdnb+MoRSUNqqlmHro0yljimSX6Bt4lK1
tucY1Y5cbxq+AO9TrkV3DG4uGw0cAs8hqf2UmF5hUKlgKik/mURDVCoftsneqfLYbDI0bhDSDbgl
bkrA74Vwi9r9zKTnOnQcXsBEHWWEQvGMge5x5UCEqmcJViMSbA4YOfEJO5H5oEGK4GKkjxhl3WTs
/Z7rJy8bbYaJaCl7YuG7O9lMms79Ew6tygW09ogXEJYZoHIS8pZIRrIerL3EG/tRqkgSr4n3bxCF
t9I2fhOAeyI1r5QK1WQcLzBOED6g6OBhJ/u1Y4z37bR6uvi9yKmPr5HduUETln4zr7Sq2Ha2sbWq
JYY25ckrg0vKbSpIw4X/TuxZX6mR7UZJASOzqQ1RLaYarxoKrOCCnlFt6RXPRClUwNCWsEXv808U
9EABL2IC1KiGQ7z+kMUnsarlXRL1jEVBOX/5U3aFi9qaqUgFXA7lYYR9M7zjAd5jAWbN/wWf1mbL
SsO7aICKKENhWW73VS/3mZyqnCs62VI+auQNtn3PnSdeHfa14Ff16SnIxhUxRpaT07IFdIFK7dAW
8I54S3EA2bGIwBNjPSGkF98CZwNzm6rB3mCs6zjFV5gjPjX/yZywIkeEXXbVcoueJtBz1mYYvmPT
JugnkkWfar/3NxQKg2Q169jSPlVuMG/RaIHj3E3cGKNbVk9yMtZztlMyWgKb/rY/l6Fha6JN5evV
l3nT1fiHmUdJPXqMeOBYoBWV1xjCQYVLv4H1oKZn4/GVDKSgcdjmx2AvjRsIp0U+yAb1gDPmHfni
+ppgt0r/g02DKIMCZV2ma2Yuieggpfa0BsANHJS7tIVIj7cq+HOedwE2ZpZakW3/OedRwORj4E75
KZXgGoP301XlMSBGDdufHy3xDoIN7331Gq4+e0f4MugybOWk4+afepqBnqE1EUshn79ISxiyl8gk
QDmAGfqHPVg767c3NW1U9e+DjXrA7tvAArs2cwMGB5ZNYUj1ie3fPjYgQZZKqJQtuGyJjT4RYaMP
k8a624eqUpynqd15gMy45Csy2G2LXHD1cXYjkpe9bYpNQUg/oR4EPjauJPw3oZiyz+zdq4JeXvO1
ULO5HxiMk9xEd7I5qNPWU/K3wJpJcs2kyRJvaTmcsocpw3nkbkpH3Ty9oNEqD07DATN4n+9Im8wn
dErXeyzUT6hix2eJ5kt1zwXtxneTFkflxMaA9S1PSviFw6Rp98WvxpX5KGZwa3aVDzZoIhAwwHiC
QNwomCg08LcvP9zTcslWLKt2ugEBF0C0FAbA5Ubr7bm/LqK9+1budCkrJRN9FkM6Q/1z8YSdND0o
Ri10HS6MjczYJEN5Bx9EGsbh/YD5CnasvwF9yd+3n7OkZzHGC3Nl1zL7e+XWMwuA956Kw4bHJRB9
NhX/edYgbpbR87ZN8HicOOkcmWebGFx7LCCT1YkWZ5b31DLLUEkb4jhZVZ63hvCo9INNrHlacvzv
uw5BwCZtvKO2EFdKhVA/6Mcc7aSQWCLgDWcfSEWwSvrA6nOYzp1Ixu4WqVe0rcxg1/S3qJGRVoM2
AmRHF0gzivyCT6rUsBaHBRGGdMz8uQNfzXNwqI3OfXiKd71rZvwqd4btYaxXkiD9verxRT/MhVmm
xZ9IHo4OfpmpSDwpwcCTjyQcSj3/K1EOCwnSJmgBGEDzcQ48Ea05r/BE8RCOZXVjPiTefS5k/3f3
Ww9VoI551udq+Q4Lbww6G1ZkJVLImgRJ92xWSelF2xepTvh/JUg/Zx6Sc1MHegI1HCacB/+3R5Vf
v7P0lm5ecSbnfMtzMiGPef5+OxE1xIHKFUe3YALvU8RWn2ajLL3jfNcyGxDh/1gkPMon4qDsQXQ2
zooA05MjUBleBUF57n6QMM8Qi86YkvEjFsasQXGn+4ec50OywEEY1WB3t5QbRF0+Ulk1kE2Ne3je
atgGrxCwkRvrqYRs9k7gpJjxUqNWYjYmWGnaT9Sjxs+zw1wsOokpbG5cmhpXmcFpICFxeNKGCGUe
KnpwsovtoDe2qhP/QYXAIB/4gztxpPr2K96WBeYX7rPZDI+MP6iv33FTNcTbqad1GjQHv+bZOzk0
pPhKwqA+PIxFCVAlQejuntjLS6jhSeFPGzvBTEzTg/ErbNgyWvw8xlvX61AunQwICf+6Jh1ZBRbO
ZeHX5w4/zsKp4JE1aXYcxTpIRj+T1xHnrSyw3+N7+Dqp/xEiE3dNkEZc6R203QmbjOfV4SEdyeqC
LHjnP59lJn0ASMJNi1LWkj0QgYV9DJNJnHpQbNqSmWTDGn854UAUHPfh0SHlx9Jkl84y+irswCzq
9bCEbEcIGg1yNZIoIJhQSQoQgr2XMHeCG8GXjNpe9TtQDqQqWocYtWcYWcyuKTG9KTc3NFv0zCiT
CPC4CsdKMC+6PwYcQoDptV5ldF1FIMsKJwoy4SnB3+M5ipYJuZipdPezMELlQvMwWEo/SRBTIAei
RHtkcjlTrEb/MEgIwUY9dyYpQZND8rmhI8i+aa3cKC2Ls6xweZGpbTOkgXI8veeIeMcBLbWT/ZbK
YJ32DWTDA4+lJu09r2KPpsdqD4Ty14Lcp6FQki/hjP1Tix4mBnYUx5c2H0Bwc9LA2aCM1HTf/lpA
pH3soail3LVd003hW5PprSaMcsW497IVR2vrWr2d3HI3Yur7rIZTv8sfEYwWcy0iYncmsiqK3Agb
HjZXrPYoSot8WpaG/6d0lPkGGeAqtr3bs2DVgFkRr8XNssjaRv2aQ8WIDTQ8CC5Mz4bMFGlP85xZ
WiJ7bhIQ/rcNwZXzhZtqiEq8WGIaTTQMTCnQWiKaj+bc56Ylx2NBkT+AAGltqcrTviwJ6A+sj9ay
VpClRLbQnyLsRAQj8EBGcx8CnEezFaIrhGxwWo84w51JLjzWK5/VZ8sX988Pcux/aiLuynk33jHI
sErpS3R/u5zXeAl5cEEmqYeF3hx+hZXpTxZgdVrIM/HdFpQ2L1o4e+91NkH8EliRQ/HtA3oWZNqA
I6+w4mNPvfYXER92Agl0Y7Y9jYSC9KzhJ5sUBgFmrFo0oNA9GfOpNV7zrm2GG0oBBtGHUf63Ube7
x5+91QnLHAAJwGSYqV6Jh3rBCcR8VxBXwW+vJcaRCAE73KHLPhLUTkEW5ZzyvqG6JLV5g6Z1xR2L
U3xhoRHg0lVM2HKRBq/NOstUdVF0ezmFnmRRqPudKgIGKP3Gu0yVWFwco4vyt5YwptbbBbxXPIqc
irYM3EYZom3NXXFbeMKtXBG86UCUVJMecOC9xvRT8aWe2WJqXSp3RChiVNy3fCkWMvhQu26viksE
3SZp2BQYVThr+NQnSVISBSI7jtqGRWPnZM2+kUywsSY58ILsoG1tEKbtnPxGiQOeYFQqI4/DdR//
gnIAhWOk8eHUR+IhdG7dUR2OU/aaYqRi2eXQyBmiVe0FstKe3Kg5sJQqbE5xfXsexqWbKVFW2tAa
dQ1r5h7zaFEXlnI3vmSA0OFL8tnPNEPeOg3tOEl1gf5Qmj/GosKXIsx9YiclqEgMp/VmZicTGEgI
6So7kRCSV5QWNaZ+q/eMAzjQI9BnqMvgZ9unu8unhK7yEOsR78zJ6JJWpfvWZKWtbDUA/5HwAgE2
fkMF/qxbew/okpiHHM7vTyrBrQOFLB0aa4xMW8oeelH+gSUSJwQb9NeN6Q5SdJdLqh7PoDpRAkeX
JNOYA1LyOu8lY3sh8t9ZscZdGm1rYBkhAVErV9N9VPquD0ePWJakGmJropvrCIwLdTZcRGc7IlYN
R0RSwr5VGXfT63Hgcolupi2IztY2uumKuSuo0YSttGd3EZlI9DMFCHmMdItXiWineb1EOyYYlpNo
rwVYVA2FN/27ftizKzDTPQ5gpVfa3bk7dihoxSiY5nwOUILBN2vNlO/9uh6Obn124sMXSHgPiOyS
XxMF4PQZHnVrcoweYj5JakvtJDq6X9kCy9oVS0dXXJWcYO0azIMirLyC3MpGnsGIDmrQcXh2qD6/
vGG+hmWCZHKDfCW6VuxaQgb/xWrWanifE3I1iVigzzaAEB/HNMIcb40XKmGVhqKnEtF13drVulQ1
bWux4Ep3stU/rlVA9wu6JbgbzA2KehthPMjZWrCyZs2ExB9SbKSaK5QKzkU1B8bEUkHe7p894t9N
uzPFKBD5XJRAEp+senCrhmbbmWg8svklu75TtwQWokPGzVu7QQ2HJLzDPWxlhe4h8krFG+i3Z1Hm
37tSr8gHLKCMBMeGTspmDWwgoszA13inRgJ/yFNvGwM2LDXz+ID9svzLwu/8wWYLA3nE55UbLDXB
1vOOcK3k6sYo5o7UH/zgfs3/ScdY8QQz3JAf7RGoZSkKUKD52b2a8BhcZ/svnaKyP6Wp9dYNXCS9
XD93QQH0lyr3SVYfVB01xr4n1vPDf8ZMOOE8NQntBwg8RWWTcRBYEeTK2Bwt2Mv99T+Ppm32vkyc
eT+nFw5d33EWw3S5kxr73TwltAql73CbAJe9i4NR4EgVPk6RQ67M3gH1N07An07ZR6kk6N4XLiij
lV3FjnNyuXD+h7s2LrttyVxgmtdIolOyZyrNVzmLlIXe0NfzBcwePhbgVRpQ0Uq3GCQHyLXy5MdG
B4AR04h7GPzYrf1GbLwFnlPb9FGy5O1Y84Fuap4g2UGvQC4APEcVofbnwRHxy2GF+Qome5moBPAi
Jrj8LlZ5JuNmnpMaAZs+r2uB2m+USS3ypHhEWpsSy6EvsDqbmCgcb8lX9l7N5vEQ8b6oEWGeFPCV
vQV0xyX/TRdzzu9n6HqienvQBepUQ4X7ktZqJjLPMj4nD2AEysnLc56oeWqdobUSx6t91i7Z32bq
kt2g3vLwdg0lwpZXkscrheIQaJs0K1HJNzzxWSajRRf/KjSKRyvibvulRvFNs04q7Et/qpELM2E8
LwpheysZ8e/UEoqC3Unp+s2LHn2Stutlt4GuD8Jdw9VhFCraZ4NfAsQh1weiU/Ypbrxs1H6a1Wze
mH8oPD5i/Zcy6FPzvIFtdml+1/9mAReG1CebB0i0vMDZv2Ti5NEl5r5kvlE0QfGzuuRZ+Er2rY4e
7SDm2A6hgGKoiDd6YNnJMp/g85XA92qpmahSGJSftu7pKwCmjIMOZEYjFr2/irM5TRp1Y8T1tHxc
2deCrXb9ntthQvkKRoodqQSOiqlqoh58lVWY9vAJtuy7F9YUUx7GUZHz8VSabPa1ibxZoImD2D9Y
F17V7kj5wGALg0oWqmLj0MtRjAgVKmCxtVEEP9PpbR4NA/uEcWngC8Zn1qTFIMbXwKD0LVeqOuWz
UerMf9yFpzUh9MZhcjheUa1whl0d42+W7DC3WgfjuudSdkE8JG/yiPddsh4p9p8wujKoAqZKX0LG
ahXa+/LW082Db412Co4w75WrFqt3tpqCHlG18GkEc62EboDagauUW7BxP1+ypH8N55P6erg9jSOU
ktwzzJv4M1yi/rwmoCapxBDNALiJGTe01kXdefyHnyAGZjK610rktqGIwDlXU+4tPYbJ9nX+mDAb
UIM7DIqxx0McrR871R9dZ9yYn6IjXOTe/Gln7r5NOUh1NFJ70weG3e83bPfrYSSMxOA2fqLrmR8H
X9tY6UxhExze4ZWskMq+URWpaZUTVAdaROWUcoLQCd+ytGi6+FVALu6IZDQ1O3/Y2tL4TG37WvTV
ImwXYMyNJkRRsER/jdSY/ERhBvLFCqjoCvTXV4Bu8IyFLWOpdW0FxypuS4T0Tp2iN9TB4k1zZDku
Pr77n50CLwvMGTHLcZK+tAfB1VJN7O2VPZLWTs0OOvHUk7ScrorduTBQFzpW/vj4sPpDobBv2G9D
Un+9ojobyo8EWsZtldh2CZyA5AoPQBDtpHeZlZ0pdgpJDKYDHVLm9DkMCd/64cFmpdW+E8j1NY7G
8kj/5H7oCvqzzGEdMOjy3AaxGSqvgpEiVkvxh/np4U2j19vTsCsseb5L6E60Tl7fRuR2k0Wgcr+C
EN5uJmP0/pCmg1vQ3USiwlU/d3GU6mp4VvL7OQkM3Ak8g2kUAl847guhBpkZ2WVAPbHPnKE8irht
CHqJfpICcbKAltsG1hryMANrtoiDTRZhU1b9iO/dVR24LgrI2jlNcUINBxVgd6cRORpT6ZQgK1HE
LdwwFLJpQIXqCZHA61arjdI4x9KuAdsFWYz3Ow3okZAX8lkD+RrmShHDVqa4XBN7s/l8Bf09MgKq
0Ow8K72R1/bM5iuCzhQcpmlME74/R+zGNoMrV3goE67hIX8FZmvI8d3NHd5PMCyYrjyl6FVGgcSI
AUQMJTzYhNDzIdCaIlVnPbq9XUOOZ9FaxnqskAiQK1rSPc/hGYlUk4VRmbwg+TOYuZ8nfYuBD688
JhA+nFXcrC4BEjlzD6xaI8UUm9x5LQCKecpnRyX5PgWFOfIj4lbxsYG/d5BL/rvPahYl/gCPwfwu
9ULUGPfplJy5iW+OpftLWpyyFETnj9GDxXdqvdjtGGplPQ7D08yNIdxqcf3jqe65sdBKYM8dS4iU
2OOYmQkWB7Cg8odn91d/l4sErOCN08NtkQMCxeZyeZ5we/3v/diBObWlKNX/MBeSZ51T6gEoeBWi
oQzoJ84lEf9qnplRlfFp+lce4JcdZzx5DWcM85I3chWqU91ff8QB/la5nqS7fJY88FqS9ZitIeHM
uyZBFUx+y0s2Bsmhopy0suOwEoYdaG0s0fBjfCLrgWZd4ysub508nmHxZr7vdl9iw/L44Z7uw1Q5
qcS14Y7mDNcMr6dQ8ZUU/IfczPyBmDMGkek7MsWl/w17Bfo5czPjwy0M6WbpTJTYLel/l8/ofPhw
7UVzwP3P6ix9D1p5pLmidn+qQZ6O8tAP2NuJ1lXr3Yr37m5cNzaHR184aj24eAvzo6Is0VADDMh2
bOV+EK8na628BID2kXJ+6q1bJO3/ynHjaB3iss+eztkxpT/O8QG9lLYguRN6EkdihrE5qPEgoNNx
qss+gTggE4GjBJURhXTGR1WVlycBqf2pbnukTKPI/b/socbjo5wB4ks8RJFW/CSJ2CcQSrLDAKQA
7gLwRbRSohh+v+B4BJLYlVibajPhc045/q6BSITtu8BqtLzRgMQKPXWJVa+UQbcFYlG2KoNyL7GN
/cVDHLe6r2g5JpC2EHddQH1VtILEtAKFEwjFS+Jt9p404P6MbcJUBuiZe4DoZD1XK2hXcuQXD0BK
N0s6jPdBvVM37/Sr7EOhzkz1HblBrtT+Q+S+OuAVC6J0YzjQOT9wawQs02Gs6EWYGlTLAKpTOqWk
3UA5UjOHcnJpJz4tB4/pLXt2ZrnhBWkjS4fsbFkFmnOYeX8PnMNTtVvh+wLwnYdYEAvZ8f3W2lqv
blpbnLZHCCKCQtYQW19K7XHbRFvfBKgPkmcPLsDdlHFVe7Xf5I3gw3bU1iS95RZcs6QGyCYsjjUF
3l9b49uHaeFAkJjoW4eDsY0py7q9WwFHYfbecfmh4rQ9QPzYjKV+gUN0TWcnoaYfo0M8lCgqhGFq
yftakXq8un6ZwVIjRXTYFB1Oc91PseugmirYO95jOYwu+ZCG93W2QZctlTFGhFDMNc5XYdmzRc6f
Ebo/n7AuHrBiMHsLHRHoCixW1ibEVCfkM7TzeI7Uoa1Ygmvun1bXeaAa8ZEudVtWS4+18TF028G4
HSPdIRv9ELaBmmbSowKVPVSOYg6frtiGiFcE/MyxBRf3q5a9i0hVTufHkfz4UiEkUSNhs1F9//CP
qW0MEAUPfqhKyR7Cw8XRPlCViuRluD1FixFTxnnpl3sE/e9NvLXLu8PHwAZQocYO++JvrIsEvIAU
U/bPw2q823MDlgBlZCPSB5wMy8cuPJIoA8U/sAV8i7cthBQVMXDv3WFrXMQ41f41/+psFtMl9Umo
JWgYReRtD64VEOESP4YZm+Ere3sovcnu2acO0SmpWZ1FG6+jrzlztXobG9QctJWZG4VcboNkBqWG
09lX5QsK3PwFowaNsTfJxSst+O3PB7W49GDI2sd8wMxTzNxDb1azRO4hDKDiBbqlMQuiGyeyo0zO
/CQ755np43FESgmZ1Fgkojrmujz51TtuoKdCegEOeKAn4ZQohlfu9bV/kPxq6/82twws4SkdBCbj
Jac2tH1JqHxVhBnfNjLqohsa4TMgMpa3CdQXuNyP+y8dpKtomOhmxLvgK1BHxAA3s9daf7k449na
ANQNMt5m3B1kjdiJjgRy72cT1ePV1PGNY0Mi6cp3WDtoaObvXpJV6kPFgqfqQ8IRNQeKOS50GrTn
7XfT7+nmOfGrW+TtRK18pQL9Bq2dKk+OxxDXiQ0CtnfpwTnCRo5hPT5pGtwIJC0J1zgAKkKSpYZJ
1t6wF4Sf5F4DKjvx62E+z0+3kKEInAgbfh5/SwPKz1T1UEnod38AD6IGNP5JTgp3SX58FIs4xCJE
LinAu6AY+u5SpVyNGGanQuzPqN5FtqiiuRLHCRjwR9RtspxoseNJvcgiGfDYQk6akK71YWRZFJW5
2nMAHReIEZnOCN8neYnIVZoWT9+4W+ruMq4jqk/5lxG7cpEvTriMH27PBXEjIYWQDuyHYTnZNNqn
q/Itx2bINezH5760dHk/g/VGTgLG2eOjIFkioHgn6B6cStSWwXtxODlvmcfLIDKNUKbPLQ3CZNMG
rSnZFUiPTKNx0E78RMUQvlpX71u3XFngp/N/xa3U3adD0i/36MKeQ325yG83sj/44Dr4Z4kjm/44
ziiZY6YrdjDYRoeaWbqpeRkakIUslLQGmmo/6LYAmuwwW3jhxeKEiDpa2ZVH8+2J/ttArurK/0Mj
Tz1bHz+QxOwcwqp95MUcBxVhRzs1xSU8PRiNUD+rfgFNSBZHxWqUi57S3CWsUZW+sC+TVMx2IgC5
44kBN4ctW344zBdbCde9ZTNE5W7A6ms1bvY2R/kA2+HtN9iemwzhM/LebCey9Yeh5OOj4TD9V/LD
hN3RVsTC2Aot6YadS6/0fjbrN7kmCIv1wlNQVR3LU6ZPywyMmXCdkTNufgeosSDQCaimdG+GX5++
FE+WKHalb04DRJOI/NDjCFWVF8M92GM8RFUwFVlqNq4YPn54s8bsNenQfa/UfVNcPk7JGJ4/aZVo
mzkCQSYWITi85ogSnI4ojl5uYedQ+wqX/bKsvTsDwvou5GtOb3w67MqD+1ApkzxmCJdfWaFOjsgO
qy02OIiZEhG8ilLh95mkCJSj37cvoIwnKt/Bi8q60zdiO6/JmKFtOQ92xrQqYqWR2abVAJo8cu5t
qW/jrw5IZPS6yAWjVkhM0iqxivhN6bO0/kDou4EWUR/WtyMboqPtso4yeVE2G7+ys0hnoADp0bod
xs13vRIMJVvKu2+GsX+om+oqaVa15oyXKNE++65ibED+pWgnxXcL7rIgko7LZrM1HSGp2xMQgLZE
ZKA84C0BqX2hDl+40FhHv7qi8fMYHN8l57ADEz47iVskWdMTCmMBfD0lMcMFWhpCnQJvc2jBG8vn
0GdcejTQ3TNjx0sAY5isEbsQ7B5ETQAtH6kd2KlGBsJiSgubhzBzal0E6LmpuML2SrSE433aYWpq
I0TVfYSnZtg3K0lzkblE8MExy5rqfcgW/5YAUmbw2Nq2zMq3kyPsfWr4PNdIojR2fesIaax3LxmZ
cbsrhmHe4vbDRydY6XdPbk5Se6vz5mILb/sxYblKSyk5SHYbW/MIYTbvZqPDEVGoGZd3f9sEtKnM
LGXzsf5CiILjJE9oa32P5kim4CrUorUIHBktWAkkPJOFkh6YU2qmXe6LwXCifQd4fChTOk8z+uK3
LvSG7+k3kahZS6TC97QcWWDMLCVTWS7Nh6Z5LSoYITeWFoZxmHcq3ghMzdspLHhaz1vNhQJQoFyD
NnKJRN+uKl8LHXONMZkSYYVjY/B4vpUJSEp4/5bA1kbgp3sSxqfib4G+XMP8GnRmpOfyhIV0Inr5
IIC3z6V/TlcD60saMbrVnD+LjrOn+eyeDq31PRSwMnmua/NXcLufFi2ZFbnZDH9oZpr7LOjn9UVz
pOY7pDJBY7kXzq9dvEb/T9gBudnLsTJF+FRYGA/PurkgttVkoebK0am+8uzG5MTPSbtBE8PcNPVj
SWcMY102f43mvNYCaEN0w56QQSUenj1mQ9XuH6KsPMe0Czv26zVdY4tPyJdbWDuoc5Bqeiegt1Uf
q1Sl4hnYUxoxgiG58lpNw9AbvKeqNQs12iXWxLdhWQQYbU8fAvXUgYxKAeFnN5dR5xNxBzfUwL/+
I83jQyktiXoyfgIVkwhgwGIlnVukxySfqbg/pbUPMEczrzLUfprIKdyF7w+pI3GrACUOozc7T7eB
l3umhRY7Jsk29igSoAFcccs1NjIE2yqL/H67XlmxlU/xUv9/Qr5btQDv7/B7dxFAOqIYcOeCC81U
TxxjgEZm+y2UzcocnDvxrpbxu0HxHsNzSzqYGbtg4/2GMAbuP7aJU+7mNRLbX24UT4VkBHZVxWTC
xRJlmAYyj9hkRIuYLr0+BtdyI/beU0gXgBeDBrEYJUeNE2maWFYZToyuGDdCS2ytBgoVBUUc5v2m
qhGElR6/tg+ed7W22pNwNL1dUDjAY/SYUgBchFO8wmkt+auW0+HVo3k8iRhhyeo+5Tx13AOhp+0z
WAQUtDroGAEzPF5Du8T3Bfv0wbE/6K2QjkAcgI1nAoOYSUOySSiq6kyTazIhVFxldxA+/H3Z1f81
X3eGmlZ5tR8q6ucKJMc9E5DPeefvyFshP/+bz3mVllRIchWQtTVpOcYQAXHf3s6XUyMXjtk14IAY
PSBGeym82OWTq9j3jaRhAEgiDnJko1jgOaSD5IdkXEOiudxrRfDMonN+aCIkyy2tLhTEPyEqn6xb
BdpfbPELFNXR4DDJXcqWykjGly+9qhaT0hLhLFvwqPXShk81bUAez3g78TA803iFgKZkJxivn+We
axqes8fYmGkggxWQtpwOvGlBSDzJM0h66HXaPay72W37u0gojDkNauIpvj3KvogGICZ4T24M8c8o
mUbdOIimP9ycTuuy1yi0tmZmvGdZYnGm5XZmmYZaGokSyDmaRxjmAgjymx/GqQQ+ZFMjzxO4yChT
DT29aBeh2GNtq9Jt6CfzZ7q/4A3bytPYAm51H5hvRRI0HE+MbG4Od7nkC+vbl9qJ/DEay/H24RgG
FVHoiFT0Tm1wZmVet0Q1nrJ7EmcfzudDp+szW3KpxolztEEIsXzf+XvZDrviDiXJpnHv/nnkjLGP
rOLcOwLssqS9ktdncTWjtVskK5PnTJR1WpVgkGx4kRFWdxLOLg7iM1V8PP7s2n+FPBoBQT7K6NtH
qYS24+FqO/ljDXPH4F3QtQaeSIUD25TiZFxYEFXYRgs/y8QnT9tmOGlrFtsCtJvEa41uBdfOYC9u
JRys+pFkwIj+EcIg3IouB7Gy+ilXLJhDtfkvQ1nZb7XYWClNGB5AxAqA/JEShjfUZShwQlrdhooK
86obe02D6ugEFUIVjBG3N2ZWo4RKsn4T/pbsFXr8WTogPoiBWZ4ws7NxblJYka+LgzWNog6kLv7u
8yMJqded66FlRvKPKvCKJ1zG5Q/473ubU/nzbXwvD8HvKPn17n60mR4u5RiHihPxQxLcmEgepbcV
069SabY/PllCn8zLezTorecUzuk6COfKwww15FC2b9Ob8QxMyilpk1eAHRQErJs9AXJZQPJmifbY
//sO8hLcOgc6rTglW6vCWFAZAD0FEw/sKc5Og5/2W4WMDmTXdF8rAWmK7//GsIHLFZMYis3tIYFz
Z8AsFfb1TeuJ1ZGqYlhMOAGMjIu2twGHLo2wBijjheKGlIyE/qDN6m2OUVj5iXuNR9kPfjZ72Dx6
5dTYV/rBmNqrdTQpel/IxKAhidMJuFwSw1HEym5vBHDwARzjsjZziPq2AE74OLT5rzb0ojadvp0o
KvcVKerzsIoBDmjLMfLaBDmk200gGRsry/qhTvPTqKhTR2q9dk92tz+A4sFhjbv7Gaj5AxS1vhPT
R+gqAc5l8XyHiIT+GxAMf/OSTkia5kO2U/jKFDIuAV71zHJop3Kxl+FOd+hUd/uBjhPjL1C0kqjX
2fFTRPSB239b9JTgCX70TBm+SE6I6bW9aVnGUUg1nipAsuvrZ/C24QbomR/JRRfQ/r9hYZZXEUUS
QZ/fscf0k+vqHJyhk7rTgdBbsYsjh8u/+b79Z2QONfWgFIs17rMJWxibBL03Z++2FJ3GYJtVc8Hq
/kw1BzYFCdmnF2R3apYVRElototI/Ky6Hr6WwmemHbXZ06penOvRJOdImmYvfNG/Dg0kIBlFx4ia
9exXahwZdd49325JwjTJeFOzBeowfjLhGuDr205Rqiy7PU8adcA/O7bX+x4GKwMzfTVwREsRhFTy
+FJkyTrF9z+nxHvmy0l0V2Fk5B8ZFtw3NVIvqE1y0De+mbujD1syVBgvMLnMNfK86Z/Av9NeLkdu
IVJpE0k1QXFJEIB5KnAa5s+wU/aPdT6vpTcElt/pGkp5wS1ErOTrwsJ5yat67zAkcD0vdsV6GjB3
zd78/xyBAfJx+YBlaCvxhWA2B+qM1m7gPPCwquB99DBIKHycP6UAMWX2cBMxyEX3DM43twJckTRl
bBNFeB9Vc7S1/YmcT4jlby3O9tvgw5TItivVvwVL4Z7sJT69Qo2LLtY8eyz7tffwdI5BAY5I31sB
zwfVx/KR8X+uI8sZCM2L9b/EVBlr/D3TB/YmK874N2RwA/Jewz8R3Rs43c3Yufal7fvWlqk6b4Nc
2hIyPUN+zPDAMdWw+hRVELs22oMeEKEhu++4te7c1Ljy7kg6zaULznr76Cdn1Eh+YygsuPFlDnG2
zkBjkl/96Xi2+HL7VM2GTegH9AHKqK3SPpeSmz1FG5XdGF5Ljzz8SXz2faVH5gbok0TDRuNjwpKV
R1r7/R1niKHwXlaQtvx5spzXoNcWzti8GbBSEKBWS0BTV6Qqw5a3zfKb5A7iKgGGBniuY+FLL/Hg
L5eCyHqL4KngkI180Jw0r3KVBFBHV79Xn0x2RBCU0AM/EPzdNEIEUSxP2QCtyywQCpsFe+iDIWx/
P+nAjIRatbTox6Fg7UG89d4zxwC3uDKhvIhoPFCEtIEbS+Rpreh5EGtW5nMGXo2h4bnVwDzAAtVr
VJXsYibJRA7Jw1gnVgpEvQBzsa3XMDFqeiyijtjiUZoMRMW6d6m921g1b61eiXeSAq+uBzZ/iKzL
zBefRqS0ZVpqG1cqRJhsoMarsA04R+imc5rKr1bhbud4bUMnmWqUnil0fcDYHWIgS0GywLc1HSi7
ciG6j2k+d8gmJZwKEDSIBrUM3LE9pufqq+fvWVubLIoIA/L5f35aQ7LkGFrNWpSTZznpiNIwajTe
lg+ba6Fosiwm8cuMY/Aw8YwSkBa1bBJEmqikdMEKcPlHiAB9APRJ9AsQARRcKe6UYJv0ghpLC+KD
x3V77VFhm/QysD3Bh0hLozZ/2pQJ/BgW6A3jEmHjdrqCWZID9013heS2X5MAKAtqN6NUbUBnXRJb
Zf24kxIww9OqXTv9W6Rr0bLyZPKqmIQ82WSg+cUj8NU76nlArvMWOpIT2B3J75yXJfb9dp0dduJr
3qIfgTPP5F9b7QFfqrr9b1a9SyU86XcYoS38mlNAOkj7Yk18E7lhasG0lDe/CkwR6eAjVQu35NBg
4FLf0cccAaxWgH763VOFMQB8P7g2CAXxsfSRWO3DTc4aqSGQdZL1NcrWnl10THJeqlwo8SliV2Cg
07YI+mWUOyIexBNXQJOz1US0pM/ynLZJvVwwj8S30zdXkkp+wSEvVvitpW5hlxiFveBBN0uUiiQz
fX8cYWn/jxtMamxdKV9dNR/DGmGM1pbFRRY4SxkBjNcFIYBE4s5/oe+3uvpjhXOBjJgmLt2Tyu+P
eczL+7/dOgo3tu3oobTPE1Re9xw3Wtd1HC1Uldf2Wnqje6vuG0QrzBXayo4eh4J+yougdV0tFPIm
cgsny8tHIejXMy8GUaMM8csUuY1LPWL7Ln7BCyX8hnUfEXFfo/m4a9acrVOqBFrhH8pRfeCucDjg
BF2n8mjjmOeLu9/yu38S6bnXYsrIbVCbI1gnoHC6ImjG38r+D+C21YB4n95crzsBg+mmsdO1QAi5
bVX/yBmpstfu0p/uATSX1BZt7qsDMWMJJ06xJkFFPGj2ogMaKqeSE7skV/NhDXwwWFom/Uidex6W
d8xP9npzEtL6PmhKa3xZh910caiM98EHu2Zvb2oNSSuGcZENCIq3qwqdEi5PewQTz0cZMQKXhD6w
SKtBqd9RS+24C5F7reaVwfA2iH9sU90EbFDp9smfuxDoGyg1Z1Ws5tFOBPsZ3+WdjkH+t/o435CK
jFiLERbr1LC4zDQOXKmbUDBrQvlYHrI3IViWUrNSIA89qSczcVvGIkdd8MV8UOkt6HF8a+383K0N
RehA1XLue5SrHKChex3xYeXNwud+tKjUANuRPtDn1rU6u9P/PViiUK+BriOJqLb18v5EGNBJ+3+x
Epi3XizG1V3abv67VGefs1K9iaivKlgqy8IVG73df8aQwsdqzUzuWkoOH0hkr/ycwxksntUCjJMz
DkTqdgCMnLUfEUJtt3uEbgc9CUvlvAI1OUwjPipOpQn5oHSnG2xALanRrpJo28eJeFiP42zjWTOD
Yvuwzo6MIv+EI89JpOzSfHCg2S59A4HcRGmEEW6TySQprnf01vkpAS4WXKF1WNJnaNpgo2FGcyjl
4encfCDjQfZBqFz9Qmj9QTlaFyZ51YYrswrDCY5Tv6K0gGeCeW7BBfWqys4nshgin+zqhOpLnQAO
QJXtRRX7RIDTWX06aMJ41tl+9fxt9DKRRE5IZ7Uvd/J46Q2YbnLncVzXYjFfjXq+atM36NlF1DZ4
aV/g8o5fO0RhW2FLHDDtHPAVkZ0wbSn+ZoIiib6HW2vvKlG7/ObCCu7YZhmCFXQO9ki1Sw6iUg6z
vXvmSyjF7qxVofKVZ8oZRFJ2Kpaikmd6f//8EN++dMQiGaLQ4xhQJ+D2h6USeWUwWcrcBdNorXrD
rTaJEHiT7szduZ6wknoljAS+6uw+O2sYWWX8q8lWlY3S3f6zrivD7hslRDa9N0FY+M+YC1NV+8JT
mO9JTfdnv2Vh89O5CTBSX0ZDrTWeL0DZvIXE+n0TAuGBUQ+GUwtE5XevO+Fnnt6weAydAdKksLSG
2yp8RLpxoeeXONL4hXl85hrdngIyEo4+rwOU1ejwxxERCAQuJybMcVSXA5dXOu2cbMl+Cji3n6xy
gw1u7qb9QsF3o68RIergSkM3UMn7IdLSVdU2vG/v0QlBNnNmCempCeVRAe5GkzQ3lMoAbZlvWvzn
ig0QPEHzZdHWAkBsyrAfCkAeGtLEMkyac31eKPCT6mcgHbzBLKUqrIQLFNuTbslvD8SxnNjSgQ/4
2XiNaGzGVT7AOZVRJH35IOilS5zD0vt1Ejq3viscZkS0mDVzJ3oI3sEtpicISWKwevH6SCSImyl4
0SKDH1NtokCAxs/9GR/TzHR8UxRxjVs6kAri2x4trONihOcDddhEjJQNEt+mnRceXcXPWOMoEQl0
e4TSOoP/RhcVI2hZBZfHtQ7OdIyjIYZCsOvK6PACcHAMBtNEV78vSARkJbYqqR9zVjTR74DQMFiv
9HQwoixRttM0crJ7YdJ1Fp5ssJD9UZ4P7Ejj0u/0KzzlwvwIi8m/3Tydu/k7F/ep7lVV+6a0XRiL
ueGPVSWEpMC7RlJuu9qX2jGmcA9ajSX1kQ2K+wxSFHn2bVBjtp5TKaGanGMZFGqk5MRfXnl2XDhn
ErRX+FqtCPshJyNJVtqo74sgTAhzq0kTfNZPSQNXtsClvl2gOcTB5g2/kzaueWAA32V1HfL13cLR
Stro/8//u/tuqku4mcqWiL3mxOepDqKfEHusJEN9hdV4UtzHnUQyGsDgdQzdzNHFRkr8gYJyA8hq
cZlSz8GiA94dcTaDsfDFRWlKt0uYr+Y+WyCN0UELb/68hOB0+QXiU1M30Fk0Svutk6ErywjflTRv
TvMXFK5g2KWF2pX9u2AhIAuVxJ+5d7BGr42wO9319iV/iwnI8HuKUAvVuLu5M+0dZo8FQ2wpvPkv
mdrdYtXQgyzdG4+Xi4T85ojsHlETJmaHQeinFcUcaEUDj/9+1Jvz8PTupM0EYPg/FKkxE4w7/KAd
ENdXBawxzgEsr7AjBV3f3XcCZ7+21yP4kwv9FbHN2rRr3GNzrf82/yPfTojOZ22jLgbwG3l09eYM
6cSz0Faxpplo9KnclsljinaAp1RmwsWVGUHxnNmaqpkjrU51k0PzkFsl3T2l4VyW/ejE+pkRDDUR
PTZjAyrC3SoX08yoFNPl/HcLcGPtYLd7+TVLfBjHyD55BRrdCqQ+FMlH7GkJ9v1bgLFWM2v00FrN
nVnJxEwc9hQ2VgDrrhFTkumdHCmDjsGjYLXJT6nt82k0dtWJTH/MlwusT1p/0wdAzs2CX5x1pXqS
Cw0PjI9C+m29iyUVklFiTsX8ewB9eVCF+Zxzkhd+I3ARtChGpka7PDgXZh3BFD9uqGtj5LGjlYwI
orb5JPKKbyQgwbsD8mfifMYkqLu34pYL3e0SETqDft2czFGWwLlZAxTdxR9QAUddzEZ+CpZctooV
uCHGWLXvc02LjblMa5EEfF4ZYB9jO8yfC0cXBWEicvoHcpbA2+XnFSqLkoeucKCznt0jSGGBp44f
b1nXNL0pLCnzEk/6eUIK2nSri7mmsLbuKbQlX4HBkzCDwonaSK5UdFh2i0qijVzHqq7fUw+NJkGw
6k/ifzfNxNkzstrmdSYIQ4y+7+Icex4WrfKXnMvGFjgFPcxtpZNzeRGM4E3tyq9OfkYpNGfJMijL
JIIZr5qFzmysfDwPwFj0XmqyOzqT5MCA58BR1do4pWuJ9OCQJ89pXnKYrwi2aj9a/S6n5ZntTESj
xxhwE70v79vEKgKOkTZ1JrVNLmdKDFuEAeEuIZFwdD6eH5Bv+ccm83zWrhiOxgXQIGAXXC+VOdGm
3os7sShdrCNjQEIYCF2khhTk9cBhrfJ1gaw9j5WRhBVvk5IKeNzsBsdt7r/HmdI3RWnTQ9/RBOAQ
/4937I/7Fb1kMWlEMA/PiyqETZ+lpR7fRYj64FmfxOOxZ0wMDSMBr4WJTCbaHcB0P+DQfUbm4mxB
2IhlFeeeBPU77fkd5bcnDHcZ1zhOk1YbcVIotc3DMfu76N15iJVMqVEhV7eq0MyDbh/VitGx7vd+
1SQLK4f4JT39ZNZ538sNTVjXIFmSbgVxPGdKovgwy0qDHVGrLjBfcEkfsAqqdyjsJnT+q0hQ8aBE
6IEXrpAxH5vQYIAHF80sZINaE3G7DfCdUW0SBAK6HYn26ekXJFi010vzaQKiiUDMeMkDlAFlTg5o
aSoKlGn/KoFfJPbMMcDF51E4xEQLMPlTnhjkkMw+ZYxwSZw40UsV87zYjk9akAdVfo0rl6h5CLhF
dpCZM729JFW6FvWWjfjp5knpuhsey4OZuPmFwBgmaYJLU1fp/UvHaXHExmXx9VA3esGAXHrmipyC
g1Z03iVpRan6G632ZaFZHvi/JjabYybEckAPzSD8rH5NoxXHpo/gS5uGq6RTZKCK67EKEWUlgAos
ndx9HKVU2htVmupaL0avo2iY+6izw5ZEva87F6st5lGdkbsRYWY9yUescuIAh6cSYJ9J93Jvk9wz
1nK+gmkE3EztKqCMJsPXojvS2pQgJg9sohRu6Iq56u/6NMRcvD3rDDrFsvvL5eFF7qlMluIcO/fR
q6mSzU3gM2B28VRoNBTXas1+7p2Un3iYqohaC4OyADcSbSkPOluLIq3qub4wrXY5c0iu682Ta7Lr
dtj5VbegsfLQ/grM9hj2PqtbN3RblRIoCb1EcVsW1tdPamwkowZhboiZp68smtVx3axcdFP0k5hx
br2/z8GG0rkGYCZpnJpZDdXt30cx0xzh2/cJmOeQD8ij+jU+MTqmAAAvKr7oWo0fK3lOAHcVLm6F
ab8vMAz7SphIURmuzj8spZ5DWefDcw67rdakchRqswwy1bzzAvdz9HFsws/3H1VnjazWCirzVArf
+5qjNtqNcFCNclGhO08LqfX39GoFZiepdAl/LXTEddQEs7Zxa9nxHa/iA6hUFlWU0P1D4vtR0HdT
FcS8AL/TBb/aSh81VPOrLgeJZDgtJeme6k/vPKXD+w/LwgIj9KC0HTC0HHGSVLj2IFVCXJmENZjW
z0QhCVuzFOgGu176UrMR+QjUsNA28+MMRAtnS3zBLtvatbbEULcCfRrA5ZPbBlFZtPmlCPYJaKIg
oN4/aUNPpbENzff0h6/p8aeIKliTT9GNupg3B1ejf8wC+AsDXUQAszeu/8bZSljQaULXCSGf/N+D
N7Axz438xwfAPiKK0FnKQ/RvK3uEypLw3tz2xNaAMGdwQDz0rn+50E06EjKHSTIKE5MgRJLpplXH
QXrwKON3DATZ6CMY5aVMMllgSYWo6D5CndUq+S+KuR//oLLIyEMqFRIkVnzIKc/yKSDrtUdAA4N4
zIehJz8OSiz0G0P3rS/nPsZ2rWoK/Ua/llj3lXz6nwlW56W3DamkcHdvv+CFQxHjMuYABtD6J/38
4Gg1SYP+M2o+cU6ne/NKXwU6duKpkcdCGrcVnU9OcY1mvccvfyWaAQ775hOMBo1G2T4geBw45f6F
jex9aawuWwFLMiguAwSjISZwBBlfOImzO8oGMwbbwr+cNatGVlRo9OArRwh4f1QVZgZeYhslzAoG
niJkhmzo1DhtGntV69HtkxitoULy6eJTDUL/Yak4Nt05WpiAp0zq19Ro5ijtT6gZfk2Ku+LX96Ol
DJq00ZerHhCj0MkZ5MPFBvDyY9U2mLLnAp/ySm6heFqNxvbqEUiABzkv8y3T9p6lCa3Kdu9UBAjG
a+66zpZp1ZiAYdlMCW0yJINRxch9vojdNlA+IlHOaKXZwaE6AgkZVLKdwVmsyKxYWSQ/VrAPUiPw
VAc5cw4hAGWviYkvRLfV/Sy0YbKiUufn2i704/nWxg0j58tkmcih/y80PqVf6otXryB3XxCAnNAQ
wWUYlG0Gp5sJgrFPPpgd2OyYLX9/1yClh74o9k2KdSCw00r4K1lbIWFR6vgOHUiH30pxMof4+uF8
gaeiiJzr4DwgX0vE38n/dsHnNy0WVdPcAMlQLahDnydfWfoLvoFDbHLvOBEtTStob/yNN4MP3bWu
qUBr0YsaSVnKTIyMBts1eqkRVfIMaVdgr9ER2kEMb+sqvd0ywvkoIcWIn7sQBge47tMTYVCCxt9C
oAxJbmqIGUCfKt2jqxnmX0aK3Mlek+hx4dp9woEyx/EHSFxvKhXs6A0RVE/LZ80XM/eHuvt+JTBa
yC2BpbmU2JbzqyI+kECa+MIVI3/7TY/VbBFjP2anX21+WKsZZhr20pU6A0pIJiT7lzRaQHoeD005
2OJGFLbq9ISGzCtT1g3eQWkbIoyPJA3eDVKTYRwH2wyCfRJGv9j/n6GSM2so1mVOeR+TsOhdYOI0
RtOBjmLP3D0I6bxNLJOfd3t7MOOaM0ZD+X4va2PAQ+qAhbPXnfK3rQLTspmrisZ17rkeybauR1rm
Qza0cc5EUkrCOjfzPiuuiZvUjtKIxeTeZUP5Kek5/jdeP42kVP3SOPUZYuRS2baGBKppgoD59gQt
qXNgvglRC9oELtCcEsmDo0/ZdTLbSdo58oSTxpM35dnjcNNI7HQ7wmZNDQEIrUnoJZoGHQDvjB6z
NzHGw9YrTTRr6AkhNSzoXaZcJGVZXnsLb+fzi5gZAy53w7oFoXKnv/P5rdorPVxPTS6+VG5Zj5ID
4jQBKV955jaZFUkDmGL2mdGBxmzPSIIu4DUwECIEfH5IqCr+MqouTP95KXhevDZdr6swefjpaY6C
WxjACvJ7SNc4aFee6KZ9WhT9YKJY5JSwgw14pTE7ZXeJ2McrolVhFeFSYSKapiDU2UlWCOhWtsY9
6JQDxYfNOSgygDcvdbYbcxWpvSqo5ejmsbp0mD+MD8zS2Fh/L1nn+BeJN5NswRDYky6Bm+OAZt5I
bd/zW1qkQ+W1l6J1aHIVslcQ5L5Cm7NZ0OlWzZ9ffXV3rUkCOOPASZkLjYB0/se2/HEgrBfteVz+
uh32SXWY5fcFnSlkrDdRSnKHh6czKZfp1+1AXM5MSgbDNYUZFWRD24tvhWV5rW3vnfPnw4YxhDZJ
kc3CdcmTgEawqZeCI5K+H76JveBMSBamGJTmV+kLAlMyufMt+QwcfD3HRbZu5q1VMmWphFDh771q
mPRx56ACB34lqwSHB5Jaq5jiwWXgsnMDiIWtK2j2O3qtdw/3uoroo22koDbepR+h3wBxvHaZ2YC+
vQWxjwIwDwudYJdny/pFuCR/KqzBIH7jSerlnWQU4Wt7GGrEiaAa61v/rvktkfQ99Wt2JeVPUq72
Zi3i0UoBj0vYD1QliDulEvtJulp74D2+MuHh3MY2q6HaRPvdvyex/Ej6Mxp92BeFL09rLX43AqcP
Z/cHv387E6A0BrJU0Gz7hgs3j+0wkPpHD7eYYmSNGJilAak3Pm2UzxFtLXO/042gTNZh8r1GP7vO
ewt2cqGjO6Bw7/vnCFRxD1dZmWKJBnQRRAvsTA3iWpf2cTg3MoMt8SkIK33GOkzOkCXuiZ6OL7Gm
xE60vdWcZyRTisk/HuPfKSzaf1hu3tLcS/vYbN+F1GfipveTL2g218hRKIVk6RIZQP+eTD9Z/W4F
nPtzOiseIg5TKQfQ3ZCBuV/ELCr6uknv959woCu3RPUL8NNVGAoQClc8/EzK8TrlUWSMunN3aWcE
cLL0w2myhOPSf+AYL9qUF6Rh1Dcp8D5mR2vLujC3B6xIdTGSia+uQBSuXmsm2MbH0fRLveBhkDj2
vxIcFQ3gzYLcmgjDVRm2wet54O3eWKalDEKZi7/5ZZyKNDEymX+OhJuN7Uvly5BbinZBG0SfNqdN
i2BQS2hBL/ltCfy+praWQhfje60J52+ho9c2cGo88DyxPaL52Njz0hMoEZc+/2EilRoNyu81kHgH
f3bvyzRSyqAGAMJ9WaUZYh0cRl6tGZVOtLOLFJ0RT2z6ca5xywTyG5wJsvmovkzyOSD6f4aiSChJ
bJL7ap633lq12CuphEwI/T9tWdqaYR9OKQTGsQSVbOrHGrkyvfeB4nM6Y0Dasi+W+qCwQI8AzvP+
LqCjwU4+BLpbz9w45DrD8RT58nYiaAmgKL0XVVvJ3zj4ov0IKhrqFkXV/BJaLX7NQD4hzRdHqMfU
JFy2benh2RCO2POiYvO1CrkqgGLygpvG1nP3QW9I/23SayN+XPPvWFiG7nUQmGkIv26ZR0lgw6yc
QDH5LjmkwW3El3Eol3qvoKb+49hp5Q/Cbx/yxucEb8LStJ1TRcgqiqVXlBDKqN49WahH6Y/6z19Z
z0cuqkWPt5VAQQPUIZ/2SgZ/6SDnNi9TC0O4r+EzquJ0OzC9Dkbsuw7ZOrx0TeuEputpECi0ca1v
FH1cJfqQrXCxS+3cxne9wG+B95lx7hCvS/jl0F5FqdykRsmkJcV5Nz21T5eMNqcSkWJ7zdoBOAgg
38gOyHnBQny1MBZ1LA2A/f0UvH3m9N+dB7BJ27euM6OqiUSRGFjnWf2UDNhCBZQ4xy03ZQsJa2Ra
5NcxhUWbSgwj43p2hmcvOjJbhU6CTJTAOtsYuNwjdnMQ4ZEUY9lAOki8y7IDV0yAkLLgX5kaQkpj
QNhzVMwNwdyHvW0q2NJm4MxxnB2ErITXNm5lAvo9Ea5QyqpCQdLtt+nu0kZiJlnP543GdXo4xDdE
RCqnhwCoIgCNaRw8yhH+rwy3Y9aiUoNotYg56bDPQehInzKFoJQGMNBDNknNxqFxNPSinwYwvMHJ
BtlYLPpNY8Pc0YbaKEoE+VMsh2UvTC/e5MqC2D2m7SQHVAUpTs/a51WdkgCrM1ukKb81a3nEW41N
pdS/vS5HwPgvYrx7apsVC++XbvrrLG5p4rsMBdC4Uq/tUSvhzx+vaO3mbY0DmNVhxL64z3Z7A227
MjpMKUsRPAhPZPnP2D40gJj6TCQ0+KHhRxwQUe/4j6nsUBwcr3ZbvoIGU2km3NC6H0zhHn5b0ieO
u1jCKU3MGc7F/dRqt2ewtDcyoDOcpLfPi0KZQfaMExmrb5AiaDongTm75eh2vafqr15pJtysMayn
vP4b2s8ADboMKa+PCMnZrzh0FTTRm5h7JnoYhSKavQVWmdhOYMpQolaxFIWcb+fbxdVE528ahUSu
bKmntg6UJ62L99TUTXkQS0nT95uk8Ar73e7NiX2fBp/1zveZ/G6SUFn5UfvXogJxj/dAPUj3aa91
Ufg42IxbYAAmmMpllURbJoUdnveBwKhGp01fYCQdBFUkXyK5hVIOZjpc/W9vWwOwkemQgRfBT3S/
VoB4sZVec3EbqHURWCZ2MMo0jpgBzdODucCB0xqR/ij5yY0T4cN0GRQNLcTn/J7UPFlu0Zjiya7a
hlx8mm+PsIxYM4W3VYSlbRRNFT6/xFhz/FpIxZTceMH1z7eBb7NshLJ7G3vwnySdTtLept3TMTz2
/Cu5CjOx80CfsFJ25A/HtLHdHGZlrcJQfE4rHmeJvOlTRrGC/iwcxbABLwBpKNj9NhOcQb1c2n5p
sqIf22qYis+qHAbMRnXGkS/h/eWGsNDYs7JpF9oHNP0cJa+7+ue5GBZSIx2dstI0eX0RXtga/WxQ
KPWirbdsSNgC3cVY22coBkYv+NBfCwZDcIQnySze+7qw44Nnj//bbfg6cvMTt/go5EGEAjjuINSQ
ygOfukfMXhdEMkXWk6AhtJvoa5svXPw8iRxMMcuCeR6VM9ZNC5/9TEYEaP9FJM8q5xA1e56xRlNc
azeyhu333g9hVCQh9ELiZ3Nhsetv39EDpCqRXjnaMcWgTd62dqbCKXfYVrOqk+/P1bv3wpsKFZOw
Y1CBCF3r9Eu50sf4JuaOJibO4kO+e2y425kpvnMHXcz91g0IqBnG/K4Si8L0zyIZdWr1s/+nh7O2
g1HY0yYJieTmXescdYJXRM42tpXGDHC6fBBE4P6iIgLD+VlbKF7YaPJrgSZbu+djzYy/+Afdo/0f
XYqLTmMJ5oG8KFX7VM+XLslah1I9md+Ka9PPn0ZDBhtFqVRumErgWxIA3P6PTUAGJ/h4xLPGXwc7
mTQMMds8pGMPg7XOrwISM/ftx65FOkUeihCWkdmI3ypR84ANig6MCCWX7HIONowQwmpwzUtdG5zJ
0a7fjAnTSGAjXiR1WkAh9ouBSqwawgOjAIVIQIV4+xl10LKUXro6Acx/ZEIT6AZ+hfBhE/M3SiVV
6ghg5nAphAO0l+NvbkjVuo4/zmGnR4B7NY+MeCJf+xuAOgjDnJA2jjZlyt2430nJcZLSZ6Q7w9LW
gP987GVEZCzSZ5jOFnsBoyL8ugoaGia4ldnJmwnlVIrplv4efv0A6DEai61CREnolNaXoB9eguiD
H5rRC/2/73piWuls81vjhjdQSmdq/7d3A1GZyzq1Zi45iAmzz451VfPDoJyp+ZhiJ6qDF8nbvz8y
g6NmWLPbDehSm3J18WWuMQUfb8V20Rz0q8oV0QtWtptctENY+r0Wkihc2diOwn+fC6p63AqTmhCi
2U5wPRJNVyEvrjFvArKHIZv4B1UUUT54nMO1CEwVwiaVSNWaYFU1ZbdjazMaDzyDod+u+Tqxo8QG
s46qcsLW5Tst9eO8kNvp1HcZgrARq8mFivYK6CaBMERNsBlCIOcoCH63Nc0bhxmVuMO4kgvs0PyD
j+hKTzMQcrQuUnldVXqwdMWV+P3lSKEDOZD8Wartx65szYRoKvKnCF7MgaRRJj23+/s5t2d/sss6
a631uCYnKwscQF0ZTglF4SxOO0lrMeAMww2BY2f9OU0kOLmhuKk5Ij+fw0EMeRr/3aOLh0gintzz
FfmuGIPMpM3hmCsDve6qAuZmhubUXhDq6QApoX/seFs37p1LP2w2VP4rEX0A15O/QzdUeGHhdXH6
WH6i+2DlMurq17Pxx464gHkPxb8HP0F5ILEbm/nqBUvDwPL8DphvxlFIxApX5fT3zygascXpNgUr
QNfPf75xQauPz4ErDDEcCn6aPUy8FGBsJcZNCi6WBckn0DZIKZW95Ql0UO6wBMFAsKY2imYpTy6c
BubskdNy6nDnVUU9mKrjuH9yVQsCgOo3JLYHA+iqhNxEn7BxWTQRHOdXjwZD0yIj2mW56ho58QU1
TTzrKxjWXZPo70MYgSu50bS2cUps4uMM7Bp2SgFQT44eBUCxERFj7aDMQbIyERpdp2Wwq+NwxBti
sGWF0FkGsFLTk/cyglHebFkOBshMvW0cDPxsQyh6CyTpN0vosdI0IKIfjHqFrXCty8b6gDlhqnnk
ZLVAT9owFQtPEBnIZ1fc8iKom7WI/IoxAJNUkfGjo3LG0lhUVSeF4FTyr2rIPbugGj0LoC+b2Fch
Jr7+EWsGdP9PpUcHhT0Z2UqLkVzmqvjrXXobyHm/VC7H4qTfsytAgpRb5LBWtyUqoFRHT5MvaVxQ
d+qSV8oRwZtZ82GQbj9OMb4ewTdxzAS7RN1MNh8liPXg41r8vIKJjqORhZkKeCpPxTRj1hI0wfjL
8/1jcoMNAYZEjdhNXOgCbCUXVwZIzDp0NnyxeswLM9qv/TgVwvHFvhPbYhkwNzv6PLnZkeR1ODDn
QtlCfNfTZSo3rzkfUZ2Pn1ap5UnwJCdzV1LQ1VFDG8YqFfRxYU1S6lo9zvHIpwC2t8irGi4r7JZF
/NS5L+BW7YIEQteZ1ddF7iwaSHyk9CYxNNq7lT7l08yTCXSAfHYUH2TwexwAdPBkrDtzuuVWqGX8
lV4+ggbIIfXOyoC8jiZhHw5TNqEfBHFy2H645apEZre+LZa/AIwV0kk/srBTbSEkRf8gAvq09wf5
qQzK/kt46WI0ZJHc4/F91Jh/rJP1gyC3IgytxVUhlcyS14OIvXBzfxzRnqCuHG1caaJVLUyyhXfH
8W62Fr3ngiwggobb3dIYcbRsMZUm0d9NCQXU0FeaLH8rR9V2Ufn/+BJsn4VkTbZIJjdObCmUekVr
YzWZUummJrMi4W4mXjQad+6Ai7XU+4P4XUGfl5DQkXWCH6RobG6Nw9wJDDdMj/6ZyZJNmSeuPRiU
bZ/QB2E0tzFKMBVqE3AJ+o3FZSvit/HkO7ThvBzgWuG0S9WiNd9N8WlNli9sn0qhK5d/nRklqnia
OO0MrUJUC6Y48w78Y0XG1UjITayONy6iBWbLyy8hsZAjE0CnuOJ3oksCMdO2V1AtHls/1Buuer6e
qPZx43A4EL27RzH6e8mpdBak9gxYxZ6B0ZRGFDxkHssl6CR/LbYPa6Al0Eom4zpWGvF4b1gLF+sn
j8FSwK72fC5BCLSL/v6NUi1wfRbZRun9QavwNa5UFq/k2pofQ+Pg/1WgtSqk11Wgi/r7Kq9texmh
Td0BukZvZR9HD5boauNUWb1tXPaYWZXMmq/r+5hiboth57x8EZlLgfYpGZhL4MmyHVsxj/NwPRab
IIlOPPEDCChbdb2iKqG/LxBpMkNiHDOtMaN2HdCRSI36t560SX1G1cXt63waE8DksHGLzXJNt/0O
EL2Mkd7HDUCXXt4WSjGmkdcXpzgZkaG818kSrCk1C8YWeDZqNCQ9hn/tHXaJQOokl1ffWM2JzVM9
mXDHH4Bm61bWtvDcTNaznSUXpRbU/vXioHrl+Y4k4uZzb1XK8qK6XGo/Mf31G9UaNe4QGIziCJZ4
0SzCMdMp9wAlFSpMzZyx/xWBHZggje/Cwea+xGBFQmPwEm4ayRyO7wIQ6cEhXDsPhsDJmlUWYWZB
d0gSZt1WKqWDdwwc1R9yL30Y2qmUx4M9mbCezrPVDloEXknB+JOQAb5TivM09jXhZdXBUIk0YCbK
y8ivwRTv3nPAwxavfaIr+ewMOkhRxnAXFARLsyErMtHaO7689FMy8L+NPUOfPpdCHRgCdhE9th38
V1xopuN4JcpJTGdvxYpmOlM4Rfg88W9kkP54K755iJNjdO5aJkiOz5zwYh1YjLeb95/hVAG/5X7r
p5vBIoYqDQ7a69sRdvdq80SP5KAEXHV1AY+ZY7npe2huCGWdPu8/nYABNDaeE3itNAhAHfcJQUA6
+69YUzV1MWaVaTx6ypUHkc+fQAR3xGF0Z99rtvcEdELuYHYiaJt0drRwGXMneDLFoXxVjKKesEGx
PVldiydSAxrS9osVbWh1aHucJXGUOGd3ExEIX8AajJGtCWQSIeDN59FkJNS9Sny/eaDVKdwj1nVT
p51p3Iz4a5z+kTrSiahkTDONbGDJLQub8xIdgM+zFW1fpBPUkUg/61zjiNvKlq2jHSSgOOkqlD+s
blLbX1Ba4aqDReYHHEXSV6c10fOC4KvvINOn3inOZXOPIy7ec53EkPcYQAXsjuJ4phabYgeRyyZ0
U0JW2WJc22+JYPUCAuRcY7G3eqP2Xxxn8ei81GqYC1CtkwwbeYwPBzR5+z19t33NERWVDWM0BNkh
E7IEpBjVurxkrnAcRABe8TQIasPUW6v7FNpal00Q9r0SXbRXl9ZQNa/Vvr4b9MRaIr15btvIrey3
rUR9t/+LttMdOuT36zxqca+1krR7wFxWO66U6ODQzNHNSQySTqiv6XtzRC1uvKcOeg/NLRF1E5KB
71fDXOIW1/FJyrMcTb8lqXUU3IEwMpXJTJuMl/hubA8hKcQHbfq2Z017befS7ZqjYNBS5QnuYMkH
PAiG3k8GMEavPeov2gdWEr3eSUs/fWaSYEMuicpJtuQsIr5y11+IdVgxFvrID2BMNxNqlKz1Nrca
fpklPeimPInTvhBwTGopIsNUFyZuQ2OVViaWVZSWOVsg5+vgrdtms/Tt2gVrH8/j/A8YOF5xSC5W
FuAAmyd67qJWyN8KUFzJjIHBQLP0kbenHmc11zYyEPGHw1nkab/ijXbSyh34DSd8mOfqbQUYPlC3
2MlZyRntXWOjl3rR8RLLzfIkRF0JJIzSccaY9TavBef28iErgDc9PxQJUBgIHZbBzgzq5bqVrhXZ
tidGrw4iPGrfMBA572EuRSeIv6CTkwAQWpwmFu/xoNUalrYmb5TQNpPdOQ8RUZZpRkMOqUY4QGDM
uvDxtcHONzppM3jxXPh+7UNS9fgo0pS77bmDKZzrBEt7nNtMoQgx/hQKoAbdutDwHGl/tTL+Y+Nq
PtZVU17vr7lalhm7RVRbe61u7HEUMfDHM/xkaQENYyqaYBYZWF8fdsHM+3haBAGWFlvJk5SVmEib
otjmdwXSLd1r2TChkMeIv7FXTggO9yP+eM5eijW0Z/kCC6SOXG2zvwuhz4/KUhLv5KIiuwJY6xrz
NkEcrDwIVC9niBk5wNAYpo2WBQQQK3o8WTvUXftGXshaSPoz/zEBOZb3g2TNx0Dm0baJN6C1rtSz
zgWWmrDg58YnEYV/AwuWtNGEKGAVvY9acqM2xWp1IxLOiDJagnB7VdfXWXdF5NgTFDObfnPfBsvF
thcH5Pge1CDNMXlP9uWUvWlNnh7u8S+Iby7KoWaeTgs51B44FkVKJJfFajmlIj+IVPPSqEdDEgNP
ToqIxHWTAyfbje8BFFcJNXZ8WvdDXSwROYcSG4yHhsQGuN1Ar99KPv0JU2iTm+95Fod/HnoEDgOf
gKPPu13eeaRw10nzrNkzmF7EvnqgtbRqhx1WHDRyGkFii9rH6M2RDu8jYvpb0dh7p5sI2IC2a5TA
NWkhSMcZjKpEsZo5VNL5GPwPBZIvPVCVzseAY3/7tDIqUrkavRKS26djtL8MzuMbHbtOYplOiIlJ
lub+LyJSzjA/x0MS4gdiGPhtQwNUr6SOYTDvwyYt8E4vmlOnGjKc7ZvR0XwKBHuCzzic8U/DmqFE
I4jGWZqefpK3OKj3iXbtmpVTBbBpDjujo1MJytWNsBNvTYBnhIPk4QU4Bp0eHzmdoo0Vvca6wEFv
HJt4X2gLthTNsyYKTAtYDEWTFVu76A6vL23jDiMFlr1uk0ozKb/82WeU1tug+67PEOGIJS+dbx3M
Rhhnwv8f1RCa9mBi6cUNivE8YS6v+XhCS5tirv6nLzkRyyLS9AODhZGhhk0Uc8+xk58/sB91OEJz
nPfldyw1d+EqWLewGHG9yF9oGyxNO0ARIV2AvUwewtAuhS366Db/w7mZe+3ok6VuNDsr6CpP1fK5
zXNoOZ2OtnkZt8/Md3wPeVzwmzKQQcFeTRsErFI/XW7nGGhBgljpvICoKOKNDGjzevB/HVkZDKqu
rBsnyV1AJVSiiRuXgB41JZdDgdorZBAMbQTiNonGf/UsZ7ZegjoZ+alAeAIxx3By95TOaYK0kFnA
Glel5dNjamcINlxnlNodS0GyfacKf1jy0PbmiRhGiPjRyEJHhVUEe+z/P6KOIHR//Hua5d2xn5Hg
ivAbd9pVNjU2aX5nAyBSXr/YFp2kwaRXke2jaWSHkl6kA5cnsvxtxv+AuzaCQr8Wa4f3SBfReA5t
flfK7jS9AiW56bEtfMfF36N7Jw4+Jf/LZo6Bqa2E4ccY65EDBOYiZwI97Fq1QLN7BEsxrz7oNOC8
ienSCCc0AwqiScLCO9mFh2LMX5f+mnTqiFNoW3YY3RuF43ANKm43v+jQsDKdx5iPUrFt3dNFEnis
8TWQvpK1nMJeiGv/lu0mOpibgBcdOoj4j1Y/aPfAG9ephckXuJDUTEpDkpq/6m9uG09xHnZyaWlH
W6Pji9cSfBa8Da2IbU23JuRuzo73yxMn77h4m09NkO8R68M1OEJ7SqJ2ou7n3djeS95sRgDDg4PB
md87euTfW9OA/XHm/PRCJCU4T4no2HJAFeSz/mnkic6OXV5JJUKLXdGL7fhzZEHd7asZ2+d4CF8n
q4Sxuu0PhwS7xLX1qgeU5IF1TK12xAqxKNAsfqo60GzglnYSuQGeA6tQFlsl+VZfbOiKl4OX8Q84
ITamva9Lw07FkAknPUTpGzGXzdRMvEQFWoj1liqOKMFhNuL7mZAJEYlJDa70Lpk0OX62wZ4PFNUz
X+BKFCTl3lqT4FqajsmZc07/N+QKLCVCjU601LCqMYEqHpQSt5Tw3SJQ9uNloTeJCosqsCyOTvEA
l+KfhMNZEsY5iP+YLOMsM17/D2lkXymd3UDGLZSe2Fw0iySscirPkzxrbsC/7Lq+y0F4sPQu74uA
m1WLzL/V7dyl3+7VQbQk07T/BxlLhJnmgeZGbxu/xXzOy5FKitm8mENGWg2wkzYe+rxgMuoNNQD3
9jrQmupLLS6TWsEApRSaOZIrGVwqfxK2tArdHXSy4Ox9Fj99gcjXnP98H9hX87xQMKMGvDhKYPKD
S0wlSCBVTnFalbGocft4D0qQlAQO48+Zx1BW3cCmbQ80atUQX4QiDo+lHKY6SGiXfRVy2B+VlruM
59ehxW/jLnAQTIQgzDKVSeGb3dGIeuH7xht8BHuKwUq6V0QVA4DPwuMl6/UNGX7CcT+v+QwOqV1y
j9bsiFEsxABx8LJ1Vgerl5SuvQJhjYlJIR2boOyhsjXWMUAbpzfv7i4UDYBP6EE9NX22nc8CJyO2
SrAUE6W1+eHKpcug0s7PUksvUONU+K7GmcR+0z3jVHAb7JY877WFPbGBSotpP8TA6E4EhjH0aTkS
5isRW7FvTYOvToHX8pQRbqSYLEEdbrlP8l6Kn3wlxsz6RPYSyqca5xKrx6HCujPFKI/HjL+V79vT
mXT96K9NZJ34vnX8nSwlmlyosCA4/xxA9/UVeXRjsL+bN4zvfASU040+XBJyDaQMzt9prndFFUWK
m79ir4sfK0pbJpeG68CKq9/aBT/9xJifGW3l+JzZQ03RubBGuHJM/US6NI6YbmQy9lH09Ku6NXo+
FWoDJoaKHH21ggw1l3dOrUMDYCXR1Eqwdu6vfAw1roZrylD4os/bAtZ831a4y8PVduFu1Ux52UwU
YWUHEYhqltbG99WzEhXHn8L65nGP48NM6zWVsK8V4SNcXxW426kDD/oRtkdSik7spTIGuH2ZdiRM
sog5s/PbdCU6IRCPBdKRhhmOP2Irn6AT4PNvRTwyQCmXEhfqcbitOT61ORAwq57Npdhk6G0i4+Jz
E3k1VAVxgNC6T3KAkJSsmdoJar2kEP0vHciX3UzxAkC6pTWj59L2H+9PCWN4aefu/1sS8ZqOJfzU
CM/wZmHP67/rRxlHuq8XSZXmFEgSk+21yBdf6/aSrlwpQajMYKa/qFSaZYqxXGJaxOcYqwEXI87Y
9CC9VybKzP2KObGxeQKYXT7woiT2MvnU8ynJAE9Ci6YAo8Hg21ZX/wvM+hV2KDEWDAoTknLfcHaY
v2N1hCG+mxzh4uDSeTbmsDBFoGqclqpkPxppcrdoEtC4xt7P4apgHab27P7SpYu22wMowOqx+WWO
qu2MYqZkZtyKu4OeOVDpwLVmusihJG06Kc53KjUpv1cXBqOmpIvg19pjwjEz2A2becmvIDo7pv91
FSCKPkuIDKLR07yDz1xV67Rdw1hfqd2qanz/7jmQmHm4/MkR20Wzon1juqv1XRqe+UMFVJNOkdj2
UVQlxzzPVWqmscN1mi5qe88L1waAb980ak3bQFmghmcmgmH9PoKQGEm5Ec2o+hgqK1AjMLslgx9O
KU4iM56I/CowtW8doUtH2bHZTYGB+LYLNmvdhW8xa7OFdxtJOUbe5WPeClRl6Da7vkLqj7mlaHcu
5F321kcnt3TLfjQD5zZf17SxZgo6oRYd+/k5o+/bI1WjN1QOBDP1QL9luYUeduaVwlTrR7LTui0G
9wNraRn1im3xb7lBpOuK/DHpgn93BEBsF3ximwrt6+MGK1C4Mg+bGBYq9bNegbG0GW+x8682UVQf
y4CX/FfecktR7L1rVora2nvjHJ2E9a708NA8aFDUiK4h4xV4/oGfvbCtOA1vAuBrOwcdGkbkmK4W
nDIiMEzjsF/8TI140ZaiaWe/HDusT18MrEUYYQRfHmuOxjM7CY5V7c58AhMoGbQ+nrMNeAxJ5C29
843k00Qw8VjzovmnNh93S9EoOCq6mF08XSA3yF02RWvDetGf8v48li5OUeLfeFi8QqxrHHF6kOhm
/k8HmFiVqQymGRhTgTIEUAeCjARQCMfOwFvwyPs3LgGwa9tgWuOWY8KNHlgmR8p6JnyfTwdTnbcl
+d/de9gnxBVgoUuB4rhqxvOsomUlRE5R3oVLFVIGDu8pSI+v5eQq5HQ62bBuUl6CH1J5HuZPsZ1Q
bHUNA0KIJs/weiA08gScmVh5uH/EalNxWiGgUQ5zUQ3whOBNBE1/EJh04wihRu/xVNIU2Yli107F
SqPPxPrIRiTeaNbIVrYLiNZAoVkcMpxv4nOEK3S0SN01seojxdKA6PS+DVlyqjPJXZ2j0dqVKKYX
bIqzUhOrfQ25cU8H27L8KmP3U6EjB1TCTFie0jfOKg26C/lG3cGSRy3PW9S34RMob0mH6YpBWQCE
4blWnCdI4uZ/hej4kRwU1DowZkRnYpbCcsIM721Z5sZjCLB5j0gRZIZ+jzhT523Rt/2NyTsGNZtY
SZC+rdvuP6ACIdn6BghzIT4zcFWbuWc7VfAPEAcLtxIxQSwI9ab26oQOPQHFbW6XfsCOgA/3/aWi
zKC0mP5Ot64b0VqdwQynexK3X7zvl1oe/sKSGnQYTmvT7OYcPGgqi93sd99uVGUZtc+VA3fAONaU
1o6HtQHj05uNix8ZuAdQZjgrWxICHKa5czPlVuv3LNwa92Oexc/csStbvoA22ZGR0Q74DesiHfky
RuvABl8a85mI85uu0gl0c3VA6SLmmmt+l4oAY5TuFPD3j9KQBFETy/u/cX+puwhb6Gx7tRWg9jpI
ndTepYhWEn36wp5dBIb7Mp1N7gDM0dXhszEfyWkbCDDmpNZbsfKydwNc+ZPnJKV0N3H8Z+OPYg2V
JENLUbDOFscHi8/eQFM/DFgowgfBg3pV/Hr0wbwv7aY+XdLj/Vx6ROL6c1wJou8cqpQDaLS9nD9d
jW7s9fraLZnZ8YLQfl0w4nbjTdy28ZZ7ZvXxP02NmWH4VnrWajJyKxybumaewva4Pq5pgOPdVByS
yskDkXNcPL9okCaOd0NrO6oXLpcTXqtEZUl/zVeShuEpOsBMtbMAjtpn592e4FtiB1BmpYs/lN4O
7AGgvhE+VACQOFiP+dzt8GgDxOCy6tCs4SHYe8MCMuv9OT1znUgP2fCbqrey4+d30hcjJoSaruXR
W537I1XR48YJhK1cy9MpqqATTMM0u62SBYZGiWW5oYyBW9HUvx9yzMFIjFLFDAJ1Qd7nt9hfDU2T
ubN6rwhwWdv50sE8CRAcoRsZ6fv7S5/ByAJ+eA+F9PI7xivymk5IH0pWZK7rW+Tnu5+Kk5SPph5s
hvRy0Pf2sMv7x5KwzuapwMMotkLfghW1WoE8WjLOdBTIuFWy86tulFu3Q9mY4PswMiZOVvQdGLFQ
e2iwMVagUVvRxX9xjHkivY8lWYbkW87HA4BV9veWcWJ8QCFBC+q+vm1JcYQP0hp8+ZpGyp71o1Di
vUerU3Mkg4AlzFEPsnyof/xLwJNgpRcz6/qgHZm3Zqvt6c1fvGljllbnCWlf/yPyCGHTIOMwOgQp
eT00J1Davj3RIqASWyXgmBbqmnBmd0MAEOMW3iCogtytAx4jx6vc32eQcfeTKF0NXW9cH9rnX/qo
5OCnYqIaCFtT85Gs6JMxVxc8ddtjUd5lpqpgjUZ2P2xNKMrU2+mxJ6VaJF6EKUdhu0LcWdv2L7sM
xozVAoZw9oT8pdW97f/XEMgv+o87npod9jWL8fcU7F525MKbYgVYRR5vu8pumGhDyCMxdxIehv1j
7RzaeJi9dj1mwuZ8ga6z9qvDxclrkNcl7Px2tHAO+OkmbahNo4A0ubkAI3FrxH/A6uSMXTJUA6kz
B5D7BEstfdo4xRCy+XOh8dO8YN6Sv5CQiD8YokrGH/rr4kbsTbwrKSNVNojR725uqY5KiLewerrs
MJjOnEV9VkJR+G6NT8WPJ4WjeFcUs3Ly9IjXIdxMnOWgODXCVhfcnXrDURavVgsewb3WfUdlMTWg
MUrVS8kPakB/LUFVGPjFgayITF01z3NXtTjqvded5bRm3K/CVm1iM3Xlgt2m8aL70F/EdKu/GxnB
Uw8U/WTuI8cmAeLGgK/Ze0Y9L5x9OqBu7FNaRX/VzBsKL5BSTeCTAaQANH3DSWrt0CnbrPw9N2Ir
bgpeczvw2cKH4pCSwVphqi+kehgAchhZZUttwwROwJsIyef1wonQy5iYXFEGZ29QY3ZyotA8ybvW
szG+ejR0ueLMVXS3YI2dYebV3Jp73A66JcEiO1ip0QfkNGtieQLazykkjg4ZdVNr/4GJwnx4LimJ
yLcr+6V4xaeMwqPL/OSDPWhP+ls7rL8Dp1cLVMFrCE89QQ3Q816/kUvxaTTndDsN5x7ALQkFfKVo
QJPH8iohaHS9rsuOhviIPWAGIkc0gNPZPmwtpmHf9aG9haUKf4k4jeP8uocfk2IrHVs1a+yhUkQH
Q1dUZnbwseY7cx3dBoJzCCHWU5mCbph61wh2GqVi8L0XFyu0Rd9kyHZTeq41PchNOfTeCy5Fy+Y0
GfRNy5gvwaDTTolqp8+pdjcIxTVJMkO87vwr2bzzxddmYd4tVwTCvtLkf8iwIZnQuBFZev+k8QY+
I2eXjV+mZw+hEJnOBzlhBEExo4vf3uB07jTs2/rAdEj7JQB6Bin/SR6W/zb26Kb/Br+xEBCIwjNI
CZcGTzrkUO1N7c8XWoM5BAt9QwU3H22GUMrnturknRZ46TpRXi+aJ9D7q9GRlVV7HMU7CNC/7oF8
ExDo0JudVjR966wSIC1JP+jxNPeS15oPK+pJsgqWVuZjn8YJm3QKDMN1GqwmMwshbMl1nzoZi7pH
BnYzgTVDRFZ3KpmHlZBix1Lczwu0vTusuO2GHskEbKY30Y/Uf/bgQExYa3ea0YPkXjMOuz9x2xTd
CK+lAFeZbP3ypnSzYPTrMx6Qic1tZJ8OMHuYi5bor8Kv/HmwT/IlqgZax8+vWvgb7/YCGvrGS2J5
xIZWBxUd3hwQON6jjPhKYvUoTj0kArT0TFX4FZmnHQMUwcVUxjTkimq3s0SotabuR/SfXfnBPkql
1KsdWMguWmiA2WRaFw7eeI2Jj6bVRmqgVzvIpRuTnx6RjhUyRhQt4A/g7mIUneAWx/OA4QAvlZK8
RojXn2KvhciNZp+UxWG2FllIc13lgDnSpyA8yiUjgnXDDS62ofysJqoKeH05OIn/Wid0SzwodWkV
6A+VVZJ60hDzXmGi09zDiBMbOW/yBo0GC+TMOnLO/SRiaADSf9rBIAUlVtfpcpMh1IQ3gXFR5Cob
Ex3/Mk7SVsRlBqeWzg1FcmRtlsu3OA0PvzGAI6kg7MV3slYJchHe2De8R15LD7BXYArzZCXgc8ua
5ZO5pgQ/a0FR/f0YAYVpDSIDg+qrjaP+a+IPZW0BuURGcE4G2IhKUKofw/gh98d+HHGUjRBG6t4U
0L4RIzgSzPkbzhfpUo6ysS3acpYJVath9FL9ygXBpk8jwDsmeI36vYSe/JP5G5pyC/jFbE26s/Cu
ZhkUspusfnI1qANUQeNZNPO1+tfTEWchegveipONQrfCj/mkxFMkyBidk3qp4jmC7gs4JMBrMShG
6iP/zsZNn2kvSyFoZSpl59ui2udOjk7ETRqUr9lE11uBiL8jTmGnlIdHBoTV+5DgKDhAIHrZkJdQ
lNvLPU/HwWdB+9MvDzSYeX8eBSl74fkUMr5rPcF6UNd6h6vh1s1ixBT5OC9fKu+c0dZOtrVypiSl
KjxSzIF0b6SlK2h70UG62J2Nkejof7MZcrFU51D/BoFGB1S7awfaohvbYSzF8rdujRD3hhM0aXYe
I83uJEsBjGsZvRSKS7OkBOlRJq+r8Hzw4LRy/5Xnp5fTH9ChB/V0R3cTm6OasTSQxDaR0n0F1c91
7lO3sgGrcsfAOFxHRvUXJlves3oq1INxh/Uh7b7fSZ6e+c9oMj1P+ixfQtBc1tvr/pSp3VKqXluj
mI+9yuuvEHJ5+TtI83LR8WW7ih1PCioQSk/DFy1YWt+PzUvCZ2xZG49dFJPWVMVxAxgpkXusYGPA
yUaxv2CNLaLhldewKbmc3/54gcQQdjFxD9CNiaxSONt9j9o3WEp/w7FD6CrA+u7NUkYT761zEGbA
vUJsgVij57B0ZyoOm5+zrHE0a2DVPP4LecSlltDbXpYLpPrEcNJEeSrYlB1VpBaIcOQSCF3XlreY
/wLyXOVGJpRPytBkcGReyEQniv+iR7RWJpp0s9QR331XOXAVZDUNild1e/uO4gouRKluA7FF05mY
dGjVg5/6dDG+xzNQcSyvvk0MxJHR/8DH08iloFsaXLeawhI4QbbKKPCWs4VsV17kPqHXkrg1ozfv
COuMZwDShEtwaG/J0JUSPofnVHzPK4Z5kQaVx2psXkz5+1dD2HcFs8CfzTnYgw9z/QHsk+T50N6C
0vWLUh1BjyRBWB6QQHuqSt5H8wPpBhWdNpLTqH8s/3lJ2m7AVJ1V7GvjI6ouYKTjV3VO8Q8Bk7XB
LoJe9Q2LCeiM4saL6kb34EG70gg8G39i9609uNeH7P0Bzc+bDetGEjKmgyva3X+XtGSPxLNSB2bD
BwOgDGIYPx4BH25AQifZOheSy+D1BgdZNZhXE4ws+4gNxRSa/LL2eCcPHRj+TEwUvb8SRkG03Lnw
JX9sIta2cFGWTayc4Vmr53fZiIo5oGdobkGko/hh8MYZtwXMfCrTv1ol7uhH42G4lBSPLR87COiK
w6nBPS2stJxHHOtQ1BKL+5d9ydIFf2Pgq6dOxhkTxPnBvVh7J8lukmfCdv5MrPNsCFq8nXMecPKL
8g572fcwTCOxaibtLFYJRaMMzFyhQ3CuMjYIk1OOt8oSqUMb8yVcOMpxYHRaUAZcvxT85COIu/z2
DcLB83i+alwgk7ECYEOxSM1CtF60mPuwY7psD+Wh9IQbWCabPS8fZzRC2jNOPELhrhYd017iLvfE
46GOgpFCbYdveAtFBd/j1hS2dA89F6cAVcNn8lQIYrmVDv0cBPfee9YGD+Teel+GPGFrtU63NDBS
XVJejGFq00qLrULXZHLv1F+LbV5RJAWiAAWpLX+OVeFZoZUxWxyugWBkTH9lvSGKGrcOWNrlBA1y
OYHpKf2V11fvIC5aA0ASYz9EbABB2VJbw9V+AS9cGw/DTE3ASHKW9z0mo6Snvl9zaWZV6jfjA+Yv
gpPWG8KfZ5wZPYzGKfCmokBiPgoaT+A0dWz+f1ykyZ6xdiditkPGD7tY3mKS8H8WaT4VInRxOcRI
GBYHeWO3j4fD5ABw8+/1uESyMJL47D4Vq7YRZ9JiEADuq1sYYZgjDOvDJULSFX0uRZ5Ta0veOfuZ
4PfRmCs+nmbdjhsoYmZ7cIs+QlC8ijljcM3b0H63s/N2FwD1lHFWweISEsoX61R4AtKiTRYwZEJq
lfQAnJisAlQxQHRWIRVFFe8dTQ9c9K3FeF35x/B3UDj8HWCA/FQrYfBu1NrEPhWKo3miVsApoZii
kuDg04BSWfldidt1+DuOcrr7FxlR12jOVUydbjsnWeMb+uaNd1kzSJZPZxGv8npiy4PtlNslO0pg
j+ceGYLjinQgT/+dE90aGeqWpHpMkFD4OisMyZpV3f4yPGEsL9BTpQ0UMisqUXKxLwwtTV23c9mq
+JR+Yhf2v3A1NU/Il+bdlTpoNHr43Xtp13YzahaFf75yiR8X+NVW8jkavAAbVUWyUpYlG7VDttA0
3rMk3yz7RoBzY/WvkNtD9DXqucAm//hpiFpX3LXvuTemO/0ta7ijAa2PiLkn5Mf9LxJPzvgtlz89
aOdCqVrKe1Pnprt+1FxdjwfRKuA4coJcZVRH3GAulfWOKCgisRitIjbFtkreV/56BhXaae19xK6x
DLV5Bz4A9pZHuAYhkNw/S+Kp/U2o8wmgA98jdscXtqqvL35XVSaqZbIt8VrXdHhvkrES34WvosNX
gouJ46enhN8xCMtIP7RIvgX6mRvFvNo+vmInpXcV3tKkcK/25AOcDAOgld5M+lijXN3ES1CzwD0w
++smga9wWU4M/p/NG8UAX9mwo4oCmbMfjAQqqBjO2x9msbcaHjYJbu/iHJIVe3E9nEu7hTBvgTpN
KJzi8x0HlX8o/1UwzgvRFDixxrlgRbD3qnapu568QFlV/cR8YHUwRvkgznFyV7zunflxKKW3P6PY
Zp8pvYVLlEsn+pG35BBSkhWbzTw3eHlAFu2gZB7cSNb22/nWCG9ETLs9HE1oD2D6FKOTq+1D9AqR
WXon4BC7C7OECH6llW8Rby77IBgIpqHbC4I7CPKLjRUsKM4/YS9g2lA+jObfUszHh0xuz/6Grx6e
FJMQtqU12n+fiyMW0UTXDcRdfqj/T6mkh8Fvq9WgtJJ2j89eOT2RoHkQZF6P8/uNWW2mls4OO07q
PKNK7Kv/e6E4FX1Z8Q2/1snjnDauuogrpRel0ofW821xGl6lab3jFoYXGDO3El/cQejyfZawgida
i+yWTaBCO9WhNF4ZxO0QXud07QPU+x5OrfunYwhnS7dK/cYDqsW3UPHz8JILTanjRhi7fKJ3UBWk
mIMreEp3l932C/xL6qLvuOdGNGMPLMLaUtvpwzuSBQVXyf0TG/8Ls2IpXHO2mUpq9RJ5iwWEu/5Q
NDwJmMPx+bAyRZXASZaxfSv0l/EyBOBGbkFa2NToY4VX2PKqBTR8QagCv+VMLacpg8JN0aUQS8AP
L8FNVTy32WHjsnilJkkDs+cnR+vlx0I/8GhDlVQ34A4bBcskBCFuYOY30iykT6xjWIGJXGTpyXOQ
PYmIM9pLCBd2OkgzhcQdx8+66ZGi2bVxVh0GgwQG1QKqJrml1XFi+3pblztmSS6kThiYjfsOMi0z
N1xwkBkU7ibe8n9lX97EyFHaVux98vE10rKyZrQzwiuhWC9j1OJ8qxxYE0n4oIWQmFhjqVwMw1BJ
VAYlbxmlwbq1Nj4dN6E32eXMFA2WfarnBaFoe3p2ReOKl0es9aVOPWz79uZYf1j+NG/hVAd39VLT
8y6i12HB60aGNc0nnkg3/JmTp0r/mn7Yd/guVF1rwS4mEfq8U+72HvtNL3oYF7jCwGF1KZ5LBKoj
4fR/PwFiicOfpiOWDivhMNaflSnhg6MQfuRHQt+RoeKnCINebO7mnJwi3UKLJDZnHFCUANb/UJFx
CdG/qKht+SEJ4VyLUjZ8nroN527q6ktwazOiF3o6l72mOgwChyk2M7mjOHPVrDTVcj1bCinNxEMU
Y1v6awD+IGv8xovEkthtcX+Kr7NJAHt3kLvdIp04VTZEBm84noJ8X0/jARlelkieJ1lQgLZpk7tf
VQ7z3JrPCHPVC7PRFO12jWdQ1ueYZeZvSky9yChLbeJO4W7g6XrMf+XukX8K5tRAUS/c8/rmFO7p
Lx9pEiRI6J8zli7a0VkkqrUBebdRhCGbApb/OBAgEEQ0hfjx6lrjEq3BTTdkefR5ygtcKHPnmR5s
Hsxi9MYmX+Jnf0OMfqWTcIVDpubQl1MReg9Au7gtpAdfPCoHZfFVXEVVgHAf7GMXd7VBKypkbNfn
krB8Afsfkuw6Fj/HkzHhQL8Y1YGn9RShLK0gdwvALJYtLD8HGkIAEtXV0mJAzTBYFK5Lkh7egLD7
3F4xvdFa4w/YaZ26TcJ+N3jqU41noaeJ0Yu9KpNLL3sYNEnqDOv7ippw/enoc7tHDxFP2vUG/vwM
ZmhLRwPFWvOG3fLfcbwaoOlEwPTh7rdYHvmBYOLsEEZgqeheqkbOb1BlDOsOqfYFVjWpIvI4Uq4g
7yaoM7v25kmIOOuzkLFxyR6KHguCvenzlcCst5STmJMmpmG8QDH4PFa8ZfNMIwWtmvJWQpXZitqA
nL13bFtLJDq8U6akpZfsvKpAdoBF+sm4cKAXwqNxI+Q7QqwHcmdR2oaXDaZgORsulaFJQzzNV4Ak
VI/jFXcEBYqrNUO4Xnyffm+4c6v7BYgFEmgtEwErhBgsyeQ+jR+bIGpXPyxO9eerVglrB9gfx27F
NANxAlcm3oPw5iWLupwPqQOopiAyzhXg3Af47K+hwtAOkquQuQjTNuEW7+DgH/fADjfi11xQJqc4
e/ym9mueBZ3R/hpsUINqso/Tsw/kz21GukZyNgovRKy+jWDjmd0CoO9C/xgS2xqqEAxGs1zLiAfp
5HFs6SL3RlICXQkVHJqSSmhdnDp/QBNM8qBm0nLe7HMUZCesSZfyb9NbF0Wkcq3jdSzVRwETG5B3
LOFK7NuLqpIBNCdGqhWKX1lA50MHs4k44zvWCkUgrhXkIQWNy/wYk3L8T1LhObgiitbOlMEKmnyk
8FKRhgeEgSCKDmKc8MlOYwB4h+nfSSTGGeXJOSzWTcRlpa1Yvzdbvoh8bp4U1BRVcoEN+nckx8P/
5F37UWeVbgtw8bG/RT+40YTWdyuZ9KwR6zjpfeeC/CUIJKB1g7IP6VzLqcVGwFdZo/dPcXTmo8JO
6JRQEPG+Yr3lZqX/9CZpYw+rklfgtV9fULpBRcs8AQJyqSJku1HYhdN5/0QtbKWTXtN6r0NyfZbq
xr1swICz9Tqvi4rBRo72PJrMP6HOJ1F579x/vSjIchzHH5N7/ML+GtBLHNgD+Z+owI5h6ZRpCABe
WHHUulcyjfIOSAWPAjl1vHT+97su0ZZU3cf9B/LniWVKdsak6UPATdJ+sycR5qVm2AHYwIjSuqd9
yJjSHj3q8mCJOzSWCnIgzGw+aGrhaPrOk4/b6SNEfFXT4O9nFmssRSyPaMZRohizH7Ic8CKtYj6N
MTwoxefQEVTG974dmzv4AtCRJrCPA1P3nq27F/QeNiFOonhLvhzM3LXQRzJIruouoZ3urWK81hms
GAYwj6kC8lKQf7D+KX+lURqms2x0Aa4noyE5F59f3XKL+RJgoHKa52xWFbCmmC6gvp16BkZXAjgZ
jM0LglaZRvkN4SyZ/SWpq32hfJYVbWMaO3O3cUZwDkvaoRk1T2fOxDO4WjGd+jq79wY38K8Fs0D7
mWHT+ICWpb8PzrBdON+f15dp5ytcqzRhVO7Obt3WVGnpJXN8StldG5t7Zr6z6adHzwSYm8zYcCDF
iUwBeTr1wyjfV4gUQb4utuC3ELtMDSDeXbzkiV6V2/YVimUcyTVfB8BcWOM7O1e2z/T3q9WCgf6+
uj9KfjRbWO8urHUcNj6c/bjIr07OeOzumpSKqBp4IuUzAR/OhCBZd5KiRfodNmu4aaL2uv0uASJJ
e36jXrq68RLj6XZWLoNZJWWmF0fYmJ0mFsA1PDuQ4QIPREfIEwqTZzENZB9/M4JtYWRdK8gStNGu
VYB6tI/SddmY9IZHMr7Hr7+lBSqyWLcf3K8KXDa+doW7HEHIILXAFGNMBRP9UOCPUKlRhpm8drKY
hp5pibdfpjQabTkrqewXFfUwUhOGqzT6jW2s+5BAingaN3p8v7sGq2VSat9g0l76nOdFRajbXawk
tBYEHpSDP4e1gLGp41GmxBh6gzHLkdeUQuZAg+1V+2naUV+RfZTrlWrjhS3oyXjMp1DLGXA0egIA
3Swbs6g6cFmJqNi0Bg/tmXwHodAFvPxhZ1Vm9Gm75A3X4gd9TRKqS352yfnRVSIBCIL98zCM9Ov+
m06mRQ7aw+FhwxNDDNJjAy5mNYBU7Quk3VpOnTe9kyJuzR7+Db9o8n1oQ2FjuZcxaed9uihXt8c6
sBLtBrU2fytAmvWqfeUh0+tg4ioUmc5GtCIZjlm4vkDml8+ug3qfSW3JPwR3w3hPTYdiuqg8GeXj
Tz9w0h3yQAJ5x4uhbJAMxRpPSlmHxKF1NCukEhdxN7EpoQIoMresTPFXCtLqVVXhJYOkNXrCE1k/
QjL+rEbhWweXxyyEHWT28zE3ypbkGsHpmlLkcUbjR6pioLBfclMJ3druYVFWx85HkMF7OqOBH8bB
FgUKPqJ6EFy2bao0jzN5L+G/PJHr72z82QzO4d/NQpDri22MfG13Wf13CZ7QPI8LsoYUcIZEtX8O
JgHOkKo3azBMN28ESTuj3T76pGgmB3baMy4+ord4zVGjI7puHKzMBnyEszHSsaMCvFXzQid0KjpU
ckCzL4PRJuY0nT3LDtRQHAs6yN9hyVqDlMhjsTGceHAk1jxdGi14lAlofdBXeGLuXuEMAW3WYcom
p1sipq779i/wYtIvKEo+MYN0pCoyL2oMROQEb72sHU1d33eU/BvHc8KnzvSxS4+ctG9JG1bHqCrh
oRY87ewHgAD54knjyAnO/pmlhUuF0EuqxUU9hRKCMsRKZyLWA35BBF6bqFffS2NedroaBm6OiRc6
9soQSlyH21+QJk0S8kGM8hRyUyMnpaTpYZKe8S/w8qBFqirztKd2nn6Svwn8H7/VNFZkB9QsCX5Q
Znm+ebhT7rTYNUSt7Kx9dqR7oLqtGoWZ2jWo/xlO9qqHtkuplDFPoU3G3S3o+dv/p6BZ1xgd+uvu
rerXHzPDkVj1kh9SajyrZeXtRTCWdUpvcr9BuqifvW6vVKooYAnilD0036dsKTvz57lC+d5EP58H
YEd14rbjXRtL1xB1WiNWiG+9l+3Xz+udCwsXTSywPA10ZWxl3qGBwdyl5g46sbaFTw1j6E/4jDqv
x1P3Wuckhcz1kga2oJO3md/G36JtE5Lz/uMHIhjigTRRUtJcK+iWU01UvdrFUpiC85a/fHWfz7aD
ErQ0GNXxucT/YyQORTMFHRhBACxbbDCutE1LxFaWfBysGTK9d304TSLE7S17glSB64HYyNV2TLpn
q8IetWU1mqnPYu0vutSp6eRVAJ3k0baC65aHH4/IrdlBkYIw6FBItqS+2+sEU04g29M7MGuVPgRx
wlbpR7aBkNDE1seivxYNE8Njorcfsm7YS0o20vLfL1pMH9h4NXfmlu9+0FHSBgOe5CozLuRHiWht
ROznF0R/dN8M3intQ0wlxlBA88TCYheTVgUUl6Bj93+nD5184FVgHfdXoryQ2nTYcx6xwZgDpFb9
msWKV7Vh75SdQSc9z64bvCtUEF7+oMWwUieK5Rb+Q6XT4QpUxy+T+H0le+yEKQJHNtpsHl0mvExs
gbDyCHuU6SUiCmrI56AEFzQvMxnSI0Yb2nrX/MUQum08NUVqS7og3XCAd5b895+huq8RQRMKF4Ad
VsiE7FN49L8UUS7Tt8NtyljO0whMI2PIx56VKpJwRzyLusq60R5cXtcfyQcvDJtQVD0d/X9vpmBp
tb/0c/mgd0XEjC+k1mWLh5LX6y3Rk3feZ2kucPdwKeIdNpyGlxOIRFzIh88xr/ASicLiaM/yd8kQ
d7qPL7H0ztKd9GatG/7CagabQ6+flJnn4vPTA7kj/v9skgdKd7ZJsKVhJvCG7yTh0D1ErckrckLS
HE8Rh1Q5CjVgfOqqHmACOX5Gwk9AMtoXDfrHyKGFNQ3qcPfTULDlhi1ow7DNu/N8kly7qXpfBoaB
ewqauYknAkwXKix/kLDJVM4S9IHGP9BG08fqaZI7aOqi8tA08oYVndjdGOjL0qH7i+u8pPrY9TqM
TdwP1haPI9ML4479+DIZURr6+PqOqgZH5WJoKOXWaBt6Ay8484Wj+jmHbgNPFP6tbrepd42fAtAv
Rfur4MNz9HBXIarzRJI1y80sezkyXaSw5Ms=
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw1n;
use gw1n.components.all;

entity PSRAM_Memory_Interface_HS_Top is
port(
  clk :  in std_logic;
  memory_clk :  in std_logic;
  pll_lock :  in std_logic;
  rst_n :  in std_logic;
  O_psram_ck :  out std_logic_vector(1 downto 0);
  O_psram_ck_n :  out std_logic_vector(1 downto 0);
  IO_psram_dq :  inout std_logic_vector(15 downto 0);
  IO_psram_rwds :  inout std_logic_vector(1 downto 0);
  O_psram_cs_n :  out std_logic_vector(1 downto 0);
  O_psram_reset_n :  out std_logic_vector(1 downto 0);
  wr_data :  in std_logic_vector(63 downto 0);
  rd_data :  out std_logic_vector(63 downto 0);
  rd_data_valid :  out std_logic;
  addr :  in std_logic_vector(20 downto 0);
  cmd :  in std_logic;
  cmd_en :  in std_logic;
  init_calib :  out std_logic;
  clk_out :  out std_logic;
  data_mask :  in std_logic_vector(7 downto 0));
end PSRAM_Memory_Interface_HS_Top;
architecture beh of PSRAM_Memory_Interface_HS_Top is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
  signal NN_0 : std_logic;
  signal NN_1 : std_logic;
component \~psram_top.PSRAM_Memory_Interface_HS_Top\
port(
  memory_clk: in std_logic;
  GND_0: in std_logic;
  rst_n: in std_logic;
  pll_lock: in std_logic;
  VCC_0: in std_logic;
  cmd: in std_logic;
  cmd_en: in std_logic;
  clk: in std_logic;
  wr_data : in std_logic_vector(63 downto 0);
  addr : in std_logic_vector(20 downto 0);
  data_mask : in std_logic_vector(7 downto 0);
  clk_out: out std_logic;
  rd_data_valid: out std_logic;
  init_calib: out std_logic;
  rd_data : out std_logic_vector(63 downto 0);
  O_psram_ck : out std_logic_vector(1 downto 0);
  O_psram_ck_n : out std_logic_vector(1 downto 0);
  O_psram_cs_n : out std_logic_vector(1 downto 0);
  O_psram_reset_n : out std_logic_vector(1 downto 1);
  IO_psram_dq : inout std_logic_vector(15 downto 0);
  IO_psram_rwds : inout std_logic_vector(1 downto 0));
end component;
begin
GND_s5: GND
port map (
  G => GND_0);
VCC_s4: VCC
port map (
  V => VCC_0);
GSR_30: GSR
port map (
  GSRI => VCC_0);
u_psram_top: \~psram_top.PSRAM_Memory_Interface_HS_Top\
port map(
  memory_clk => memory_clk,
  GND_0 => GND_0,
  rst_n => rst_n,
  pll_lock => pll_lock,
  VCC_0 => VCC_0,
  cmd => cmd,
  cmd_en => cmd_en,
  clk => clk,
  wr_data(63 downto 0) => wr_data(63 downto 0),
  addr(20 downto 0) => addr(20 downto 0),
  data_mask(7 downto 0) => data_mask(7 downto 0),
  clk_out => NN_0,
  rd_data_valid => rd_data_valid,
  init_calib => NN_1,
  rd_data(63 downto 0) => rd_data(63 downto 0),
  O_psram_ck(1 downto 0) => O_psram_ck(1 downto 0),
  O_psram_ck_n(1 downto 0) => O_psram_ck_n(1 downto 0),
  O_psram_cs_n(1 downto 0) => O_psram_cs_n(1 downto 0),
  O_psram_reset_n(1) => NN,
  IO_psram_dq(15 downto 0) => IO_psram_dq(15 downto 0),
  IO_psram_rwds(1 downto 0) => IO_psram_rwds(1 downto 0));
  O_psram_reset_n(0) <= NN;
  O_psram_reset_n(1) <= NN;
  clk_out <= NN_0;
  init_calib <= NN_1;
end beh;
