--Copyright (C)2014-2023 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--GOWIN Version: V1.9.8.11 Education
--Part Number: GW1NR-LV9QN88PC6/I5
--Device: GW1NR-9
--Device Version: C
--Created Time: Thu Jun 22 22:32:13 2023

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(12 downto 0)
    );
end Gowin_pROM;

architecture Behavioral of Gowin_pROM is

    signal prom_inst_0_dout_w: std_logic_vector(29 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(29 downto 0);
    signal prom_inst_2_dout_w: std_logic_vector(29 downto 0);
    signal prom_inst_3_dout_w: std_logic_vector(29 downto 0);
    signal gw_gnd: std_logic;
    signal prom_inst_0_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_2_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_2_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_3_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_3_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 9;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    gw_gnd <= '0';

    prom_inst_0_AD_i <= ad(12 downto 0) & gw_gnd;
    dout(1 downto 0) <= prom_inst_0_DO_o(1 downto 0) ;
    prom_inst_0_dout_w(29 downto 0) <= prom_inst_0_DO_o(31 downto 2) ;
    prom_inst_1_AD_i <= ad(12 downto 0) & gw_gnd;
    dout(3 downto 2) <= prom_inst_1_DO_o(1 downto 0) ;
    prom_inst_1_dout_w(29 downto 0) <= prom_inst_1_DO_o(31 downto 2) ;
    prom_inst_2_AD_i <= ad(12 downto 0) & gw_gnd;
    dout(5 downto 4) <= prom_inst_2_DO_o(1 downto 0) ;
    prom_inst_2_dout_w(29 downto 0) <= prom_inst_2_DO_o(31 downto 2) ;
    prom_inst_3_AD_i <= ad(12 downto 0) & gw_gnd;
    dout(7 downto 6) <= prom_inst_3_DO_o(1 downto 0) ;
    prom_inst_3_dout_w(29 downto 0) <= prom_inst_3_DO_o(31 downto 2) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"955595555656A599A9555565555599666655955956556AAAAA5555546CB9B1EE",
            INIT_RAM_01 => X"ED3FAAAAAA555559555566A6A9967D5659F5596696659A5995555655555A99A6",
            INIT_RAM_02 => X"F0000C0030003C000D557C0030000C000FFFF000055550000CC00C0002BB4FC6",
            INIT_RAM_03 => X"00000000000000000000000000000000000000000FFFF0000001800002400FFF",
            INIT_RAM_04 => X"A7AFFFE00AE00FFFF00030033FFFFFFFFFFFFC003D557BF8000A02BE80000600",
            INIT_RAM_05 => X"01FFF0000FFF4000B03FFE000FFC000000FFF0000FFF000000FFF0000FFF0000",
            INIT_RAM_06 => X"00FFF0000FFF0CAAACBFDAA00AA7C00000FFC00003FF0000008020000F7B4020",
            INIT_RAM_07 => X"215088000205400000FFD0000000000000FFF0000000000000FFF00008000000",
            INIT_RAM_08 => X"C0A8008000A801A900A801A900A801A900000000000000000000000000000000",
            INIT_RAM_09 => X"000000FFD000000007FF0000000000FF4000000001FF00000C2AAC7FDAA00827",
            INIT_RAM_0A => X"00FFE00000000BFF0000000AF03F00000FA000FC0000003FF005F0000FFC0F50",
            INIT_RAM_0B => X"03FF00000000003FF005F0000FFC0F500000000AC03FF00003A00FFC00000000",
            INIT_RAM_0C => X"0000000FF0000EAAA0000000000000FFE000080000000000000000FFC0000000",
            INIT_RAM_0D => X"0000000020000BFF0000000000000FFEA000000000000000F0000FFFF0000F00",
            INIT_RAM_0E => X"F000000000000000F0000FFFF0000F000000000000000AAAB0000FF000000000",
            INIT_RAM_0F => X"0000002FE0055000041BC55000AAA0BFD0000AA00AA7C0000000000000000ABF",
            INIT_RAM_10 => X"A0BFD0000AA00827C000001FF01FC000055E0D730000002FC02FF0000FF30AAD",
            INIT_RAM_11 => X"000BC5500000002FC02FF0000EB30AAD0000002FF02FC000055E0FF3000000AA",
            INIT_RAM_12 => X"000AA00BFAAA0DAA70000C0000AAA0BFDAA00AA7C00000000000002FE0055000",
            INIT_RAM_13 => X"00AAA0BFDAA00AA7C00000000AAAABFDAA000A7C0000A000BAAAAFDAA00007C0",
            INIT_RAM_14 => X"70000C000000A000BAAAAFDAA00007C0000000000AAAABFDAA000A7C00000000",
            INIT_RAM_15 => X"C4CF1B8D38F38CCCF3931C6C713B33CE2738F3309C313C2CB00AA00BFAAA0DAA",
            INIT_RAM_16 => X"70CE31C6AC70ECEF3C3BCF3ECCE38D38E330F0FB318C6B1BF87CE73C71736B33",
            INIT_RAM_17 => X"92567440B65E51D1674E10518508E34DEFA13333CC68A31A28CCCF71C33072F2",
            INIT_RAM_18 => X"218125D298D144CB27640AC918306C18036665645499431844B6754576547564",
            INIT_RAM_19 => X"015CC763B101E4CC18F6250106401F94079330E3D89405725406585391913147",
            INIT_RAM_1A => X"727667796255DC251135605437148A3043425148A34965509333D0198B18F635",
            INIT_RAM_1B => X"D1D19155192247CE3476544406811041464607041A0741913445914504162552",
            INIT_RAM_1C => X"506D0C825308E11541B4130D0714574702D1E1560B2430080674766456466015",
            INIT_RAM_1D => X"066CD991F289D9D51115DD19D1DD1B0AC151D19DD924564544456705D4F23C45",
            INIT_RAM_1E => X"D9E300E3051C157055015597478CD191DD5DD19915530BC1270D9955119E34F3",
            INIT_RAM_1F => X"F1804448AC511D289D087737C8875419DA300676728C019D9050005765004011",
            INIT_RAM_20 => X"76679573DD13DD41F4010005C37674A145170517179C55D0D3615743494552C2",
            INIT_RAM_21 => X"5244D09134100C89AC81A8EE0D9936640DDA7754D516441511B2350240D06777",
            INIT_RAM_22 => X"180476566749C3476707299111070544380C0320C0CCD03010743000D0F79D71",
            INIT_RAM_23 => X"75C760731B142451A7A155A452B00AA15469AA2A69A068506273446899115595",
            INIT_RAM_24 => X"C274246375447437666A1D591DAF24A1774666A95599D1D15525441C500DD3DE",
            INIT_RAM_25 => X"0544362635598C5951138D5E6C514D01A2455C98D40668B122300247A8770991",
            INIT_RAM_26 => X"92261147CC14720A0702A28A2029A717A49032132016434685C8115618560A3A",
            INIT_RAM_27 => X"D11844483C15515A3547744499D1D2483777665CB0149282B96605BA00B8C04C",
            INIT_RAM_28 => X"47048A355148A3208403138410D09C5200E08A344075716151655043689581C9",
            INIT_RAM_29 => X"5155455640505551DA05A205565D1417481D10B48355D4D08C9F39D344CF38A3",
            INIT_RAM_2A => X"9415C9E85F79D719F061520626B76453DE675C76278C12347FC520528A1DE550",
            INIT_RAM_2B => X"15A2567790C213744E9343474D1914CD11EE8D3DE75C59C3CCC8098804583059",
            INIT_RAM_2C => X"55119D7443A286821444451153664564674344881005774481681E943E68372D",
            INIT_RAM_2D => X"230C0D0307545444422022440828EB2091029024893409249A228D041D356441",
            INIT_RAM_2E => X"76756499276C3C995E382F1686AA0DD95C0460D25D19D0D234342864648D0300",
            INIT_RAM_2F => X"10100F1764646089D059811DB174648149130C230C0100AABC50EDD9DB1B1147",
            INIT_RAM_30 => X"2C8D1CCA00655745640F9B01741D19049C0A00050048030011764676089D0D94",
            INIT_RAM_31 => X"832065574464091E89526C2C0D1CC107320823A2564B0B03473061CCA30648B0",
            INIT_RAM_32 => X"19900247A2664B0B03473061CC8014B0B02C8B03473041CC8200654B22C0D1CC",
            INIT_RAM_33 => X"B0B0347304732883A2564B22C0D1CC11CC8120E89992C0B234C102841901955D",
            INIT_RAM_34 => X"73047320883A2564B22C0D1CC11CC8120B02C8D1CC11CC802065065574464091",
            INIT_RAM_35 => X"91D112715264D5926C35493607040770E3070C1E335374190A25495091B0B034",
            INIT_RAM_36 => X"3624144D8614A53C014A534810A53C01CA5348D8905183745C983641C5C03C4D",
            INIT_RAM_37 => X"519C34B081804444B56456454A3BCCDD534DDE82868ADD115592861460060062",
            INIT_RAM_38 => X"1DD74775D8141D0DE850005801005001D8D519748263814D1D9192475464499D",
            INIT_RAM_39 => X"19191F20B366455445282C9D2C9D04106D59151158057476645544414444775D",
            INIT_RAM_3A => X"1D15410C18551D0235505106095D580003AA43169651926015D15D19D591D10D",
            INIT_RAM_3B => X"D0935057424995064416C1116B23691501A4015AB2895D591174677774340444",
            INIT_RAM_3C => X"0129505E5976029879D4074A134A88A4262090850701888741C101C040DAC815",
            INIT_RAM_3D => X"2372945444DD2655628159593404A06A01474464824ED019D01D222784106041",
            INIT_RAM_3E => X"32A681474701F3CF7CC7F14DF44FF3CF7CC7F1000A0695510790244A11111CAB",
            INIT_RAM_3F => X"30D2AB33030310812E00DE25444D95120A6348218D20A91D04A91D07082E9A1B"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_0_AD_i
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"40004000010150445400001000004411110040040100155555000002FCA30089",
            INIT_RAM_01 => X"4555555555000004000011515441140104500411411045044000010000054451",
            INIT_RAM_02 => X"00000C0000003C000C003C0030000C000C000000055550000CC0000000115540",
            INIT_RAM_03 => X"90A200A2000280A000A082EA80A20202000000AA0FFFF0000000100004000000",
            INIT_RAM_04 => X"F1FEBFFC0FF800003000300330000C0000003C003C003FFC00FFFBFFE0000060",
            INIT_RAM_05 => X"A0FFFAA00FFD0003F01FFFC00FF40000A01FFA000FF40000A01FFA000FF4000B",
            INIT_RAM_06 => X"F03FFFA00FFC0C1FFC1FC55E0D73000AF03F0FA000FC000001FAF0BE0400003E",
            INIT_RAM_07 => X"30090C0900600008003D00000000000AF03FF0000000000AF03FFFA00FE8000A",
            INIT_RAM_08 => X"01A901B903030088030302AA0303020801A5809542558300C157417602708060",
            INIT_RAM_09 => X"000000FFC000000003FF0000000AF03D00000FA0007C00000C2FFC2FC55E0FF3",
            INIT_RAM_0A => X"003FF00000200FFC0000003FF00500000FFC0050000000FFF00000000FFF0000",
            INIT_RAM_0B => X"03FF0000000000FFF00000000FFF00000000003FC005F00003FC0F5000000008",
            INIT_RAM_0C => X"0000A003FFFA0FFFC0000000000AF03FFFA00FE800000000000000FFC0000000",
            INIT_RAM_0D => X"000AF02BFFA00FFC0000000000AFF3FFFA000FC0000000003AFFAFFFF0000C00",
            INIT_RAM_0E => X"C0000000000000003AFFAFFFF0000C000000000000AFF3FFFA000FC000000000",
            INIT_RAM_0F => X"002AA07FD0000AA00AA7C000001FF01FC000055E0D7300000000A003FFFA0FFF",
            INIT_RAM_10 => X"F01FC000055E0FF3000000BFC0BFF0000FF30AAD0000007FE0555000041BC550",
            INIT_RAM_11 => X"0827C0000000007FE0555000055BC5500000007FC07FF0000EB30AAD0000001F",
            INIT_RAM_12 => X"0001F001FF55ECFA30000000001FF01FC55E0FA300000000002AA07FD0000AA0",
            INIT_RAM_13 => X"001FF01FC55E0AF30000000001FF51FCF5E00A30000010001FF55FCFAE000300",
            INIT_RAM_14 => X"30000000000010001FF55FCAFE0003000000000001FF51FCA5E00F3000000000",
            INIT_RAM_15 => X"4A4120951041051405290454129051043D104052F48076555001F001FF55ECAF",
            INIT_RAM_16 => X"5114514614514141049141041441051040524220912485209450451851516090",
            INIT_RAM_17 => X"F37444A897B055123FAE18E30F2AC105F414545014830920C241445950515040",
            INIT_RAM_18 => X"B7863303F861CBF503A489400430AC040068686878364B3CC804786584476494",
            INIT_RAM_19 => X"C1C414417BC1720D140437C03573E8CF05C8341010FF07106303B860E2040A08",
            INIT_RAM_1A => X"80786940CF77ED3F2D28828A28738532B1B1819473C7DB2104373C124304043B",
            INIT_RAM_1B => X"5A1612121EF07B8C1477474831011AC914080B000404A15A84251001865CFB2C",
            INIT_RAM_1C => X"909F30CE63CCD10A427CE32D0866B74981D111F9841C71862496858684859892",
            INIT_RAM_1D => X"1A781952C1852D69E9A1DE1D21D527010D1691E5EF079694454A798998D33C42",
            INIT_RAM_1E => X"9EFC2CFD083C60D283820C30CBF029515D11D11DD51C37F007C1E1E1212D37D1",
            INIT_RAM_1F => X"FC50486C901D1998D60A49150CA48A95271435A7B24C0D69E0A0035A782800D6",
            INIT_RAM_20 => X"4747751336033646CC82200AD0784B434AB74D21177C22E4EB708B92ADCD31C0",
            INIT_RAM_21 => X"281A6A06B42A0B46DDCAD4DE0BDF37580508AF07D5A7569919C37727C9D85757",
            INIT_RAM_22 => X"6F3655556942D04B49252DD252D8048616B0CC1300C42AC030965438905D75D7",
            INIT_RAM_23 => X"F7DD8710353524D33D30A64490412101594B1305479C1414D0C048D0DD29A9ED",
            INIT_RAM_24 => X"0879079044486A14546A1D15959A2490454456A551D959D1D5956B205AA9E3BE",
            INIT_RAM_25 => X"048714150845F09DDD29CD1D18210D01D1C2D0D0188004430282100004492000",
            INIT_RAM_26 => X"242BA188301A7D2A8E1122A600A51F043CF255545427834BC28F10A5266B2415",
            INIT_RAM_27 => X"F31555AE145565AF186A744A9D96E3C71747475FE28CF0CA87580A462A8604C1",
            INIT_RAM_28 => X"4905CDC4905CDC46DDB6423CA4686C6518C1CDC490667070B06640407799C181",
            INIT_RAM_29 => X"A083820FC81820C3E706710830C32DC4B712227009E2F92980053F6049CE30DC",
            INIT_RAM_2A => X"14698110D7DF6DB65381A1091567A6B3FFEBBED82630A504BFC6A092471B012C",
            INIT_RAM_2B => X"B742B478740D10740D5343EB4D6F1F0295440CDB6D75D6D149C94E089A68B4D2",
            INIT_RAM_2C => X"0C383E0CA040410104848121E07848686B73E88A00249788A3922555403F285A",
            INIT_RAM_2D => X"294627030946844860A228000C90551000094F104418008207D1C60425058682",
            INIT_RAM_2E => X"49496029057D14E92717D52AB66429E92D349C6C1E1E7E711C9C143414A43180",
            INIT_RAM_2F => X"2BF2C6D479459C0E1821422581454688A835C711C70344A6542CD9E9E055A265",
            INIT_RAM_30 => X"2409270B20945844860F4B4846A1119A19C92F4A208ABC289D479479C0E18218",
            INIT_RAM_31 => X"8020945844862521016864A4092700C9C2048C404869293249C01270B2096392",
            INIT_RAM_32 => X"16188948405869290249C032708223929324490249C022708030963912409270",
            INIT_RAM_33 => X"9293249C029C2C8C405869124092700A70802310161A4890248082C425825161",
            INIT_RAM_34 => X"9C029C200BC404869124092700A70832F9224092700A70830095094584486252",
            INIT_RAM_35 => X"2DA013537366DD5B6024B2C9090809638C0A7029C140B40608C1042252929024",
            INIT_RAM_36 => X"0A090B459928CD20C28CD2C828CD24824CD20820242DBF4B20DBF4B20DAC2049",
            INIT_RAM_37 => X"5E1C84700050486C85454646663500D22B42550949895599999A7F2BF2BF2FF0",
            INIT_RAM_38 => X"1F27C7C9F02C25455040884082444C825829251A60915105A1521978548775E1",
            INIT_RAM_39 => X"2129ADD8405848684924140E940D0A00C1A1212126249787878487A048487C9F",
            INIT_RAM_3A => X"3A5EA5105821D64D2FEDD64D851E148442C608045681515B925E1A16121E9AC1",
            INIT_RAM_3B => X"E49B418B916D9595561515115C154405057C195A84455111104447EAF3B03D49",
            INIT_RAM_3C => X"012954505614229EC05084AA18AA08591A11EA0514015404B202428884111062",
            INIT_RAM_3D => X"03845486486E1884AA802094D800C29C0068448673F9E0FEE0F9222C08081020",
            INIT_RAM_3E => X"1319C00E8944F3C53C41700E0083C3C53C41710289C992923F603E891251111C",
            INIT_RAM_3F => X"7C12A9320300208B2C029104448DDD222F9188B24612106D0A106E8002111C65"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_1_AD_i
        );

    prom_inst_2: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"9595555655569996A555559555566665995595655655AAAAAA555556E7700CB8",
            INIT_RAM_01 => X"B4FCAAAAA955556555559AA6A655765955D9665A6599699655555955556A699A",
            INIT_RAM_02 => X"00000C0000003C000C003C0030000C000C000AAAA00000000CC000000AED3F2B",
            INIT_RAM_03 => X"030CC30CC024C30CC30CC0C9030CC324C3AA8324CFFFF0002000080000000000",
            INIT_RAM_04 => X"7007FAF40AFC00003000300330000C0000003C003C00315003FFF7FFDC0006B5",
            INIT_RAM_05 => X"F03D5FFE0550002FF007FFF80FD0002FF0005FF80500002FF0005FF8050000BD",
            INIT_RAM_06 => X"F005FFFC0F500CBFCCBFFFF30AAD003FF0040FFC00100000003F43C1C00000FF",
            INIT_RAM_07 => X"009030900C06003E000400000000003FF005F0000000003FF005FFD40F50003F",
            INIT_RAM_08 => X"00A802AA00540333005400E4005403930030C1800300C30CC00600324300C006",
            INIT_RAM_09 => X"000AF03FC0000FA003FC0000003FF00400000FFC001000000C7FCC7FFEB30AAD",
            INIT_RAM_0A => X"0005F00000BC0F50000000FFD000000007FF0000000000FFF00000000FFF0000",
            INIT_RAM_0B => X"0FFC0000000000FFF00000000FFF0000000000FFC000000003FF00000000003E",
            INIT_RAM_0C => X"0003F0005FFFCFF500000000003FF005FFD40F5000000000000A003FF00000A0",
            INIT_RAM_0D => X"0017F005FFFC0F500000000003FFF05FFFC00500000030000FFFF5FF5C000000",
            INIT_RAM_0E => X"00000000000030000FFFF5FF5C0000000000000003FFF05FFFC0050000000000",
            INIT_RAM_0F => X"002FF02FC000055E0D73000000BFC0BFF0000FF30AAD00000003F0005FFFCFF5",
            INIT_RAM_10 => X"C0BFF0000EB30AAD0000001FE0155000041BC550002AA02FD0000AA00AA7C000",
            INIT_RAM_11 => X"0FF30000002AA02FD0000AA00827C0000000002FE0055000055BC550000000BF",
            INIT_RAM_12 => X"000BF00BFCF53FAAD000000000BFC0BFFF530AAD00000000002FF02FC000055E",
            INIT_RAM_13 => X"00BFC0BFF5F30AAD000000000BFCFBFFA5300AD00000B000BFCF5FFAA3000D00",
            INIT_RAM_14 => X"D00000000000B000BFC5FFFAA3000D00000000000BFC5BFFAF300AD000000000",
            INIT_RAM_15 => X"000000000000000040800000000800000000000000044041000BF00BFC5F3FAA",
            INIT_RAM_16 => X"0002000000002000000000000000000000000000000000000000000000000000",
            INIT_RAM_17 => X"C912209D2772CCC253BCA6FB6C97E0A151450401000000000000000000000000",
            INIT_RAM_18 => X"9222000562243ACE878BD3A13E84A73E881838281906D91468803A00A21110BE",
            INIT_RAM_19 => X"2002511B1E200021B2515E2381080168800086C945588009106D22200844BFE8",
            INIT_RAM_1A => X"8E328000A112BD98C41484091EA47D940C3C1C32EBA610214585620424B2515E",
            INIT_RAM_1B => X"4606020A02EB1B2C8033320822102D92684840CC8840928E40C80320828A10EB",
            INIT_RAM_1C => X"E7CEB692AFABF8CB9F3AC9542EB0820BA94BA43BEEBEFBEF909381808282BE42",
            INIT_RAM_1D => X"43B60CC2DB64A42CECA0060068482CBB280A806CEDB1B083120B0BA8ABFAFE32",
            INIT_RAM_1E => X"86B076B1C9AB258C967659850AC30A8A86042042C2D0F3C86B20602020EFA88B",
            INIT_RAM_1F => X"A0B43893320A0AB6421A084321A089A4AEA3A2A18F21A8A86BFA5A2A1BFAF28A",
            INIT_RAM_20 => X"18194AF942C942145BA2E8BFD8181A863F6B602FA16302C3ED9C0B0EB6B2CB2E",
            INIT_RAM_21 => X"205928167EE190942090032D902C8019D0034EB4467919ECACF8886B2A662928",
            INIT_RAM_22 => X"6EB000030B3FD80A0BEB48A602B8C009E9FAAE9BA23D04E886AA20BEFA514514",
            INIT_RAM_23 => X"1450B8F840CB45559C8488A3A614A6C919336C9133C51339D2EB0AA18A6C6C2C",
            INIT_RAM_24 => X"2428428680082B9595A0529ADA2FBA0811C11E088B438F07DA4E0A2136CFA986",
            INIT_RAM_25 => X"5018FAFA4AABC1A8882724AEA10E5E5AEA50A9E5AD04C008F41C4C4C883B4133",
            INIT_RAM_26 => X"2207B04BC10CD3401E88A4ADBA04CC4CB6C8000030B0BE0BA2DE8CB9F3187171",
            INIT_RAM_27 => X"EA40089DBA2020AF8938090902CAEB2CA19090B4DA72EB203A18500B4A001032",
            INIT_RAM_28 => X"08EB6B209EB6B00044110AC90303030CBECB6B208EA28E84AEA29E96AC8ABA1A",
            INIT_RAM_29 => X"B49AF26B27652698AEA2E86966142C20BC82B43ED112477020003F2E0BECB2B2",
            INIT_RAM_2A => X"1F0AD3A5271C6182E88684C0C8818295C70986097AC10CB0BDA248B43EB72428",
            INIT_RAM_2B => X"9DCC1C7AB23F86BAD8FBA41BA82CB830A000081861453FDBA060663D0923360E",
            INIT_RAM_2C => X"69898E508884A2128083A020A81808183B840AD0129093AD024A2000002C16B3",
            INIT_RAM_2D => X"ABAD8C886A938908920B404CA94D4EBA1326E2BA6E88A5145D1B6225AA8181A2",
            INIT_RAM_2E => X"08080120EB3DBA60ACB02E880801C060AD80BA2A0602C0C9B23299585AAEAB62",
            INIT_RAM_2F => X"4F2F6F111910B25465C690EAC9191820918BEF9BEF882D08BAA3606025555800",
            INIT_RAM_30 => X"B62FBC1D96A909909B0F4B54137604DD6ABCBCFF862AF0FAE111912B25465069",
            INIT_RAM_31 => X"E896A909909B98261465B6362FBC15AF07A6E10D09BD8DABEF055BC1DA5AB8D9",
            INIT_RAM_32 => X"466EE61985199D8D8BEF056BC1E9BCD8DAB66D8BEF055BC1E8AF2BCD9B62FBC1",
            INIT_RAM_33 => X"D8DABEF054F076C10D19BD9B62FBC153C1E8B043466F66D8BE752F6B4A5AA426",
            INIT_RAM_34 => X"F054F07A2C185099D9B62FBC153C1EAB0D9B62FBC153C1EAA5A96A909909B98A",
            INIT_RAM_35 => X"08DA5E2E9E1F687DB2A0A288E0D1FAB8D063014F06BC0A522D16ED298ED8D8BE",
            INIT_RAM_36 => X"C0C1C2A888EA6DB61AA6DB256A6DB2B2A6DB2B070B0AF20A21AF20A21AE3FEF8",
            INIT_RAM_37 => X"8A61EACBB4B4389301818282AD8B210224A2AA1A1A1A8A8A8AA70DBCDB8DB4D9",
            INIT_RAM_38 => X"9C07A5016743CAB221B213B21457BA1CA10AA24A860686ECE6C26609A29B4826",
            INIT_RAM_39 => X"6028283EE81808180A4EBA12BA1FB832E06020A06F90908182818084180A601A",
            INIT_RAM_3A => X"710CD227252AC21C433EC65C7ECCE163A43018FBB0A727BC4242060A06028210",
            INIT_RAM_3B => X"C37D9C0B0DF6567D59FA6DADAF9DD94D5EB27F881128A4242818180005724008",
            INIT_RAM_3C => X"2B41A3328200B41EC8CAA090A090D29852886CA490E110A0A238343BA2E6C302",
            INIT_RAM_3D => X"999104A76856158488A5252E08B2D82D89399099CB0CE906E90EB4448A515945",
            INIT_RAM_3E => X"858B228545452001A0482141B4483001A0482A40D4D44A4243F240AE52DAD66F",
            INIT_RAM_3F => X"0208027A5A4B5AD34E6A7AB330A8882B4448AD1122A4006FBA00620C8900066D"
        )
        port map (
            DO => prom_inst_2_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_2_AD_i
        );

    prom_inst_3: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"404000010001444150000040000111104400401001005555550000023463F1BB",
            INIT_RAM_01 => X"1554555554000010000045515100110400441105104414410000040000151445",
            INIT_RAM_02 => X"0FFFFC0030003C000C003EAAB0000FFFFC000AAAA0000C000CC0000000455501",
            INIT_RAM_03 => X"010641A64240C1AE418EC0D001824342410101EA4FFFF0024000018000000000",
            INIT_RAM_04 => X"F0001FD00FD000003FFFF0033FFFFFFFFFFFFC003EAAB0000055F17D40000000",
            INIT_RAM_05 => X"F0100FFF8000003FF0007FFC0D0000FFF0000FFF000000FFF0000FFF00000BFF",
            INIT_RAM_06 => X"F0000FFF00000C1FEC15541BC55000FFF0000FFF00000000007402C0C00002FF",
            INIT_RAM_07 => X"4000110A840000FFE0000000000000FFF0000000000000FFF0000400000000FF",
            INIT_RAM_08 => X"01A90000025600440256004002560104015540154055015541554154005502A0",
            INIT_RAM_09 => X"003FF005C0000FFC0350000000FFD000000007FF000000000C2FEC05555BC550",
            INIT_RAM_0A => X"8000000002FF0000000000FFC000000003FF0000000AF03FF0000FA00FFC0000",
            INIT_RAM_0B => X"0F500000000AF03FF0000FA00FFC0000000000FFE00000000BFF0000000000FF",
            INIT_RAM_0C => X"000FF0000D5550000000000000FFD0000400000000000000003F0005F00000FC",
            INIT_RAM_0D => X"0000100007FF0000000000000FFD5000000000000000F0000FFFF0000F000000",
            INIT_RAM_0E => X"000000000000F0000FFFF0000F00000000000000055570000FF0000000000000",
            INIT_RAM_0F => X"007FC07FF0000FF30AAD0000001FE0155000041BC550000000000000057FF000",
            INIT_RAM_10 => X"E0155000055BC55000AAA0BFD0000AA00AA7C000007FF07FC000055E0D730000",
            INIT_RAM_11 => X"0AAD0000007FF07FC000055E0FF30000002AA07FD0000AA00827C0000000001F",
            INIT_RAM_12 => X"0001F0015E55B5550C000000001FE015555BC55000000000007FC07FF0000EB3",
            INIT_RAM_13 => X"001FE015555BC5500000000001FE515555BC0500000010001FE555555BC00000",
            INIT_RAM_14 => X"0C000000000010001FE555555BC000000000000001FE515555BC050000000000",
            INIT_RAM_15 => X"AAAEA4A0820820A82AAABAAAEAAAA820AA820AA0A82820082001F0015E55B555",
            INIT_RAM_16 => X"E0AAEBA82AEBAA0EBAC3AEB0AA0820820AA000A4AAEABAA482C20E82E0E824AB",
            INIT_RAM_17 => X"A19998BCEA622222899E30F34E39E2A0A09282A0AA924AA492AAA0C30AA0E000",
            INIT_RAM_18 => X"068215542828BA19092FFE42290E23290888B8A8AA2AFC2088BBBAA8AAA998A0",
            INIT_RAM_19 => X"815455504281554504554E801551553A05551411552A05515540A82151550001",
            INIT_RAM_1A => X"8DB58000859A6B0E06188CC419ADF83ECECECEEC92CBAA215514A81545045546",
            INIT_RAM_1B => X"6222222A22A1BACB2A999988132212FEA89C9CC88C8842A508BA222249A84A20",
            INIT_RAM_1C => X"637B28A5BE8F90C18DECA0E61998AA8A076668BA8820A28A189988888A88A862",
            INIT_RAM_1D => X"CDACA66282C6222A2A22222262222B0A822A22A6E91B98B9A9898A066FA3E430",
            INIT_RAM_1E => X"2AA4A4A4E223089C22308A288A9332222222222226A4CE54DA82222222292183",
            INIT_RAM_1F => X"B4F88483E82222EC223888AAC388042629088A8B8A0322A22290C8A898AC322A",
            INIT_RAM_20 => X"88886AB062B062331AC2B0AAB08899C9A91ACA2B286631D23298C748CA7A82C2",
            INIT_RAM_21 => X"2C8407212CC762FFBAFFB3AB22AA2AB9000016E9A92AA4AAAA8088CA022C8888",
            INIT_RAM_22 => X"291BBBB989AAB28A88DBF652EE28E868D8E0280A023F3B808C0998A0B19A69A6",
            INIT_RAM_23 => X"8618A5B0ECEB3081888C3BE88EFCFA9189A2A829A27373633281897265662626",
            INIT_RAM_24 => X"2088C88D88889B4888A2662222AA28A488888A2222262266291A8823EE500461",
            INIT_RAM_25 => X"E868D9D9C2AE9366662E866773323636773323636F888CC8FFC88CC88C8BE212",
            INIT_RAM_26 => X"2A1A638A933A87EF3A08B39B206688D8A4A3BBBA98988E8A42390C18DD89DDDD",
            INIT_RAM_27 => X"B3EEA48A28AA2A6908948884226EB28A088888A1B1E0A206D988CEAFEF2E333A",
            INIT_RAM_28 => X"88DA88588DA887BA66998ADFB3B3B3BB28B288588D999D8CBD999D8DA1663636",
            INIT_RAM_29 => X"BC22F08A83A308A2E91A90C228A22858AD627EECFA220AAA2AA0952D8A8B2C85",
            INIT_RAM_2A => X"E2760E63A8A28A22A28D8CECEAC8888C20882088DAD3BB189BD925B339222A20",
            INIT_RAM_2B => X"99CCDBB9A03B0DACF782C88AC62A2133200008669A69AAB28222623F8463ACA2",
            INIT_RAM_2C => X"8A262E8A94CCD3334888922224888888BAD889FF22589B9FF08A2000002119A2",
            INIT_RAM_2D => X"66083808C08948848267FC889F7F79242227A4A82A0892CB2A4A822302488898",
            INIT_RAM_2E => X"8585A338DAAB2822EA253A1408CCE222EB08A022222E8780A0E05C8899980A02",
            INIT_RAM_2F => X"384A4B48888BA83323B233C2B088899C424A8A0A8A089FCCE8636222E0000599",
            INIT_RAM_30 => X"A82B253A0C088C88C80F0FE08A5222942AE821E90CD984AC848888AA83323F23",
            INIT_RAM_31 => X"A08C088C88C842232210A8E82B2533294E82B4C88C8A3A0AC94CCA53A0C0ADA0",
            INIT_RAM_32 => X"23211088C8848A3A0AC94CCA53A0A5A3A0A82A0AC94CCA53A08CCA5A0A82B253",
            INIT_RAM_33 => X"A3A0AC94CF94E884C88C8A0A82B2533E53A0A132232282A0ACF3FE8332702232",
            INIT_RAM_34 => X"94CF94E86A4C8848A0A82B2533E53A0A9A0A82B2533E53A08C09C088C88C8422",
            INIT_RAM_35 => X"1AA08ACE8EACAAB2AC688208CCCCF0A594CE53384C8CD9322A49922422A3A0AC",
            INIT_RAM_36 => X"CCCCCE92222AEA2832A2A2832A6A2832AAA28333333AB64820AB64820A87A4FB",
            INIT_RAM_37 => X"632319B0BCF88483C9898888BB1AC3601190AB3B3B3BA9A9A9A21A25A2DA25A0",
            INIT_RAM_38 => X"420090802333323AB36233623333623326365D89CCCDCD925221218C9ACA1632",
            INIT_RAM_39 => X"2226A86880A888888BF92420642B3122E22222A22A189A8888888A8C88890802",
            INIT_RAM_3A => X"EBEA4EA3E30A62378AA66237366D63F3F89B3CD9988DCDA9626A2222222A6A32",
            INIT_RAM_3B => X"D2B288C74ACAA92AA4AAAAAAA808A8D8DAA062A9AA92222224888BFFFEF18B88",
            INIT_RAM_3C => X"2736A3E2A20073698AD96840A440FECC8C8A309A688EA8A48233333B296A6231",
            INIT_RAM_3D => X"08AAB88888220898489222AA48ACB3BB08948848A297B223B2267388892C88B2",
            INIT_RAM_3E => X"0C8A43CFCFCFE3CBECCEA3CBECCEA3CBECCEA7DFF7F762628A22889762AAAAA8",
            INIT_RAM_3F => X"145557FBFBEBE9FBFE26664888922227E0889F82227E321B3132104888322229"
        )
        port map (
            DO => prom_inst_3_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_3_AD_i
        );

end Behavioral; --Gowin_pROM
