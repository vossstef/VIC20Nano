--
--Written by GowinSynthesis
--Tool Version "V1.9.10"
--Wed Aug 14 14:08:55 2024

--Source file index table:
--file0 "\/home/vossstef/Gowin_V1.9.10_linux/IDE/ipcore/PSRAM_HS/data/PSRAM_TOP.v"
--file1 "\/home/vossstef/Gowin_V1.9.10_linux/IDE/ipcore/PSRAM_HS/data/psram_code.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
Of+y9LO6mD0nYLoRz912qVNOlLfUNFhIzZkDj3sxuQ+rtLICiuZaHaT26xfZ4EoosTbJPeWw+mDI
tDd4rhBePJN6Pfd6qavwjgux2ujz4zBu3kWcq8udp8c+KJTpEgwfFDasEPDqEjqk34dcVRVBuBsj
zMBnC8nnviCjoHuwJpFIG0J19m8ORnNhCOvQC8/v0d/oJFkIQ9grhShQuuYWPeFdCbNxFrQsXl12
Co+0KWkfqXIHW9wEEPW/pG7cHDq7qgv/Mn22aoIwCYVP3X7/AuXK6IZZ8eftCJtotXsLbLJevcTV
qIM0qz1CEL6/a3bwxsmYQYfGh9fTDGIotZ68Gg==

`protect encoding=(enctype="base64", line_length=76, bytes=310448)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
cGT2Pgjf6Wnl8vycK0TpFQsAslEGr9Pv9tkw1k1Rzr2w+TIfsfagABQwD/QWqYaXVrCW5nnG8A77
qZVQeaBzcx0+QQkMKqof25TwJs8py7qKgutKbT6XXaZcYHdD/UFTA9kFmjyqY6Xdy23t0LTgQH/G
QSAJH6m/zMSgD738VLaJkT+gXeB/JD3OgvpvmGyxqw4Hd2xnyr9cTOxCfMHxukCUnVGLvVwN+vBV
wKSKZ76Oui/X48QBHZetnKGXBugfay7L7DkjNlMJ//msbDChDxt4navqMG1HafKsuEl54D5b5ech
/gCuUxirZwsP55yumTH1tjrjitVseydsTDfu9Yk6zaVeNjEHHnVDo0CLXl/BxbFvf7psgPAGDV4a
wwyPOlOLtcwNc9K6ZiwZw6gEOFa909pPqYADR0OXXzLj+cgBTZaQYvBUteuR8WHhZJhFkmGM/vk1
Qbhh9ieJnebKlykiKP9KmLJUA297+DJ4GkEWf9RJTxPe3RBwgeib48RLVtMBwq+X9OA3sZ5Wr96W
vu977N2xFF5iI5zezIauwAo6t33Jx/j1kJ09mMBYe4lTuxZcR32HCPiArFSztoiuWoOT4ScaK6nv
UYMQT+N1KsLg9bcKK3hwKmQxrgOHp6RCoU8ml+ItbJG2TWrnIwzEixSHdpEul+Jo4jr3AxhoJ8CZ
2G6zlkx4HHJuEO0b1Q8Sro+LCUf9LYoOzY7Z8O8Elx4GejDfsh+Wy32c2UxE3rf4VnDSh2srky7s
1dsIoTxHqilE24UMtS/ZVLmmdYkRRpd2BeM9gUJCl8L3jh/oxTxVGkd/SSysMqvm7cHrzJKm87bg
C+J23v/Ej9W3Jc/s6sgXj0gBsGHDeguU8d8wU+J3rG00LR6IflhasYYUBokaPPVMH0dC3gFWX/Uv
s3MiY1L2YVqDwlmhjwplMwTNXjEwMMe2tj23XPtiPx8BFHpDGrAd8gLbw2+TfpZMplc4rkQH/vll
KLQ8Yrx3BHJo7Dn7j8s/GROEExe658SnNT6F3olzuE26EX+BR9vxhJ4bC3RxuGVYAN23j+itf/Xg
CxdnjbN4NVktxCKIgCUBoYMPg1D6iVyqFp4ZXp7JmH3eABJXzQUVjWSaf8+0S09c/7dTSzGr9Cgw
vJRoylRGOAdVknt5N9pelERlnuHjzYY83fg9V04s3TgSsP7goJtCxR5w1Ao1bm40YVSWHqN4tEcs
M40KQLwd3NMHpSdaueT7j2NEtWXMewEtxbdJS2qNGXEo1RPRisZfUobGrTkC2eNJWpOGrm1yA097
7wyGFGQkmsg4xiT0XCe4NuPI53tqQrmDSStkwsBomb13ulk4VedvgzmqsWtLVZWa2j/jr4A7XB9W
qfxBEw6QEEsQ1o9LH8m6a22czHmTIFL1htd8/FHnD6p/LO0cI859eVAB3SrO3/V75q6cxk7d6gzf
WBbB5DIR5M2lDzg9AJAR346V87UelBqpW1CwFG1In2ELb4KlMLzMkwu4FrMuWXOpFCjFHiK2MxcM
orBVb9Y4K1KIwBrCqMwcDSBToxB1TLSAs7a/ATfk9DnFJlZjSS4zeT+Wd7oLQMIEkTAJ7C+ah3+d
dpfU9N3H6SxD4RJKRtd4pcRhjO7TK6UL04/B0i8mU2d8sVElCGqh1KrXlvV5X2i95M+Q4Mvsldhb
azXHO40k0iR293fmEY3x0d6xU2zlP78tuAtzfSOeYGmncSALCp15IO+4lDav9KxQNE08w5XjScsZ
RzIulth/lZnaFhCE8+dDt0ZKxrSMZ3UHTMZE85nECM1qp4XqC2lH5cjBvWJ2rtTXhYYeEmCFcbpW
qwW24SXoH4FDKqSnQPpu0sOXgbN/od74Mj5Is+qyx/GZMtzwYpA25uXVUomEsKyTzJa6wW6f9Oqu
himYncKFpQDvHVwqCB4CViivNVWliTsZB74Q79u2tpLO2Gxl9gGERYl8PktKwYXxTwivzsMaQsFv
cESPOJOtom/sAO9ntScW/q42ZDFLwspZeY45Xxutj2FPSDC6Oum6/ehBMblUdXkEFDVRX+pGs/7o
DFEYR/bsFAWUwr9udhgt0FtoJfHwtyxqhkmTKSCTzk86XIVkwJmwQM1SfYbWxud7w4XBFYZqWx8Y
fCJDBK/nMhGXTVZffdRxdKq6pu/+Qyf9//3am8t+3QpEp2r5disM7gbV3jM/CYGTe/qFmIT5Nssv
qv6xCBuXMIyRtPomO4xZ6z8dSkBP4l77/FxSmBhmBX71B7p00f0XYnJb19tQMjM98vpleG8d/oFK
y+3l8gXmlKh5f0eEgExDhOTuC9PWaZ3NwQ0yzs7zbnOLgIY6leTtqx5sHmNXnIAJ5m3vk2Ylcppn
wZXI61+utlGr7+3jM63z/92awTwDJcUkx3C/DxNIUhKBnnFTB/C6COrn4jGa9jWb/KLtPPyGCnNp
Vhyf5VQUsz10IixpSfKC0iEWuK8FmEBpCI18tHBb0VHQ0/VGcIvi8X4JGzwNOYpYEzTnsNOqipNm
TApto6EwgRIGUxo1VDd/AoOaTO/zewfQYE8fKmeYGoc8lci6RZZpvbqwGKRBs8jpBBAhN8UrBEui
hrkyvnolqV50VQSOmu37qlBHS4nGFF32BPubfthCctojBALamsJg+mUouJ9teH0uq0M3M700OG2C
zWjN8+h1rphN8zKa1hhHWVXl6EDufZAD7HOsGvvd1qeCz/YuDgbmDb6Xha68g86kBLaxeSeqbgGY
rHVA08PzZpfFDHIlVTfaiYR1XtMKD7whgzp1XbEOJsDtSjryJLnKP2A2qzAoPnluzNoWOOqy9cvM
vL3sp0ThYXzD842bIUZyCwF3H5m62OiKZueee7ulmI++6KezkEKpSQjHMZF0WQGJ0W04aQlRAXHq
+pHkghg7mgXnJ+nPe3KVPmWvzSxsitEsTjKeS0G4OQDe6vQeDZ9Oady4xHXLqsEgqHAr3CiBPc+g
KmU3MEq3Yzd1XsZAzs/jh9gLwgu3LiXJdTAfjrnPvD7BL8VP7JQAB/xLPwkIKwgBR3thWhHbcNI2
XPlohdgM/p2h+7Hp3Q9wNQ27CDAF+ZH9HUIECj/6IIvXfrlzd8Tn67Zh8q3i1G84ragTb8WTlUCN
xH87kb/3mTrAN9c4FDJSlekFsVDoZRP01Rs1m+TyWunEYm1Rzd1NbWquw6pwLt95uHDYBtOcvLTm
NFgCF9wjYBXX5eRjJ+sccVcomHIIdM5SY0rtFrPgAEgFDMX1J9aX/6TmfrfXMbPVD4AYSYcWKPw+
fY1NTiSdr10JQbTt6Wll4M+RNFiS+sk1NJXPg/vpSMbNQktClWDXoWikU5+Kv9fUf2sdTBwDPKlf
AKYH0+lVo8AiNRUnY/eEuppMJ/3pMSAioC7lQV2a4JtOXSy2LQUC8hUf0ddmZ5hR2UyqKOW8AfWT
zmJ+uQD770+K1WXYLL8v+Tov5SHwK72bd1+o6pan7cRFPxNzbzfY+sJWpp5owKSR/mMA6ZdMmDFS
2e20Q4jfTlfM9XyAWt5/BpI0O5ScAG0O060znaggB0KxaDTy373JKaBE5gIRWXqoeGcYoTAvqhKg
d0/2iYqhQfqzhul6ke+x7jxCxr0IIuQptvLs1ERE2IK/LGPO1FrJAif6M0weVbCpKdBKuDQfjtvG
dHtA68zR0dLnURNKtAlui9PRB6WaeC5voxcOuJyiCcWS1OMdabIt5fY7xe6GZOnpUTcpTemh187d
zpWxXyHI/geJfP6f2lJR/86gVCea+km2AZoLjZyU38lA3WI8HPtxGXjsxYT1jd5dv66/7Y8zj+er
aJVSXUZpmXHNNZ/5z1coXUx+xW00jOjDsmPEBdrWK0RuvJYn5Ggw73M4Gl20zIHpL0OKuU5IzC8W
/6l8dN3WmxW2M8+Rgr9snZwxmbYy1BHiZ9uPCoAGdzyvrhZz6uxAjcLk/KsXwYualM6FtJ5KnEso
G4VHsZHRfQFRio4y/Yf0ccFupYIWLq9gqQ3b+MKrRmK6bwtV4Qp4wZlTEvoH2Ohdh918OHSrCktX
gRZHDWBdlTo8kGJitmcZ1nbE8Jsr/PfuJ3Cq9cuZdoAP0B+/QLnLuyh/1cLmIzzwd/RAEWOiELcu
qFdtzJNAy9jDymPQ6J8k+L9LV8vQWCBhQzr22q0zcLYK6DB9oK+IOdqkdr1ZTUyiK4ijqlM1RX73
LW7XhSYWMuB6RD0zq4HIaz8IA3SS7sastdRn6hPqKaMy3Y5+l7sZ0sFVShMKtmo89UyGshp7HP3o
I+oQAiC9uG8J+mOTGYpmdD+l0tRkRDvu59dpuJZMi9NMMBjTm3mO68Hj/bihVhGTOyGs40p3jfRi
EFADTJS1gmN9XrFKL4dSgODrRJo1ziB5kHbFUwAdbykszqG6oCu3OOtZB/u13Lde2upWOHBP5hu5
z0DQ9gbHPgtKNWZytYtBC1qako2/CuYYE6jGv2voxgSZH7x0zqK6bHmN1lBxuUhYk2EHuSMtvQVX
Cx5WFnHN5f6dzrgVwPZg4PCaJhRtN0ZzdY96cALe6IxXlWnXUlUK4M3uUO3sGUE/DBjK5zuDWVye
XCnTPbGL33DmwSyK7/XM5eYdfbmF3gETTPzNzV014UuzWOdSfiD5jU2P6klaz3tBQ/vuavEBH34h
QTTJmBOBk7d7fg/sPBCCVH+dixYJ4UiF0MeSp+ZCAHUTgBeYAcFtVkKHLDjosysZ7qk0br4+6HA/
yaRc01TsOUW7mF1aNdnAEsJOGI6V7JKg8KGhqL0l1iCmYkz3Q6a/Onhpdm57FQug+fRQfc9262hG
qM07sDRrJCSDiWaYm6nhTPOOWzcpIq2oIUBeDwhgJ0XjgCm4zfVrn/zH3MR6/t8bKeoX+9MRdDpx
x1ExPboVIXlHy0akyEPfGnR/RgIhvtPR9c9W82NiMcxdNg+JC0TblsP7DJi3YImv7q+/K1KEhCAA
5tAvs9EYxoDGZIdn4P/HUVQJjMzz75cqkejTSzWZ/9cZWE8SQCFoyzknLSkFGYV2gkmkXFyAP17K
tNFKSqbu5hGEXGWkAF2ECgQWzegjJXgX83m54mErfU2mjLy3Pi+7gIi6VfH2NtidM/1EnlDpFZn6
JeA2ufXvifJ/japZZpntqhdyRBaLzWbDbVfBeggstq/y88FvlnZmkdslcB7VyCrejY4/EvsqLkC2
bvFAPUfYZEqVUPHm8HJ0OG4Jd+SZ/sy9SGBUoiUUBoXA+uXFlXnc1iiOJ+quzk1oxqgWOowdpDXH
f5sZqUBoqWrsfAUz+vWRkDOR8MoOvu9JKpE2vRduu+7nvpLncblxosDK7LZnqprpcjKB/ZCPh7xH
ucNxfOh6w+PsHe4vE83azq0SjxU6nvp4uCsneX088az9WmwxGwZsA+5Nzqs0CiESivQ/fdbEJS4d
KeFgCNHYL+2GgorBwy8cjnAPAY09wMUrvMFzO3wV1qQjFbT0jBbHSax9MBP7SnSkwHQvRtg6/zCa
7b6H/o9f5O/qM31XGjWcR863im3Kb9JQ/IC1TQI2RtaSWwFPUWEggGgiKVkiW09WaKBhPXJssSK7
AjZ2O180ZRAQtiND4d8acsQoy8wkSWL3eF/tMrpTnElD4Tc4H7ZNAhEX5ZuhzdTbH/aYBGbGopLS
Sy3RisHdDBi7pZi6/Dv6EDBHRBiJ2IVgGW8uVqaK9FhwgZuoLnKVYaSLQ66cSTXd91owUtTNADQH
VYS6I7j5PiO95gTkxpQYcwMPMVcdIUE229k89rocjxJj7UQsrR2RBJvB9gGd/kUj43Z6mM6bYOUR
YG2P9Te9hjOivxceWvwn0nFhR0pseLObD2Y8cSWQXpTCAdySDlM+ztUzhgNqvAiwH4f9xnwhUKvT
70W007rTSqzI4a9DtJwx+saLBBk1MLtKhDVWph1eLbCRUnjhTSQ45ocTK1Wv9wEpwPeMzmXR4jlW
L1QbyvkysLeCjEoaWdRFX1Xm6sg9txm+ub8b8Fn3ShpBSteXhGZm356xn43yaS/kTaFYm3DsWcWq
giabZVpMOGPKrDAVO1C7XzVDhVusoUfpCWnvjqyIxOnwi/F83PSLCt2G9UYfI6tfX+Tm8bkEXROS
4/92okunfIGOg4kHFrRiWfXue7dUaUTdvvPyjVymyN5+KsMv+PvVF/VaKC1AKNU6U3wnMWLzaS62
mBxFR81S/lEwgtbCsyp+jt+Tlm+IIcF3jcoBsiEsymo9PF+FCeo5PbZ19v5SSBooBx14Pnedswq2
TdGLQhoks7jcIaoDmONlyB6s+ZaBYATrG3jbvWut4WJKLOc2PNbbdX7EtwGRcTAK8rE9nClUl9oZ
T2jCIzaA8XqFBL5h/T6k492rGIwQ0vABH1lOEz4su/UvcS6Nxnz3mIAoqfzvUrnszq6ONlnamFAt
SU16EL2zkFyLJnKnFAmKasrNK+3bz0eg2vwCuenS9TszQunlGHlYOU10hP4VFax+GsjCB3sOLe8n
wisBMzT2hqWBQZkepn3H/oi+5+cA0fxUV3KpE/l7jaZhGF2OGtAl3mCw/PVeFJ6AxqFMekBX11Vs
VmgFsfR/CF7udprb34xxIGqSgSizp5dYKln0Sy6rW9htBCM++bYAiDXlgm6jOcFSFhTwXLg2NpOb
5j8psZ/3zpOcYdVZ4NuWRkFBNwadjXsqip3QjR7+hqcEiFnMFXbRA7ttLgo/1R1PxrP6k+FJxD0I
7rtCanM5E895/OSnuObm85U0850jmGIv2FmlIXiC400clC7DAMuVPbGmxdvz3clMqmKpVH+jtspg
QwWR+gUFwAvGlV+Miv64W5xJTFsW6M7xKnc1zxBRqT4xVQ23UV6U3Bhec4Jd0/N8uSdhgSNdaxjr
/atlYuwcAu7JfpNn9UEsmNRjoPU39ak954HdBpI7KyuHWXlRXUMuScdV0nmdaeiRqRwgJduqj1sP
CH5gwzTp01tkaIcotfuphrqxeRcuUtsxNFmtCQ7Bf5IEDnyAY6qdSVZZpWsFAY+W6RDIz2obxCkr
IbEwGfbBXbd80bJ2kQydpCAA7M2qjcCtQlXnSwXQUqPgauHJ4IeTcM1u1i8ip6tNpDLxeYkfmcU0
lnQWRBhgljssSWnamm+49e+xu1xaST+KEzvSFkwX6JIe1x+pnqLVbrF+ce7wtFLvdQbNtZ1+ET3e
v8qiXdvqK7+KuYIopUnq2QJoJPUK1dHdvMaceNpgNN8QFhnx+B0zo60wx30RBIxHSMTgwKgSj56x
Y27btEWOjAC+j/0TcPAUiawvNilcNxtNjSorBfmrRjBuT4FuzYIvyEEI0MgDqWepEgOwmVRmqPUu
emlpjgZdIMfHuIMTaEtoDc3N9Xeni1m3/GGoH0mhkmbCOdp9KU7WX4KsnwVzVmgrJ7S64YdS9Yg7
Sy2NqrekVz8NeGKUVeeCSEgQcsruGSi35wOat3rlUT2MYAg4H8NkWJsl9JC44aG76N7Nv4isX3oc
x57xSoSFN6oXms8f39SsvNG8ruX6Rbt9A+ou5Unqf3AwTgqQzlpVgWXOkcjrhJsKDmS6tQzv1PP2
tQvF4GiFV+iZZ6N3Hdcsm8EjPRkCX5f/VBcnnBzi6jZBnxTEbQEdEmCJ67b54QnB0VCmEmyE85e4
52fX4yRkaINCZXKIGbtP5/5z5i0y0TxZJOZuQD/92GdOuhMXFuY1qoi7LAwopdC9E6NYGG8FZQQX
T86INa2iY3zCDK2Vtc5KYwp0YxeoBgJZW2tuogwXwiGYZ2O5Uuft8+0UqQ0FB03dbK5EGfo+gT3V
V5Lkp3RRAxY7AUdY2FIlzYfabBQMsmw5ALEYil1oMpi6bZDgP2Zr9JCNQckTCPinVppJ8fvbN7WK
lZyAbHiconyeLwqT7UUPX4S3tFp51DuuXCJqj/CqwyZ6qJuZhNbkVcutu85MeUqzHPSCmW4IuXjV
m7vcBvMmz5AmzWrdtfcKjNARJmvD/HewJ1dBYBeOhlcZhHgkaFbHf2YE+7Su+mwOo+/gBwbW7zS/
aoQ3KBYn2cYNDncKjhy4sRzE9gQHXyxfITvaOZmDlUHGYFAqAxZT5jxLkmHkhm1YvKrEES3tpM8i
PqXG0YJJI5F90Z4KjcJQQozMXtfZE6h9G8Pbz3v/lO+JUqm++Isj2/ONqcNJG9pNub48o0dilyRb
Sq/joT43GgVkPgcFsPsJVsL4ufIlO+pGiH5USjWhPcAmtLy+kmqQgqIe0brtlvHWXd4avQ7GXyp6
V7S+n2tv7QLRiep2cm9ISJwMeDTI5CvG/IOB72fhRQy5+MCeYf+UR9DgGnfTz02IS3aJE12qmfBd
FxbONVLrL+PJ5sU+ho2vOHYM9jWuTg0vJ+wLkg9DNRTrzeOv5PFWqO+o9TyEoGGQe2obEiYojOcU
kHM0PjprLsvyV64n6omjBS2AOXqTmUC3T/6h+Q+ZkS58sF340EjGWOOGMu+Rp4sJBNDaD2VUY0VQ
Ar18iIUWQ+in1NAJDsq1O8J4oWDEluVCjYNnDp57wBRCRSMuoRNzHid/GCjZ942LjpWhcyEmZQej
AaFFnIs5G4hefiSc0JOsv2XsACGgh1GhkKvGZpMGItodqKmrKk1yYy7dgx8nQ8pAJZgVqorzYlXy
PjlLRxCaWD8LLAxf4kKueoOMe7MDsyA6RwgWyRfSytG7amM0ihfi5yI3NrgP1i9I5JsPYOdq26ps
YW5qVD7wYy9vw+6fuFbXRl/ZiGjIiCpwWQTA5Xj39prvMkieKEK9auiNsoqDdyz7yVRjTOmEH7Gt
uZj1qVhfkNR6iRkhGSi0oE+3RWcka01PmT83bFVJkn7AITQQ3jlZWNQcrJ2OdUhYoMPfWB0RavaZ
9M7e4lnA2rzhBYpJiQ+jIFdGz0bUG+secDAlq4nPKsXSPoKVe4ZaFHw2WjL9qYhXVO2wl74cWYu3
HfSu2x3wOAfB4f7LoXeFE+Bj8NEyuBOGoKRdvEsxX6fzM2AHg55T7c7okCoi5QvB3bue083+Dedr
oX0HR3Qef9M5V+YTuBiXR4G1WsceTJS0a3ZJUavA7z4kWi2Fpl+5L28MWhW/Qu1a51VUYgPWFQEw
A75TN/lnsBHeULXw1pAUHQVy7XLAh7lfltAqzGEuuA8QDdmlP9Yqi/3vGEvDMCGJak3DRIEVdZqe
feuwrO0iwE6cVVcsZa2M/YVOQR5knSDh7QLEf2zwBgoMmw9cXTF/ZMsQc+E+fgB2QYumQcovoQSW
kBA/gNfGI7haAsxrgq3oJ00V6HwNVxvDHgMf0cFLmsf9CdvvNb0WOLMSTh01AF2KhVwb5/r0ZH28
5QGWaXa3YftZzQeo6Q4kINhunFTErjji5sMRDMv3udp8Qk1EiguE45zBIpLq3xMNYkkd+32tLle5
Tw/ubkYLq6XYjxoTGiFpkQeGXx9rawVYlPsTFwh6291L50Y774C6yrFI9D1b+Z4njs4BvVtePCZ1
m8uIwSDc3udA+6H4I5KXKjVGy4Vfdb0S3tmw293sSl1U3SZZdTI/0ULbZQlEBrrp/pWnOHgCBIOb
Z2Nuvk0HUswdN2GRPRnXp5RSdYkjNcmVvsz1jFPVZF/dGiix+uHuuLb4XFF2+oYRmlYgdC2T5t2z
1mPp5lnaHLk3TKDxAQEgUpo0sDpWuNyAQ+QL6dBhaelc9GoDyvPqI5OQR8eE/tkmWtHicroGQVZ5
ipP1rGkdfLfthfumC2HRNdKEuWz0ec/PwCbuUDyF95E4A12CEU71cAmZ5XyXpnNcFkk4o5aWYTb1
gOtcpgNb0woHrmd3C6DoJ/UI9KzukF7H55rp6RQ+XWIUNGeFIy3zjxVJoDk4DWNT0eCBJEp2Q3gX
5U6Jjqt/hdY5F3XZyQorKj1bRfhiLa+ox1uTdgyTrETJaT3SujqvyQnFRtzPcvhmHg23JHkbNNlp
ROLIbC2oJXTQ8eNl4Z/FgNUlzy/m5VtAGP8+ZRO/2sy0qAarMriRMb0iJAiF3WDcLw0CvYsoDVWE
bcNn6lA0SSYbX8JjQqq/lm693tVrY/UYeWNMffoWPgufyDN2CuoG9eQ5QL11dvBJ5d2czjY/rZnO
RM4YelEeElaalsLLuXCc4573iUicmWBIjGFYgeNtgwrOEx4Wpzul5gUbu0t9LZfcsZuSIbc0t0H7
Twkq1ZyNKE6KeOxYSprSEcKeeyEo14iqDhU5ThyrcT+E/mvkBOSlBvm4UH19O8QKOk84p821rgNg
1xie1zG8A39Io1E59MhY80+Sa02JHEt8T6YRhbQYI0wW6fS/oWaAldasZyZivIHZhc5J7fWXEbgN
HX2u6iWNcHXHelJozPW6NZt719+XkJKPPr1Mb/1h0ac6XFdv1pnhct/38/gNmhTMroUEpmVKB4Oy
2jGyP+LVlJpYFoqBaufeioj0wUjjdEJLXYWqdxzcRNL4f4FC6PCxVpMKemNuO8FXFJ83CBTrXGP7
rvJ8tXBsRTIvhMKj5wUpMqQwjeSXpRDnGMOfR/CCp5vHt0GHmbLbi/llICMrSWBO0dpBbi3x1abj
9NrMVCg0JDU0OvAfE3N61Bf5iFcYiG5IVpNHBR1k7xYprqk67e9K4gTXxGqJh8YYXWP7pdvCDFAE
bejcvQd4jJ2nf4H+PxKUlS33l2K6JPP4weSZ33ruMNGsKBD+1tbPtXW6YdPs3NOcIC/kRewuXQ/N
wNd3JguPXpWATIPvSSlUqEW6HUNCHjOaFWR3Eu+4mOVLL4Xvm0djMiyOoMCv2uVkW1ygsuGfN/VP
FIxa4WMa27DGVO81o3QewuXqjrADfBMdWWw1UAUoWlfViwwJ+7Ug8sDYU4n2Cr9Q2BmCY/ogvIg3
/w3K51dNcjz1ox0pNmNSumYwfYyM55OQ+kw+xJE3TLUPcP/dxYIa9hBrEKwRkBdbwf6ici95ttcX
5ycZOSs2HvRBpbk051ewZLRqGGOGxUfRdUECK4R/QCCU03FGWF6NDVQ9hN4Xq55z4b88zzevRjl3
d+CFuW8u/CIuHVZpgNBCo3DhX9vdvfbvATPVQrVqKqqu12mO1hXt3G7Ar2e9nDpfskVfG3ySIDNV
ZVdd9duS8gIoPrrqB47h1/sBngB6DdoGKPRCZbHM0l3MmivLn36BAG9hwhJoH382keVmJEFJYo1J
DCfMINkiHZ9j6DsFOGrHlSe/HDQ4rbXs5MSqYcrEun2jXbSrPZuRT7vUMhebA2OyhasrpTm3enMI
1K39wSmOaO30UIBDije2fvPCN1v2ryuSZySVKUnyIdZiFBo64vRO2TFSsg2Fb59slm9lcRq8pX4K
cCd4brCZej6YkJ65WME8g5QAQW4L5VOkyCSWxX6do23RGrwXhT39MnZbraUhSk3TBoW2qN+zy0Ov
+bsy/b8D1BGcjGkdeB3Ewp3wbLN1n0s/VZWUCjmFgdWoFNCOSmTxNns1X7z+njTDfWJZbESsj+qA
okdANRxwLaKjvZkOItewNXt4vRxcrztFmwQGXI3vQuOtxDE2NAoOn53j/cjvvVjWrDvgisaZ55Q7
Zxi4UEtrVOuiqnWoE0tNTwgTppZQdLvtLnaBCEy+Co/QKRd57W2VCfgCFJ+WwIKrRJV6i96bpQ6X
N+Rb/X3x8HARK2ruPEuYxDp6A1Kx9MAIgqZ9EqwcxkOBxXFIcvpxmB31iOdT5BsSeJaXY31pMIg2
7q9DBPjDBiy2McbuyAm8EsHcT6XqzIfCjMjfs6VaiqnwzsWpzMKhbQZNH5M1sFkZA+U0faaxGspm
8pzI+4ZKgU5STXa4/vNARuJM0ioFVF7LAP76dGSxXHYRkyby/qye/AmlkU40Fc89zA6apF1ZK9X3
6Q7j4gk//lOZmB2FE/2YP0mMUld1jAJ7ZreerJr1APQKM+b7c1rGDPnRYENDvv/sLINXcdk2FwCn
AfRDdcK53EU2Y4/x8P4XUsyXO3tWlsiuFTXKWz0bsnjMHC/+vXrquWLc5M4O+aQ1Vq/VAGhsYW/l
mq+uSEWSDfVUwpc/myDd/5TAAtogXtFt90IXFzuSgvffVN5JmFSBYgfgkAho0Wev4ODbiqn0sWCt
nulnhJkgNn3sPFrNGwOSHSyqz+gYK3vFR3UoWRE8olcg2v8T8A7M38oXh3oI60xF7NQ7qY9akAoj
PcxQSh4lzSTaXN/cRO10gqz9xNQ3UIGu0+XY1Ji7W/+keORqQftIdZHXKrsC/td3d2ly/WXzngC5
XzlJSAbkMThSPlWNdA1/9DJqqZjeSJDu/SaAJZW/FA+HMYRziv1aqyGDTeAElGvrsNGcD1VKwA+m
Ypr8Qs/unVYtVS8qkcdsC/DgOteiG8dTJi5uCH/kDSW2xL+vo7JHF39C8opF9kxWndUFynqZ3vur
6enGxoJjIse8lAssGjhROrLEHaS/3emwulDTeSIcVrr9hVSUz/X+Roys4mFvHXrP+YWMdmebW78K
F9SRFgJ4VE0Om6DTfC93gB77BFA6FLf2zL+7ULW6V5iDzPi1dUN/WplMsiggru4MwsewVx9xNMdL
16uWtjdDGHMRxTrscCBGhzQwf2SE+XWqx69HWv0KwKoy8PZ2SzrwyJegiaLRMxPHVb9yjWfB+iqw
OFOI5vw4TOE4UtcrRCW8H1eDIpHr2btSCVT+9uFRkRLqvFbf0tfovsFY52ldknH3iZ3+V3h22G4i
NJFfNoC+3eIxOkBk7j56p8U/ezYUM7DAr8l+Ryih7vb+zoRUUWapmQUEgl4tZtPnCY8EvNG6xDZe
0qO8Y3BDFgJ/3W9IDzUe+v/lAMBvkJrgHaaYUF1ePQ6O5mljiYdJ2UTVYQIXNG1qi4msbrJ6wLYV
2VW/JwZe4E+WNB9V8UNQaU5kKsyvE42k9nZbqHlU5FU+XuXSHYkd+kQLEmGxwyLCVLoqUngMzJvj
guQcqJOTL4ZpHqUWD26dUhR3Jbkn2sk9FW8ON0XpCj3lE3l+COgL1PeS8+q6lXPfFrLyZfzdeZ/S
ppLAiIQihe2eFLiMjpMtSq4+91sQECSK1FSKLDkMQSB/rE7FrVcAtrVnV3VKsjaOQ2KIHnyI8Tko
GdbGQde+chJIFbyEP3XC4+wp9+gNXVgIVTn97v4ygRiMnizRkqOywF3IE3kSBCEAKpiUYQ/ycP9Y
hElQThr0INANCzzodV7DPSj3xT4V5ydpOS3SD33qSiAZDzOcB6Cz58UkglAIZlRvzU2ahS+2MuI2
YniStmkAukMhMbnVVEx24linV3KuvfyD5SAtgkxrD797r6VkMpv9+nSzaWc6vZNx9FakqnA1wAzA
K4zCV03aQA9l5s/qIBA2gZIeJtyG2FbFEBj6v04pUSijhr2NylCNxk9q1qRsuH8Kz2vsXCDiVeiT
MabUGfkX2x/HWRvTRV5IOrZ7Sc4FizP5M/KcAgJPfewhcALdFGt+wfARaaGuiHzGHKtnkDKeK2ld
B1mNJPsgPa+K1EgQHfOAvv8ECifPQLzlFuudak3JFnLqDoN4i7X1uCnJom17oF8fDOd1IIMl6OWp
z/M+tdOUAcn2VCvU+rHmLlno9B3VP119FKQ+GvFz0Iwn3umuWFcg2alW6chxZ0Arv3S7OpZa+4tS
SmoCjj08ok0sR/GIj80GVoedqrro/MffPDoM6/z/figFIXyBiX4lr1hiiKACUDfVPAxmcTLp/e16
ZFnM44ZJG9sEIpcLV2qfb8UuZKnJtCG01vLp2YQCUxP3yd0hIdtAAQHE+NB2xtNmwQrrKKRhn5Kc
AIqFCDAU5Sr0A3gLLrNXyn+0+ByTwIwIFO3m8fgFm5pAIHTFLasrsgiqhO1bpFFMtUYuSQltU2q3
5hqnkYfWdonU2lOyb4MbEXv1O8pC5aUwdq9Mlg8J9Caoew4iMGk1xRqBYzHYAV5CaB7sYFVJx+mw
0NdDI5jTC/p9spnCiwCAorIagJ3Hhj6NNJtDKh6lUdEHC1/pDuw4fwY7NDxiCfU2OhXnTnvfs4Q+
VPkNpobxMLbP5/jqYKs2Ibr1LAEloKR/lBM9/Gux4W1Teio7xQfRka+fotMaNzXoaYXswgboL4Uo
BfN9SoxE0JAtZWOo/xH0+zuceS22sd5hPrV63jQBecM2wkn/tsdTglH5NdiwE5/uR+RAeMVHMSy1
rqif5ZJrnzeLz+E6aYwrZ2NEraMMrjHsnoOxk8VIySJekPaxe/DzIvincUbGWgVF+k8Xz9ex7oVf
LD5BoAkx0PKkVX/tW7ZHd2K022T+DNuaBKn8pQjBd2WTpkr1oLbdolonbVk+jk/Cm+zUloqz77VX
uPx2t1tdkt4Zr+Sqk/ZAzYQiiXTnhvSVCVF0a6CXvbIi/Am9wkEOjidYUC+scR+HjGIoHYJ6K3ZZ
c3aC/Ons7u2XVUSXONvt6VjHnkShk2/w4m/f3vM2bIrvO6vnaejlH894b3z2Nx2tDohdzSpkQI0h
dr4/sadt4C5FZz03gklgXiA2k6c01XkORqU/1OLoExvxw0/D3jeCqc22i8zP7MGxzJm0aIQSsNLT
/6acmHgt/YQXtcxC0igahfG13kNmpsjda8AHV3/0Z4r2mBW54eZ+fjJeuqOTJdPMFfwj+fzsfU5b
OEvpHiGXtKwP+Dk2KtP67IUQ3LrfkteQ4AhJkZLxikZR4rg/K+iAj4I/iILVES/ExOXEmh/Eyrya
RQ6UtgG7Cc+0c1RMsoI9EmcoEXjGIL0sXofzkHta7i4O6Q1RQZbRjIzBIZZYUk+5SHEEn7liZ3Kk
Ej43neTZFzEPbIeWsUuJgXxLsM7tAU92mOWPvWfuO5g3F59WJQ1wfi5miJGvjthPm8jmhpr4srPQ
f81fhU5bXumhwDWLWJDpPSSuTbeqhkpJnhRzql2L67SLbHdvQSKFHdHLrYXIPPqvXq/WkroUh5M3
EPMPr42WaeOxJx47Je+tB7yJGvg31/QEMYDIAFmuI0S32vEXKDc5KiB0VqIRTEQRWVcIy0tGDAXx
3ZlfU+R641mD2C1NlYKOLUEL16uhOrOA1CP2bhQRjIP0Suz4w/mcZGTkqJddg+f7ngxAQPiRthfv
a2k4m0nHToQjEzYD+pZe2c6G0oKoImMzcLJmPo1Z9zS1M/xc1gxHs1u5aSGBUdMnLQ+2/wMwrh5I
SgeLnpJBWujj5gz78ju/j/HSoOwqb/K5qNPf7zU4leQGfAGXmgix0+LoCy3GQ5lXrmcCgE0EtJ8s
OgUfrWPzyZb+AHzF02ZIiQhn9/wa1UEzRU7Ke32BtH5OC5Y7diDcw9XPoneQ1SxeK3FqQrhnKbWS
UKqi2+Csz/O65KDcWM0j0O+Mdl3DfX2lPZSv4tyrgQX9tvclHtdSQdh4SkPI9Fjh1HGoSbZf5IrX
nGaeSdwKWcOuocpkB0pDvJFS1CfMvDQ3+OVdNNr865jW+ZFckGl3LIo5LaCC7YLYdTdAPf/EwFTD
PRtqFsRtkFbTGlLVC9PYqr8yz9yOcVMZ106aY2D5IBIOy6AFrrMooawCzkCvfRaxAWZC0CDBP06I
Psm+eqkOjlWQW0E1t/2/87h8mrb7C5nHERUBbAH6ZNAAfAapTsmNhgpdv7ZBSyyi4dgj3e9cAXQT
RS9pKeQTBsY1kDMcCPi0aklJ4j8K3BPQR76BFwDu9AWq8oLmJ43U3aVrGo0+udguQ5MmGOb6tOBm
ft30/vonkQiwAYVXFvLVbjo1yOvy1dP4v+4raDEwnugCABHIwOz8O7pOQuhesaHRm1v1PGnTkill
N0RDbJD1Mw3urzn6Xm2FPVRSHH++jMx/YRfpw0skAoMUA8CPtotpmGHlSyFma1XPDdkiIrolfZy1
x4HW/osRxfMTcyKx4lWTpSTG4VuMDjHmLUO1IMVq4kCZ2nf5rWaWS63+Ju6UCLcB8g5IqU4qpORs
JvaamELjCrT+MUObdr03BmCOea0ukiwEUaLFlRbalvnGSG6t3hd5DsOZkaoN+IX6pyRTLk7oBlCu
W7va+m6v26PNO+SL8FSuncMHwZva8ed9G0504WXki0e8QYoAaQ8Mo855o0pO4ps56j5WYAvie3OI
WCkmnJQ9SHIKLQrPvM1PncWXwKC9ptKanWOKojwL5sFmb3HLXTztiNPl9lVv6YFMIqAxn9PyOrjC
hrTn6O+lvdMBTZi55SXVrEInrAZ+KXUhcit42/lnI7c1rZPmtuJm24ri5KZxQ5/L7D/NXrkw2tVZ
sUkBOWQr5JSnUqVKVNl+RBc7bf2UJfPjxsyzMMJgWVGR4fpM1IhIQrhHm16lQ2px8EjkMnCL1Keh
9u1A4ByAnSDgLVjI0gkl1Ch2nxx78vcNkWMxY4JnKRcq5aTDXB75RqP0Blu2RLdpJS5ZlfmjzKQ+
EStCYnGdwPWbg7i3kra5gx3Q5noc6ot5Fus1DQYCeqUYdR44kWLihMwJgIAZ6KAbUaOc9C0sge7l
8X9Y9pvFoN074/QECEKS+iY6fVraXuTZOPOAXFRHZYqWd5B6nOwyzf2dmdSAb5MmpfWc+QXLKQCQ
/rjHyXShhSJX+RUeNuqk2QGibpcMD45SYwnd1cT09Ma3lYamf5i50XjbWIJgO8cM950MhyNJzJam
i9BEFcfgXrbn98N1T8wFhOjsXVbxIdp7h2RhDPo1cTTOIJkjAeacXMstQu4HXPhv951d4zp8fWSW
Rm/pb/v95iivYPiyyawxse8I0bmcyu8j/EEFi15GGDl4M8oTnpwwhmQBsZA/KY6goCTXuSrFuuqP
uC2/ko34uDx6eftk5jTN//ozRMqua9R/dUdjkko0wUzU/rEK58yx1BkLwemegO039T95dSBQDvFj
mytNsLyE2ZzQd/w6/JMmUDnvduUMqFGQ/H4aUp7yFIQ0h6XbkTciP+YC3k4x5x3mYsOSVguXWOd7
LT4RBvG+vuPyz3plxApqY7FDFWvyyDWDlgfjkAZJtIMG4XE9Q5cIx/KMuXLC2N5R0VGV//BI/kzw
hYwnm2MXW2RJJSy3YO8E+YLLiHHTv4NDXZ3Tvh0Hfgu5LFDbGoaMNkVBQNm34g1cnl8ZbE81ClSM
ey66OwRm1GTr9/26G9T4OiqzJ5ycdAVRGUa4aLTde4T9xUR545Xrvi5OYslPPRkUzh+7Uffd/xU6
16vtCW9vQUe50R6rE4gYQP1FylnUX4VmJ+VOnnLei1IoI16l/KYbN71PVIbf+ZLcQTJ9WU/J5ij1
tNKLtFmDJHrxag82edK0O5AWl9vXQoC3PTuk8FnQhmPw9Ha2fVgshT9X2bUozCN+EWfrdJYBJUzn
tW7XyRREqx9X2I3FJMv+RXhpNud1H3EKxO5360atBiDCjQiMxtdZbYmB+PX0KfrR+UjgZ5aOsb83
+NZSkImD4i/hoVxnyGzJjUb590iTlxyMRY6QtUs9bQzuTr916+j7erzL7Xvq9h8XV0kU+ml3s/2M
a3ihWvlqRXtsgRWdQ3JwMn/yw9iuJGOb9SQjCbdGDTyZXKc/HUsYtQojsUMWlUjPWyG62dMJdX8R
MWwauH4spOLeH62H2SMxSsvhqYBr08SCRFVkWCALja5QB8ry4bKYHHE/hD2QL+NMl8qiMG3bs7CP
uuS94QuXg1taml5rEHWCtDJ4iylEuCEwQp8BhMJce3XF1bz3vtalbVDG40HLvhYnyNhYeWWXI+8k
U6usdBL3w8twt8oEAFjsEo5/pPoE+dURA1FdI7PDWtCaiOPw2DyKjrH6/0foW2xNHFDKW/uEyshd
asy5MbhXSVA/R0NLvLICwLHhrfPiK9HpovBNcyOV3rN1UOa0q4z6x4xLf9AtFQ8DtRU/KhgLiZRK
nP7h3pE3FwaWzUvfdfT9XivZmTiMAq5oPqMv9lncbw/lEoe2RDdyNuZTQILtn6fcd3PC3VmOmtyp
7IB06ys+tbg0LBwCYzCZ1w1XI0X5uzpJmTv2pIKnzxopvQ28pRC26bKu9cxXR6U22XiBwwDo8B4E
i35/nh1NYsbWYVOdrFvTA1d7fJuUgWYN0pZJ8sxN9XoFKemAWpyzI1YEkjacofOhUjlVR9XHQXES
N7JMiR5F10YqgOzPoL+N/4pcqAIQSKwULuMAbN9zREtM6gh4Eqh+RXpY7QN6/kl2YGwXUFDtKk+j
7ixPqtCTythj/FCxcb+z3yzPOoJY3JBesY1dydezbNLX1ZVivzpHHWb4eB/yVpRHzbdz23zw7963
HFazYoROqpzXPTP8JuUvhdLaEh+GqSE5jub0d0fUvxhFYG0+Mj+o9uSrux6gNs53zfY1QCjlzM40
uYr2NgYVu/cgXUCID2JBCFF/oJyC0ABbjU1cSUD9oGmg9v/mv4nICUjuLc7+3DsP4zxG37c1BOMU
EgUwoi3GeMamafE3kiJFvHBUuL5k43roEhlEjC68oYqgo/DqbaCqcP49edRhve2CmH6Qzap6aJRi
9M6zBSRoV0/imQ95KUIh0X4F1IQVG1YbilfE/DxWXcYn1qQ82GNgsi1Rrp1AhuoWiuRA/b8GlUOj
zEmlMwtFJW13D3jvCBHt+MbVQjfQ1DBNekstI7cYHvv/2ULoMINt/1cy1aBXjOyV8A7hFI1ENuM6
DMOo6D6eY8PEFZy8kAYAULhukuFGNHZxKRyx1+QBa1MF527OLyJEOXEQX7OnMNYSYg/Ml+HcDOae
5rVg87FxVkuI7zwD71AMJrGQwrZ0vcHzNW8jvdqARqW2f5wc3kHJJ46XS7uhQxNUeE1tnSZzPhwi
baQpSBRthJtt5pCwqHpR9vgw5blGJ3IYLbKY0cN4XXmV7KKTdtmB+wMQ5+PrDMKRreB+N7+Z7ilG
GGJi5gzhuFuHMguXeNLAMmHguFO58D2uuNufT8se6TnlhBmMZjWIPJLQI3yel6xQrtfdf2uYrUlc
H2ZZZNVunF/QFnAD6T/eP6ZNQF10ZotQ7jdmJ46/H1Aoz+lMCjafDKovUJU2H0iLyGMgC/gHjWHp
yDDFLf/FlPMcg4PJRTmLD8UVMWKzBEG08VG/7poPb+xkFkC53k/UxwyT8vAJv7JFNzoX/na2kHyf
Ji39MvdwdYNcSGIDcYYZ7gkd9opyX1J7knCoX64/GR1e/tzGZid4Lq4RwzeOq+b4f8ZL3ByowemQ
/eS9usZXw4VNVOLXKUBvgm2gvvOjU23KdDdN2KYnDjyP8gxYK1/9JahWR9RU+e/7fZYGcWx9fGpD
PiYiPAdjMSS9fsJ7hjDna5kCCgMytCcWyP1cvRN00Ht6q5JSAotiC2vjyPFzgKfvtAwSr+RfI17+
HCtIfJZnlnMgSC0+stBn+ujhIFlBVHom+yFDKOh/1hF5Y8OQRG+6RrJ8/nVqQwRLIrhov0fOlaIh
Fieh3ML/9nSCyXu8HPFGPZLy6xZ9KH4rRm68vKuN0hwL+8EyLlyme/uD665fmQFPsUgmd+HqBNsn
23Vs9d4iINDIcZP0mIoNTiUGjaeaANEpUrkE/7Q2+mcbmuj8AIqDfMUyjDxwvdk1n4PwMQkeu4y0
MBR6XJJm+028cVVsgD9Uxlx2tIvceXBvENaz5tkCJS+OAbrcTcfEOlmGozUsCQ3SDMsDpysVRcER
OUu9wEYKan1KqyxW2Qg4lgG2Ss6pprjClJmEREGgOmSrUPmdz32KVpNJj1DQ3cPYnpqHBHFsfQQz
u9djTEhcd9yQKg8PTtFiHS4QN+mVWDhskP4ZfP32AwfoTODFpoUjj7ITCC3Wl8ZmsZlh1ztBZYkz
tF19OH74W6WErONKonM3/k0rse4p3Q59uQh9d1ESZJgjl+NBiabFpvKSQnkgu2+12La7iFE3lSwz
AmrxA/3bBeZGqATMllB5oJVBsIYkQaxEbz/gWbYvSNiAkxc9IZaSLSSWV1KgrjtaWrbE68E5qkV1
snm1nIQhkPmSfhIPSY+i84L9tdcVEaDDceAaP+FjSlJW3Lbkdxuwku5t25Ss9KsXDDXSimyxNalc
y5DeajUX20UIsrDdLFO4yGYWHphbA7gdoNdueHTf2Xjhq9onUB8mL3d7PSfmK9M3xg48AVByovca
3W7eFICdYsnRpn2DcmoYrRGjuW5Y8e5m/sDWotvMid6Lof9lkMhEqI1Am15FMfBD0NnpUXrFO8VJ
rrEtCbJd5E6eTJD1wSlePY37EB2LY7k98yPn3VdaqMa4Rq+KOIPep1QiF0s762hLC6ZWi8fyYTFj
h00v7IAd4F6xjdh90aylx3rn7h15XYnt3KKH3sAFgphGtkGRjO/0/+TaqK/udmJ6Tl8/je/T4Ngo
7qZGL9i7AwyTX3/Biyiig9+iDk9/rMsLRGv2kAMXy9ne8alGmP+jDkme4Bb6tofThcdfZM57dXtL
RGnexl0gHGvtwSHuTbWQ+JOux+v28CWu+F+pvQ8LAqTY0Q86MXyyMT1tTKxorKsZ+nD875Y9sQOk
0gWVV1xZ9753lmAExZYYdvTduGIYC1+uUqvIJUnrcOcqh5zORcMsYDg5TRTALFk/WpqZvp0s8u05
yJ6JeW0Tw/SVJ1Y04QjJYOtFEDHjTkok3HZKw5pTaE3Uudgt+Hcm/NT2zx+tQk5tw5d5d9DDvIvX
BXwA/+QV4yssbODL/71ThPxPw7fk+/2sW7jdGRN1NQ7mLnkWvkDMrcMy/Q16TFdVqVgtN/obeX2L
MtsSwnh8WXk3NC9cg9+Rt10jmpmiMRguUH9XaCIOtoVhHWwNUX9m8Wa0mtvoFJd28WzSc2BIj3hR
SrXs6wHnIcsgbIxzl7TjckA+0lYi9YafUVl9mf0SFhSxqXWQd81ZJVQjugRMmq1WCqicCBkyn1+O
U6hwzC3x22tNiXtPDr5VYA2QikpUMQG2yGpWs1iI0LgF8Fh3pP4Qnv4sBJvgZGt+4YxKxPPC1mMH
eyYZPjSYONlcb2upBk1F8reRpLrLbqDRys6np4c5AZdRy8cBKv3jEiFYRm46dqD/kIjF+Ks088ob
kpSDYVi2qz4WKlF85jhc+1ncbAkxpDoFxjd2Yx15tvRbb1qmqAdvFdZFsUr4ghrSX9ENCjZGT4DS
M8y1ksRQl2sECiL7Fx9o3237NggkACIJeSYbNzVYq3T14qbmaXAknEPCxXjST4dyb1aDw+yCJzTC
I1ZC/YfphOwpFdpE/Mu2klGhnNvE+Qb0IfUFZj0WmB7wA4xE86fXHiZcHt8j/fnf13tOWQDr5Pqt
/FfS/MruBQxZu7P6B5rLkyHDsHF39jTeaLa2SpkxCpIV/BISym3r50A5PqhkyOdrLp9wqx3hDFbp
EI3+ZdzphOTDLhM6raU4sasYKWzhM/pRXxFVuhagtRANfk2CjANpTgjhEdCcqha3Dt57qngs3ylG
aSHhcXSGRpazyh4uRFP8Sg2XaG1rjQGfOB+4/X/Vd/wINFgZRB8XQMbCtzEwKZ2xr4PsfkayjLCK
jhC3e1bIq3+DbJTScxFVB3x1dT4+hpEKKle2RnpOPehed+8PCvIBmWeh86VoUV6xjta9HYQD/0P1
der4uC3wzeLMg3do8vnpoj9IsRCpKvpBJX4ymbSdQuOZaqHGabUlOVqee0N1jPCO3dszBhOKbdzH
GdQcGY0Jd95lXIFVTanIcf1bYTTAZKayDZEKfXSxFRcRC3p7umbtlzBKdhJtFdFe4bI1GFgScz4q
xKvWfxLTC8d2c7cpNTZaE9n7Z7te+a78SWEByLhr0CJppIIMQZxitH1F//9rff2+AhSfnx6+0VJM
HBY2siCkhXUp9auKzgqMj209zT72KxfsYqyeMk9K5749Jhr/SkECx23qbBFURvx74ysBNow/Gy+J
HBXI49iLSbqd+9Ut25ussS7uv8ON4pAPAUg3fiCqUE+sNgGoCokoGmCEJgJUOZkwAwnZqFg4Ob5Q
jaNvJjZ6hLIRkEcvTdh2FdWNb9rzW9R9wVEedEWpMXlf4h+LxweSpvV5IqqXWfbsNEbdyMk5OmkQ
1Lum/q3CGmen21epjdB17DaHgFhjJmw3bzNlZA6mf/1/URRVad6HwHJOvvDlaugMNLi5PC6wYPHl
5SPPodpW0pJUelUUx98Xf8LYvdYOuOSqeI3d246KqZslJ8ek3HWQyDDoexCy3Ymp0wEly6gL0Nzx
AMCnm1cLEfTbAiPuTZEIvQ/jbDrEo15xpxrBeGvf7YAq9BXluk9Atno3F2lUWbvU9BOMjVYMIzD8
TiLHbO002p+blnTWrC4BisZPTCjAf2lIVQnZH+fzsFa4bv+01aKtawqvJc1lFJ4R08hFu8+sjSTb
UYeFouyNHCk6zSxxt/1Ur2Ff12GfLoNkiWyMdJ+XwCxrEUWrxjJuQGMU7FhZfgsiJmer2WW4r8hr
3jwttiepLpbuJkUyYTD1p1sthBaHx1MXOTRpA30Aen/blf2tUxAczC/RhYRUf5IpvySp02bpr/tM
eh2w6FE5Rkcm96qFJqaU7qVMth3wuAL7O7V6Id9VtZuNnMeRfYjKRbrbCe0OvuxS5lGcJV2i3A25
4RHswqEBoIwFZFUHxQiRtWuiUGxYsS55f9BeFmtiTnqsNp1EJ8qcv2uQBlrsRhb3CmBs8imF34qq
YUg1rLDr0GR1/jxTCdWY6+wkSVHFXdxyvN2V4PYmB5xpXpyaabLG51FXOHXpPUFl040NCkNu0oru
PmpKHRMQKCn9Iw03T/auqkgOC0eR5jIbi0hWPJoLrwFLIwlpcc5KpzCuAMX/TGl+ywd30n4t2ojO
I/QeSwZOx2nSiiSgygvhHGI26H3K5n18MzpJ81LeSA/Cw7BQbSdsnYHlGzLCJKropHAyDfu3H+Ty
vTCHaLbv2+l+iOtcdVVwzpSPjoEnJmTbnVAg/9MHvttfkmnPgTL76kVvTKB0Sw4YFIAnOZazbpTq
3RNtiQjW1DJa1yZc40EoawQZFpSrVpFiFlaIfJbntHbN3snOgeSIcNniuD8+/MyaT+AwErLNH3aY
kebQHnn1QUnOd13+yKiGSfKzadh0jqj/0t4054wUeUCJZFjlpMpHLcUDL6ejNRtzTnhPASLtMdJF
kXKj9dq6NWKN4tvq+vDCC3JhvkD81/gqtkDMCnmeAAbCp9xJFtVCxKl31ru8aBM7gez1lw3Ffgs2
BuFQwswZWGPoJxlFOVdwyZDmmUyGFwIOc5/CINJ/Oy3134mdgBgDCLj8ZNzr6e95eSwCTcLARBen
mz4FQwjL+s6cmBCmfCPoLepNGc0otAn1AzoLFipm7c9pZUbRGeL4jNNz7hTcY7igor7JOXTgwkTL
kP/9QeLBtkrijwYz3wnDdCqNxhXruocaKsoD5/eNsmvFvLG6LEeDRh8xewOAMkjqkbw5thvUbNJ7
4GRUb7Yblv4WNz/Vh2CFJqCkXk0Ezho/qraDBhOO5pWIXzFHVASEYxS1Cb+QtI+zkpHrIKmKyJFc
xfs6MJP9Ehhlp0K2H25SV9fMVXi88WXxmS5M7P7999NenDVx6xoJRItqzKlDoSMuc2MS2HtopIKc
adlR0XWEOPeEuZr21Tpv6hwSuyTDKKjkXAX/iewiNR4hsstD70EgJ0zFW6K6hpHQcfJvFWGNYWA8
IbX13Z1GnAT0HBFFogSu+yV28ncZYo4+K7jFDWB2FEjnlJLPEEfOEryhbphs1XHnr2lup55s+czz
WJQUv+SwkmId5zkAbSkOZMQso45hK/08Y9MLeavTVO52MM21i7wYn9GMwg9ZrC6MUvkGjFyL+w+h
yh4bmbLjSNE8bsrpQK2V4J73LvX0zxxAaOpmF9OOpkEyjqRGMlwplzYr6m1VYPUd2q/Pevhm93wo
fkyLhL7jUbzO1FDetsxspS0n3E2x+ryOJopHNa2OMuFk1aAzvuwvVOdqnoaEwnshnaOh9wjtHk3S
ktwSET1waRc9vDutvTadhIcopheiHXRtkiyPZfDWr4ve10UdckhT0QXqxMjOLvp/hOT3b/H36uwQ
OeT0ZIo6Q1lsQXKMIfP9lHxYeMmqgGIT40V/yUcaeFtAX2iRyGGmQTIwjjHMwPaIItenK5gvB2L+
pnV19oVE7887Wp9LyPZ4TN5Jo9VL+JXVwISQwYwzUj0+hUH3hoSv7SgzTrc3sPdBCfb47jjxkCbR
rK+Fh8xMQvKOuWJchUavAoOZAdky7RO/uv4h5DyHF/hofXn3O1TIcooGHnuMpjse93xGUDF+cjDV
txDQs91KS8s/D++R3gMpSlybHmr8HiQtymvSnlXv+pCeuEcHeV6D/mFvEkGNuSeGkHccIeTg/2uD
5psE3aTefKUt+qdBdiGVrsczYhUTGqMoBQfiiy/29Vm/pV1fx9KH6dSzpkSRbHUgCPojoAMuTIcw
hfgARPYhLuE8eTzhLYh4xHXh2L3oeF2xKWg16V2DPn8STD5LxJReU+EM0dLf7CTRgvInEU9aOKu2
uXlNMKGBjiLLDn9fQHb3tS2QBHInN8JV0CdKdd692/TjpADmv0nR308r5uhYqX3Gn4qZn5kGDZky
AiU/UxJ3z95dT0GW7UXUW4G19ABo3FtT02JdeTUS6O3IAZ37PI8pc7WcN6aW9ECRD5fqnwS5bX0L
Z3EzBe1i1VehOdt2WfMrnNAlVxDHRJkLfr3g+KjMW06sQErl+aVDWF7q03DloigzOuC2yP8arXfU
U+E0hgZ20RMb3Tw0Tc8BnyV3gE1+m+dys6WvFEA6kzgnluiAcH7GAY+ONVlPuIObYbRMwWjpvAFA
Z/Wq+Dfq1CWB/WurnZVLyMN1NZcv+yblks0F52Cp/svC5AX+IKBRFYqSM1I4cfg+TKxpJZQVKMO0
L15NISbBoIgpCuvzFgLXj3SOWsbCe724AEy82iF/jXNLYujfslI5HzezIVKnKiJXbzRLHkIqzPJh
ebHkG6JmtOaFWbeBXaVLdp7VA/yPmx2yZjS1dEF7yxljwDKIGTKH8Bm9wILbxkWkuFDG3dmBHvdl
6IjFrgqrx8v7L+6t6X928kGnwpCM8aLIoIGqkmvCR73GYGNznI90X31bTfuwV0RSHk92w0+TtsJ7
xWVnFt9qiSinruAMLRKFyZ36O1AITUAXRX+iH4k1GylhN057LYq4MBG4yx/QbFenS1TdPXHe/Q+d
z/mbX9W7tAab9/8Qlkx4eelEg0pw+4aA/xg5dSju1cad3u/1RvMdb7I80xfLa7WfOkm/5Q+aEEh0
jI/dd+dToB8jXYniBARI5/nLFI/+uxrXJm61ZE4WO8NsHSGeexZFN3VFXtXxS0CNmaDYPY50bTGZ
6t/90CpytuntN+rTM4f23b8/p3c2Fah+4x4T4ttHYXTzjsNLDUsacBlVolUYq+DkpUbuWtbfPsVl
zpDh/UWb68ohUd1FVrqDkrZoATSWL9L8z8XLuISJHRfQxOGf7cYVlSMcA8fxWfeWuTD8CKBIeUtJ
RU7kzWB34qOsYzevz7rYUVkJaUMMOLTGy2OaHPHCVFUrdknAs3Tqmm7NNpU0kxOjqKo2ed8x1i1W
yKSpLByFJPJcW96LzolZX+foN5Uo5vV9IogxkzaPzl1hjbXQ1LqlLTSqZmtcmsf+X6LkscwkQw8C
2nAtwMjDiDggcZZ2LHxKr9K9nVYTBdI68hvpDcbksFZN368r0kO5CgKnmgF1NkirmkiowndfDqAZ
+69wyeTKbdUak8+UemqBAmOziEuz1VGoyWMBmeCVV/pMKtGkWRwPJpAO8+jsXysMC7EjlF1ARgQ9
PHki4gQGPzfYQvGTYc6T0sFmkwlS+dag1cvR0PQpsSLu+tUleDsNGZPGxjwAdyGQKt0ypvGC5zfz
D7yFhi3sA6+jJ8py9d3rraCdu/8Wn+yKeq/JuQZ7o/P3Cpm+A3swStk69pLgTpkFRu1bykSGc9NG
vn4kHcx14jUHMfxjTJ06RyWi16BFphgW3C/0UjVlYVgexqhz+XiCTPhm6A1Ejm402JlMAnasBP+h
6ye2W/Yb3mrEapmT5GU5qos7HqPwTgdjVJ6uEaJkTQDDlZSeM6mN2+BYiNc6OeEXhVsMnRjSUXxF
YOSAhYz35flXoWkDNs0QFW8YBPm79m4DmOniTdZCOZhhxBOf0Xd2tgFMkKStIGWHpFS6xZElC6XZ
GF7gd1gKy0GRCccINpzGNg7kh7Cc6ImtN8AxmO4EbzHSj0D+iwqEQ2AZd4uHnqm9738YAhAawFKd
EoZPMRmTXgGvPsB3VpsF/9WuOxdiUXeZCa41YTxOBKdbig/RhqJumLTi02LHj8z+9IUYCP1AKWdE
hMiSkRr0++Gq4KjCy7X/3yBlhMYnr8yLpOl3tUB8nLI8wWKw1c1pgLu1ynoCbm9uJoXy7tNdH3gt
je17o5xWxMcoI6cREOG9EeGp7Yit0p4Ul5DoDyA7KyZSCk3+CPQBtHcM7d1v/WHV2+t/JsQAyZIK
cZYnVp6P41x2VKdbn2IOQ4ok8Y0TRzm9XnzcCQB0CBKvmnWpImAyrlo+wjafKPBPGxUtI+0gw2Fh
nY0nBEZaaxqVVGIXAnJG93Ht71XPZSMgKjCfWrTMEbaIvLpeJy7MpIdAwGFTGs2KUSiFpGfJ8qxB
udONZkaGykkfHL5SgksCe/yAVazGGU8LJbEAwD3VkCmJY84y7QFqNH/9H0ef0vaI7drv6dHQ3/fI
eXrtRrFlRp9u19AG+tdobmQ4CinvaIBc4wom/3UaeRWCbqK2hcK4dELheuiLek4QD/c/8m7+Nmko
OADqygTLeNUAY3bVK5UT5fEJWRoRWGjvvDm3RvaJdMpD5HLuzeVHTQOMNdCXOqbgF7j2CL9A4U0b
PHmKuvKyo8V6t+sBxfsyO0aamSrN7x7tK3V6rHGQqcZubFjq9pCKag0iWUGXMgTJQPXVCL5gji9J
vpy3+eN5sRX4KetWyZaj0rtYLsXsNcgwZ/tObBFVOLKt0jPCixfVZWirs7Aaop8o5jqTsavULS6A
Nx6w967L3t2bilLQxqVGbXlvCtPTZDXAF5LYQQdLaxjId2Dr4tipyskHDfP0mF1UL0a4+ai8o9/5
GSHRS5Vmhr8r+mTGl86KQ+gSGhCSCEz8KYYAhBQxSofamsAzJFygW/VpGjZOQZSHOI6oU6c72PWj
wwCvIXvjTtIm2/U/0K/y3MqmmouXhmeVIvcVKH4fEYjRfAenNZ8N6CyLYQGXZ8EoQ7cUUwA9YGdz
hnBBDLuVB3oysCD39BSC44Blis7OXeW8BDTfqwZ7lemqDIYVsXZ4eOL8ZYmyk1vC9iUG7BZZ3iUY
zW5Ng/O+E5uOcOU06tloFJw/CPRRm30PWDhx6STuLpzn8iC0tMOPXpw073bZL3ljN8LC8hO6O4gC
w67zfQ20c+wOJqL+wxFGH+Sh/fR8G7NxNFxrS2Z1BolWR9wIu0K66vEYj1L18TBbSXOQzDz5fmkA
PU2by7L+8joJSSuHAntp1uFKci/UhQmwz36ZQjTPGkmVvtcyb0VneULZt1ZS2CD9IYcC/Yp71Bo4
Y3Z9iQfUUukANSV/zviB3kF6XJ5+1c58mPdJP9mzI6LB9pPs5QJH4FSYfFTdeVrf9xjOJIF281tp
Xb4WauraP6xgZ1Qj0H/qPqVIRrw/jtg6rUabEOYzcfsG1bIPAf6RVbupeYSzmiYGSJgyoxE9p5h+
e+imYiTU/W8Z1LQ+Ee5hkHA+SNmo3oMIZf1CuNrOeL2Mpe2e5pbOqOSoeIUenUBVmcFQpmhqmxdP
Kk/OFTa+R9FI4z9Lt2FVXhtfWTjsjPABHbMC+efcnFBTDrRZX7wD7SZbBwP3v1pKs8lh7mxZdUfZ
rb2Bq9zzh98zPZskWlip9GY8Sumo5lKwPXwVpCE4KssH6/ArmZaRVeeAC58DXC2gHe35ZMnMAt2y
0ulGcEv/vRDMl9UC16e3wOI8NK5o5tt0Zu33kWiZGxlTZUTzrwWoaj+0DMTJOjXR9V+nyn7wgVCX
2Z+Jk3pMSX5AaT0wNrEL9uRiU6QGQtJyckbiSRra3QTQCsCVC7MEguW9uQVkEjdtmXfFmr0aOKLq
LbbMbKwWNvWFTdhrrABPZmoBH3Thjsf2afGd7sTWRpITrwlAzV4OckHXj25HMJaq2T4vVnKbcD0Q
+ai1KPgnWXGfZa7Ap7DOsEBl53SjfFlba03m3Z41RmWXNYpCn+OIJNhH6BiVsR6UzUAZK2hW25Yx
wKxwLJqpLlfNmL7ZVCJ8thdc05jjHcctfJKTZlOiAsyaqa29oX2cMIlg1kGM6wlFagGCAgPkrvir
6ODt1wh/pkaxahHbt9c9LHBDk6LwrUjkrBPlZvxQqFiiWy1RXlJ8+z6HWlV3CMjQTJLhR/+4u7XO
tb/62Kw00UMRqPlra1num4FdR+uU+FxEvGtA1hNrTCLl/cjbx9nCVIo2PRYIW5GcPRWA/SLYL75z
Y+fxnLhsegkH4gLdL3z/9v+ldfqLopqa38ff1+GsVTUbAPSWrp95abHZt2BCokKtPCcbnZtTQqdV
yi/1LZzFaWbPj3Zka+HyJfHrFIxco6P/9W67ELqltRsGdvP+qQdW2zH4k4XQhm6QUyZNRNz/RY2/
aDiQxkokqcCLoQt8A1DEz0ZQBGTTKz21wbW8EwNJaFUSY9aXqhzD6vxr/3acFmBo1uZSazjGRsdH
o9eB8M14K/C8ar/VseMsS2qOSEF6hpixomXHsuvNh92bLhDIBjyql9uEOhfbohW1tfgaj+M11cHt
G0Gior59zrio4OtO51fPsPA+3VRJiI6Q/tzRNJ3h4BMfC2bawSxcRnrNOatV1KbKG+RyoK9IOpum
rEbJZl1ljJkia2uzoaUflGR2eKzgBne9YXgv5U4Hq2rDItTMiBvqgiXGt/FG7vsan7UqdDVSfiTC
m8+CyoJYMsR1CLtwQP4aB9l3b5uzVUmdOFxNjbUI5yDy5VROUuhgiP6W0pB5iOnuvCYEqSUa/VZj
kLBReBrohFPFFPo67gr2sk2C8M8Kz0khPdOdt08e48dflwEZLgQTzhUNW/SohM9s3eh9rI3igfTm
aGiLuaopfnqzcxCaP2ihcuZU9O/IfrTPzkBY3SBfk4ZcoZWr1VVfpKUiTRUqvD4qqvlgRZ3c8PWE
S69jRLz6jnFTN46zJxWqaYVawjU3J+56PfYBKwOFfLhisAP3mBO6T2BTaCOPOM8AaKlL/2UxsYdh
2pN/V425lY1eRgIMZzTYMin36gH0YCYRoVOvc3i3mL06AsH4JDKFUowtLAfrA3ohApTeMJV5heEu
lbQzzjSZxWrt9N4UCxwq3QNd4j4HLCcgvYs8BDbwkh+lzgPQtlt4ZSEhmbDNENpXgNFMr9rSF/PO
rBWeTKRMEeZyH2yboVCFxePhi4WjoC58nf8IDmqX3t3QXbfNfQKyfMToOeRuk3xw9lVZ7PhirqN+
bgdKO69pzCKYrihPtpQFdZQX2xpJQp3MQuAEynVBOgKIrPO+kY1uz5x9gm7BQL/kVrBeVyDwsj6S
0LVd+lg9JUOglPeu+wl4x3CbGldyzfCw5JRjKalg7xnSOkXUq7AmyLplLm3YfxOPqAH0FtU60nHa
IN4y7QhYaoDOd5t+H7STTNPExlZ7cvAQGF7GAzMwbq+X5tosREv+4F4WvFwxe2kTrjKTxc92AFBo
Nx4oaqboV2KEU+aZ8TgwsuggVTRqUN/m6jAE2GCNXNzI9INwYrrZE1gGllSzRCxXcue3NtVWMkHf
K+uqV3j4Zu+rvhdOa9OBNtH6q4r24A8flG3hIB1qW526JeTX+14ZpwHAIHWKcyA+QgtaoaTqft0F
iwe0lkcrVkRzjeUIB6qaBvi+XI40X3vErvIdx6D+wUmtiLZytYZzRzJntDUfrrudzPwwstc0yJwQ
+0N+QS7wCz3V8tmLuibP4x0rVMXF3HU6v2NvT7qo4jtk0mUFHeBQuG1zuIvp+4Uw4pZGACMO4cfD
nyJBVOTNyg7sKni0D2vq9HkOt4MhuilEBh5NjIN9EcdPU43WHxYvR6lTNOBRMeZEIhUor6F1sWmQ
uYgP4o+NyRczJeRTVt6N3u7juCYSl5wZdGDfadNPMqoPKgBEucq7S9vGpqu/7hG8ou+K+S8TL+fC
1s8mmIINdb63zHJmIvMqvZrjzRMyJNFhakP6op8Da/hvdTywizfMGvRhh516K+GC0mYjaQEtt0vG
fKdUwTtrMVZJz77eSDKK6c4q3b2MFxQEa6lC6bFVleqjTg8z8Jr4RJZGwXzd470IGcNaGmk3yfKX
xr3VmI44SoCE6FJgLfgJbMQv7AmxwF7xxFotWtPOsdonj8S5PQpyXKnGQ6RWW0cQp7wEdShnR8ch
FOSEk/jtgjNwpoqHgpivDQ8IJkfMWTAT8rKJgdiwqSe5njZL9Px7vYv3/86vK2BKUhyawfsiUf9F
fl1t+eWO1zY+HIv1f8f9HH7+VtLSMMtWNBnzkSF4cwcpGmJFPK1vAbq1JS1gB0AOvYVgjPXPnoF4
o0V7zJY7rEwexXPsYEr341Ham+PKQmC4Krn+BaQs+7cUVxiZOGMDL/MUyq9KvAnNjlWq9YbrVHvv
o6lY6Wvxxmuo6PW63sO/gX9yyX0m1F7wEGgb2VEFVKkNBxdJkQgHZUQDX5zuWNOOcqhQDyAU4k04
oFrXX8JPdtoFq/noXoZuUlhBS4ZYdEbgnEvwsvNBaiPgeqvDLvTxwo0pSjWmotBq+H0JH6Ev7tkY
mBwIr/W0JQwgAO8ykjkZXP+VZn+L/0lEB9hbcdePg1YPFFeW604HzwdT3A5jHa87cxa5/MbfnuEE
RKX/2FDZzPIrXBZySKua3tCsBxLdvMxp8Y8oNbF7bmfwIQleKm04rsWNqgbO82IRLbUlARjhB+/a
SbQDLptAT3HqoxUtFffVMLUGBu/7fBy4XKPTUIwZ+JBHp3esn88l7P9o7cOkM7H7AJHxsgWhM/O1
JMJvwp3QvNWiyiv2bLpu8LLysSXXPFawiznVSy95WywGMa9Sr9tAr7BWrVlq8KKyVFauk/QO7+hQ
ojpKmheHfXqw+e68T3n2HBkR4NoRcnB0oA3QwbQKkIVg5fe1YQZw11ViyNnMlEE5jGxHGgzW1VE6
j5uI+9HuM4hZhbpMhnpfGidvnS0/QOdojhvy0vLUUzi+tSJg7JbRiYlHLYKhmTjf/1A6WHCMSisj
XEdnbyWyCtZXhTjGVjIf03fuzCO9HlOB0hA1QOTmp8C3KBjTWJ1uQS53tSMk/6vUWwMLW4zYGuLh
vOIN4QpbKAaIyUh8fuwQtclZKldRCow0MCcUt8o4HqN+XCAz/PigQwsUw6YsQYAhm5IV3cPDfqMn
WtkSNo68MC26LKCCF3gHrRcXhJhpBhSQSSCKfWUc3Vqs4hMB0bB+mhYgdwQuiBn73EMJFpXd8hyO
uQGzXE1NMp2nb/sriWettaBKS3mdwLNTXCJB+wHSo2B4CFXKRDMXUKstIepdtGjS4nahIf9txaiN
LITWvKZv1rESCjyJ/3bmHHr6VLhQe9pa2QkrYQ0aFcU4lXNeSZdRJwtkILvQIP/+NGVhvBjPNZhb
ncjI7IcNwdy5x5kLgFINMsYO1Dj55lTM1GaPF5x0h5IT2T4iKXL0+KD/TFcYQx7PneR35LbQxKar
64wNHdu8/4/k1eLbfZJZs26QgWhnPvv9rVwi5kH24eAzZKWH6aAq+Jgs7Bwfj77ftRZRzsAu53Yl
372vIuoNAXoXbU3//I2NCzayL0bThy0Suv/2e4XK3im0OvF340ab3tFxukonBsUvkaY0BOSEVIOw
/fQKL2g4KTm35OGwShXFOFa/xoRCIuYlGXq5Iwhh57LnOC1hGhBNBUaKk+VCpQtvWCbuzQmJZ5/C
R6iNG8YZPXED8ljqudLWDVHkjqE6A2mimWgtVqBT5DbHR3iTfRP7NC3sj52aZnWwGOEHZCH/vHQD
Nfn3jrBSBAto5SFapd0ER6+HOM/Y0HpOzcV5Bg7aKlfM2J1j6XfvBB9qyHpKp0AEVejQoUeu5GeA
PeXot4jUU4wLEqr85NqibNWW5QWs9XDl5Gu2w0voYjKO7J+oC/XLsk3pfodS7B2s37cVnBIDhhB7
MzZUumYga9Ei8zO3N4U5t74Q6x24AV5YhJp12C5GAIyScntqERy03P8iri0La9kJbajzkT3k25Jg
Igb27DpxJgMfbqOrg83cWeatzS0kEZH6v6T7ATAC5el8Z4y0xEkbjEG7zRPJD3voPa8THcD+f2Nt
gcB9gDk4InlBfycAuPpSR/ZWr32qRPRfQJim8/5Wpbe0uIXp1wIEgnja47c3EobI+8jrUUDOog1L
rCe2vDwBAhvuKqkCYKMhjmMB3dSucgnPH3Xwy/QsV3SJliS/16HJNbjNoq8NGq0y56OemxEnfRBH
KeP//UMp1xUxsn+1pd1aBt/q0heOTJRfsbaKhjWkuJ2cAHXo/AiQz9yHwViT/ga3YziU/VE7mOHP
Qkfp02x90nASpronbDwQ+cfToWN5gwbOrVzdvD/OSxUZEdZT4UNOtmBdhOwAL2lZsbWIDClKZdPr
FWiDLhjpqMijvZEJk+l4W//pWNHFzPQg2Ql1h5advT2nn8+i3FYYMzXkQnbWvEhPxJpHRmR64Nrk
0IU1suFg3tHNm4GFwCB0EWwSVnBessTO5BRCCG6zKBpAq3KnZl6N8y2WLfjMEUhlHSq9e8kAQosr
IW6Tl5Wx4WR9EF1FTCIcvu3rHqIrQtyWQg5kq1Uv6Ks5svGcs9Uu/DOzaozHb51w+m0MJfDY78PR
rTska/Az34R5H5lISSCntUhqlvzKnBhSKRYSwuIWJ09axgvmaI3w1T53CiA1zB5eWiFglvM4q47t
MQjQ1T199qZV7lAta9ciuYvvZoxJ83yDSQoRX/FgCEdIW3XYH8YYmzHtSCiWpe5J1IANxDaTbvs5
eOkQEsJgBYrL4W+IzPN+qIvMmtI46dA2wIw+B5ays/bLSPNihHR6WwJNgfPhjnOlOV0gDh6vPcUs
UupdckzprswIxLJUa2h/rYpEMB7ARW5y1C8hu84MzvavxX8On9A3Ud2YPT/OCkjuhHWt/8dFjQJS
b2EvHgw3HlIW9t0teRDlbjGVkWdrwrBNVQ29sSPHba5OBTeWsg2NEBtnS7zd6WiTXXsSBpitB7Fi
lPQIVARcWxrfH4Uw4g8VVvGkz2PZ9iFzehjliFI3XmkkONVevptAqObXkkeOLX3o5aES0qz1ycPH
lpADM7Bf7IHaoqGnLzFrptArjP5AattnZVM1xzWeB2XGGgZPN5O9LIQgWB5U+3E8T0tOQ3vO3A0a
449/0a+46u0xFjws1qT/Rq96KtCtnr6WHDgp6lYhVqTCQlnPTKBx5JIR6ANF5JVN6Bh+YA+baXms
6su7M5aWM3V2aXCNGlXwhhhMqwbN7tnYIfXnApfVj8tJ2bRriGei9QmtKnyFRufnAYXL5N1v5JPI
UJW4A3fhBeE34xKV4P4AVa26+4vjWT3t9YQGLjV0dGeVrNWXkmrgKjSiPTGHXKEUojXrW0YXy9nv
Jo4yNcQjrAybeuKLYDBCvrkZ8CX887AmMceJRrZjrxpQyVaM+Sn6g9C0r3DIHp7oAwwdxVkbxlU3
x2zrzmmAWAGr1flGqhkg7Ug+ssGXmi9w89LAr2kiEIDDpVkwVGuRbRJMZhy3MAIdrYDFk/v1BZQx
7N/taJza45+JCTTu8SA0kxtxIDmGAXl0JWdzqKtXpQ2LPwpyR7pOa20Q8UuN4EINQkGyyWf1b5vQ
aR1Ku3pDaPFpewzjK4uLNomMvAh0Vn7RiRjZVVCmryk4xno0gLckYKXTMI6zbnYwsU1axoyif4mu
isasrckYkKy7dNDm1y+dCjdUH5r1tISuNgil7fXQ1fH+j3d7GXjRwEt97i1MxGZ4GAo8Dbub4JFx
8mdrSF2lRNVcKVswbah7y6h8dhI7xoqPfQbihyt4pFM7p+sBMmBn3za4EwZdQVBHouiN1NAJ3dGX
ufhiKowlPPzmiQWwAsNSWBjP6CU9aOqyzfuCAu/dfIAW8JDlUdTX5Bmjy9mwzotC3niv34m27xvI
so1HWDIARN2a80tYkLm4GgpVaXgftCCUm45rOwBtMhSjYCwzevG30YpEKlG2nbwfvquX3PKKnM4x
ZLT1oi14uSp/BKACGHj2B6E9O8jD6xt9CF5D67B5KGrhyYprILjeH/lGDEHOQYKlGfkXUQHhAqGH
vZ0ocitqWHP1DKYJgj3/r6U3EB7gXmEQWbFpicAxO9SKB5eyVWsga1AwodYUWHh7xvOEeYex/OfP
rEhwF94Tb0UIZV1h79A/Qp3b+YlVdcKq0ZMAlcZtGzLT00s+Im1FVq1suYDhlSZihwgLJEB8R48+
TwbmxyxpsQlnQswUW9b28WBOja6PuAHBt/EMUF3Xeh+xxnswFQqNB8gZiMDOY0eocEw9SR7J4HuT
Qe6OzJ6baqy+iftYlxmbJ9se8Gkwt4AxzvRKmyj7dtWSivfSczBuPwCBAPFrpR2UG3qTZpgIGvNc
FJB/lQPJ0CjvunmApTuNXJXBgsS97Un9ghHE8svhOn6Pw6yUCf9klBKZck5Fxp6nxN/ngQ4FLA4u
y7a1Y0qyJdJVwdYgh8lxE7ADr0v5PJXuXPQM/4Uclqlnne0ngeutI9K18Dslrj55c5KAASx2DIo9
/zh9JWvwzEWj1NMfwbkDu8277i6ueHgPU4YL3viAazlnA2hDdJVs6ubHW+D2/K74BdNngjZR4MeP
wLD2307qLlcTl3NG/ZRtfr0IReF28tQuNG74pISxR+07PwFl4ooFULrERWJ9/zSlCEN2gjOcVQSL
iMXQqKYcr2rtLV9VufvXQZNJrmynGO4qzDxN07KqL8+sEylthQZCdYb4515FlhcG7Dokgvug5tFT
+ZBphiNJD3BD+/pnnLofnrt8FDtG809SjEZnCIH/Jv9ybFELKYDETjD4RJeWmG5OQaCuEBbKRyu1
XqI+uCX4bh0mj3WM/zB5XFWUr47XO53JTJ56NphUfi+cZaHSFJoGIyjdwADH6wYjw+/KyISaq23x
YxovUtZHzTbTH2J+bJ3jzE0QtOzA1iBYo4Qdairaqt2ZarI6CPCB6YsuWdu8Yl5Wmja9tVQ1FYEL
f3Mva8QfWRB82BR4itq6mtEhcn+6g5duyLQ1TSps+mcLGo5g2mUlEB2bKrjz0gs2VYfWr0SjTYKy
JJQla62yr25ckeLSmXd+EV9ttVctYsd7ZF9vgLzdfwyIg2H9yqLWH/Lo6rDmhrTdYwQejcjw5Z3E
DSboYUnvFVx6bfPFCNM93B9aC39B7VV3uzVHlpqzvaKRamL8Gswk+E+O58fT3YEOZwMliQrw5EkJ
w7SAptwNEFX0/yczZqYE33dATG5rxpZGgsU87EpgE9EbVUppCWTLjW/dFZE9Oxi672QYwvLtslRh
/Av1tMcvNZWEgAf+oxtdHyO7lmPQ5Ikp6rWgb7ot+rr09ANeogJqhozSWTbajKxWdO//CBPpWCyc
pfB+4UzaVBqAADRCIZ5PbEt7r4d3Srw4JHp1yEOXg8MNI5O5/TDv9DTuYMfwmLB3QPibXKfOJ8ha
EbOChMlq3cAkyPvw3S4SH4dffbbF665PTc0vM1lN5+oBEPJ4AjEOoaIo9e74MiUyEMy+f0DrH3/9
lyUv/e+5nK7RRAfoYUROibQ0nvXNkYTs36DjJlPi1ODtVg3qksxIk4PmzfmalwrR2wHnI8JSuJvs
lxqMm9KVW93ydHdKzfL/nMvl79z10Sd2lbCnQxvxlZNrG7ag9abjxxeGQ7rWsi+lL3nR9lXQUXrc
efatTmE27HeRngFwj/wnVg0m9Xfn1ZOYsRiWj1bCoBgkyayxmlIzqCJZJmpn3zdZAnrycAj3kQ4j
qKgKObF9c626Xe79H/YpvVGd3cn5Pkdiu9jiL+1/rmpX0ZCrybtHMggG9dVYlNcVApbke3A/R3/5
kCQI38xXZ1cxQtmZEtB8gAOBQRmivS6lC+XFXVtRUlKgFQ3RTlmvjlmVYkgTaDGsX52n3XPVIETg
M307DgmAntOVVeKuGjFHmhWYUy3fEZIVDhr/7/DSQcAaXuSvVXx3NCZJhtx50pO6NiH6g2OVrFvh
k4mTTfPTdphBX7+xHi/WW+HKGhYPMx40/jUKajIZfsmb63Xg+HuYt5pee0db/k4I85odWew/Yw/X
gHb6yH4USf1MaqkN14afRvqmSjxF+DP0soCvtYMfKTF/tn5Btu7OTng8uX8/b+xO02y9NKW70jc3
vWKtVwvR1/SS0BOIZn3s71LbHvm5/9QUdRXAGBUF3Qy36lv124RGXV2PEgDqJ0GvUtKzEyD5dQg8
zYeacO1BjjbzV/XRvxz1Ls5vhTMTXeeqTOCJ7JEUElvH3qPSIza0bMm38dfcCnZRytjFg0aLhfF9
E1kUoJ2UQJnc5Q6M+bwhGTfdxv9D7TPemXjafr94cj6M5SBphP2yFSU/M6qSZS70hpd/3s+fFrmy
Fs94hwjolQU3svPa3JPomZ+EZiw0R9zCrZdEQQ5mbgPexwIEHeEnUgVGmDR/wQPUtR+DgWSrSqGt
YaxnytiEm0yZBGBwvzdoHX1fzloCJbiAEQuqJ+asLdq3RtU4EnqkNsEbk9AbX4WqDcUFxBUNcHQO
Dh7vXJrzsE5BKHicN1XDhBYW+xb6rSvjT2gFuLaxfIWihB/1a4RMZHTxRaSnKpAxMXIkC8iMwjou
W+J0cyD2ms2XBVxDeUM0vO2ND/IE6oJciTp2r/LQS8c1gWIm7mZDhTyTkrso9DUV8igqyKoH98sN
goW/Vo8eevZTKZXwDdc9fxLmbzWlcc+fLD2Exy3hNcvnUf05idsxxxdhUPQjJu4zgd1MX1atKAHb
fCafSIG65TVvF/Bz/r2TJCzUevLGdJBoUcDpTlze8z0q4XSaL2fyd4EJH+LzE0S8Zici864Tm6KD
GSYttkPfFT8UoyaEPyEc4jeS4eL1313b0441TSdq+phXtLgOJmQFlo+jhcyEFCoppwhY8cZPOdmZ
mwCjHkhJ/dVNJWucWOY014/ADPHv57QlG9dskDfVC8cUeAIbFnm6WFKOv96oXIOXrgoTdMfuZuO2
i2WFDQOXZZQf/YBDYLjGaAuOEQF9jI8e+xqDMZeYAGkPQcQvtfwGPjt1f9TGijqxHOQCdo0PS0ZP
NRTNXc+9l0qqpMzj8CfUwkKNQ36xt217d4Zyyu6zpYk4TLdiMC77c3oxF3wBC6zjX7GqOVA3NARZ
I1S6q2f8WrkAIaCCtyDXgaBLRVIjCR/jf1LMfO4KEOQwMF/nSqYAPc3u/KqbGKTgnADxeYP2eTGk
+S+40XCZVcJ/41MxdZImzW6vmc/ugydYcosjBdnaMsXvSNZHgRD9eVktv8LBirJzOuh5KvEaTHMi
O7BNqy9askbXlHZFnU3Mm32C0teL/9w/vV7cdtFSDG1PyXjhv958O9PPUCJrvbL5XzKT3aVeLmMB
9vUodghUaKkfbfH8r1/m8OUHm2w3FL7UKyvhr+L0H0n89lr03nXNZaVTm52Zokfu7NiN8RZKMqZL
MOFnOA3jzAq7PcOAzTtrwus91Cf4/mjdBYaJeFTrLLJ/pBWuALBqwiT3L14xhSQJq5j8pgl/Ia51
agjZvSS2RI4m52lnZDqL80MAndrIqbtiXQbwh+7GU620GXyy3GxFgB5H/7NaOLYElUVbDPDI7rxy
j4PEycOW9D7/rLUqCrpdPh0TAKf1e5S/mfvvIT8Au4ML0yJERnMEc3UQrTngkimgg2AgeCV7PotU
5uj9TeRrFAccc2X+kDNbUBbEpM5TIE4yVODOdvFTav6hGOU5e/EbIy1i1xkauc1V0KUGjyQtCP4F
QaPEN8O4qiBRl0ktvdEVzrb2r+qQag8PLwmKabNFQFz8Pa8eHStU/iHMHN/glhE/uRGxIx/RYx4W
tnGXo2Bqaa5tSO1GY3xP1PrNNnp69mHMKAoiTTkd+w1SmGP8kXPNgHwT9cXVRQ590hOATt/UDSIQ
/tgDiRESukWKE01FEhahDRnc0q76Qor7XQ1w1uJ6n+X2MRBBswciPLMpzzlezbMvSpaxflYWZHOF
slxzjOwgI4tnJionUE8BFaKff4RHON1cYv2g5t+gnoQCMLEwcQFr6FmBBuwLUu8gblkMBg0Pv+MG
MG9StE1tP5cbLaz4R5B3Q+M84Pj5czmeSKC2/K4N/hR38ozDnfZHon9nXCOX3oinThaicmXl3Ycg
Sg0SYR1vo6rH29PM90g8OdPg38hYXoKBWysHWQa5NW0/4P/GgdYUsWyVq7W39jJf9gEW6Pze+/Uq
ZiG58MddmTwBKGehdSj+e5zaB1+/vtdj4qk25XQgw1uMIghdlyvLAi6EnlpbDQLeQHm/eB9T8RpW
HhQNMrj+T+JBVBAw73yCRmtCVqnkSwPmNXXODBocs+71DhNDRqdOhJxvU+qfHGf1icVddcaayRL4
cZ2r/c+LSVZDeVclUYZEJghqpCpS+aLmsTQnWfP3HahKuZkIYTld3YNnRXI4XO1EIps96agxO8cj
miN6XtiLXoTteOGsJcPzXuBiXEx+Y7WcQx4cgt3bPfBwS8c0UD3U4B9XshEnlBrEeXJt/9tIf/cq
uvdcgDHm99kEBso0ACO1Fwuw03TuYnos8htKxDL79XSMJDC6TT/n9cmRUqYw4NtrTAM7vblc/ouN
F9nLK+F+t5Sw+m8PApmCwA/nOudZPuBjaGq5OgVFzeQWh2agv8XL3BIIqFXFHj64I/Ok/98k1+dU
KK36lOgu7xcP2MPMctjf7ECM1mBeOj6L0htaCCPkj+OKGVY6TChr3+TTq7gN/E1Suq5AEErWhSIT
wUxFk75KGHfF/pga7H5J0w4j8bxTCfvKWYiq5fGHqs0mjc/bnfKMBpIfSRxP5SKDWhhz3/ckeBjT
5TZeS4n+kOX5+2Kcellpn+S7WA2jcLL4q8JdBM50r2UhbRulSRETXiY0/b2a34wJGPzdMtNvacoX
saBpAlS0cU3F3n7Uhqt7E3scLhnChpey05hnWPUzrGNyVHvhz892hXmsl5UTuFKFFZ0+ys0vfsF0
Z/7aaxCx4XhJ5ndR7OCL6kgvzd9sC3x970S+FS9ZvsFuWJgVpX7rOpkU7931/m3UrxPNBxCCZtlq
BDcLTjkSlVzOAvrqT1fzniSBw/KmHeMOr2fIUogeek8nFwoH/AxEtRHF0BET9F1aS7MIX9+2xVAG
ULNDYUICXbMYmZg9LEOxRhJx0sZHo7t0x6BYAzrlRti4zsjwUdJJgP7F8BlY6Wu/+C9UnyU3c7Vi
BtrPIUfnMiltqU4LvtQugc3J2K4UJoTTw1X9mda+dhllo82/wUX2ufW2UfIDGHG3KP36zvuVgzKo
euOaps0Kx8c3odmmmuw609uwBUPO3G95ovb2U1eEBF6OzMWNFHYkrEN68ZAJMomjAGhp5SIlRLI5
DJoJVK3l5yakS/GjRwkzluIaF8f/pIYibHgjfeSsyuTcCu7yqziVSDGrDHHGuTh+i7dubBCEJtHh
EdHoIGB4NpUVcvsfU22ywFbdwUCX7PYgeIQ3wxBXcC3QIKKKv54GprK3P6a1mM3dttphkSmFQr6t
Exd8roiLxenddkF5wMfQ3jwgB+6+u3dggm10T+NA9h6Db7sXvbjDTutSZX583djVPKDrvgSDLAoJ
7LpI4FRdkgurP0VSpg+IVegxFx+WJ9FHn9/d/W5DzNO3Ys0qr0Fpub8lZ0ZZcmQWsEwT6dkIjQ0c
M7nbXwkQka459N3X45VL/9zYlr4jWoaCSckALCLk/VKuMQorvUXrO2E3xhUpdGWSvpHaw1EXmu8t
6A7ISK4B+hPyhuDPeXOslBcbh//zu1Xsnh1ii6XsmxLeVO71inwSnmicSSIEzjNPqQ/yqnARXdmR
vJ3CGFlZb/bWI65LFEZ7DD7p3vrQrC4vzPG4AdKzlfW1zUT8loHDn/ygl8DjLYm3P8rpFIRTY3MG
8bEvijSZE3Jvec6RznKu8tW+Mh9pjxL780l4wtzT/LIeajTeCzSlW/4IRuDPjqlQ33aylWgaDATE
VImlM6J9DUhNleacKBzPlLEB5xMIP5zsruGLfw6HgkaDUOiki8Cb53HcN9Kf6LPyiV4KOP9ua+3a
B7jYM3N7sqnEID0VdJzaiCRnsnyl4K9C6T+iDioiYDCD4+yLj2dPj7BfdE1y2ovxxNsD+XG2UCCX
UxE66zbrwR3fg/E+82eFvq61lYUr2yByOisCU5mN9bVuP1dqD0ZUjEFrOEmiSSd/F8UEeO80EGhD
jskQhEhdrmMNbye4CStRfblphcNT8mDTE4BJNhb+HjsmXwoDTdJG28dER4M2TuEuamS3SzZNoYtw
odGewxBP44Dqxyxwloh1ZHi9vSdUzgxzJh0IIml+cBOhFE1HJ4abyHyd/GGGeauE+ueHqbkZFeIK
c/KcOImBZMxNATxzQjhrKarF0Wr+coTT5/duwSrqTHcgkGZpNdOFe5MD96AxGu/IkAm2urtsJ8kZ
8DFAW0wPN7w5TZyMWyksVzHBChY0/9mMWzjppuCOlJ8CpNhxoMO0lPUcFWw/AEd+yWkkELKxr+j0
4giwyfuW4io7LpuBpr2j6Sm8MSzU0nmmR9S7+GALTFvAA0SJGoOmIRLqTl7x8YJk9FiRZpVt5eix
DZStC7oxOXOQRB2DXGYoyRdPQEFPwFLF/rTX1+8KbfGhs7XzHWPzWUueDeZwGaNW2MqkQec0OhpY
gB+UG8hHeDAc+9J6/6WNoits2dc6ykhDk/I8ezDtd3tESqjKxjG/tSD6raikuhYnNVBBrly5bMnJ
iNE8C46EhXu/5h+7VtjXrylDSpCFRM16u2YrL8ylmpMpp21pn3yvaQ0K85ITTJUgfI2eCjh3itlj
Y/QWb18FOZh4xRIdF1Tp8r/9C7ohKYcUQHdQXdFB0YuPN7Vf1OhtskTjbiobrSaDw769mxMflrhM
JX/7b3HO1QtjVNpbI2o37ytr/c9HSyGmdLlzfPF3wGUE0qwwl05Hx2BR2/OupdETbgdWWI/yeDim
fsiBujRU5wvJ74MTxZfjWaNlQQXx8XVW7auACM6N+ppIowo6fWFzGvog9KwQEoKOlLKOvOSvs0UG
1MMFsUd5zZWRS9ae/xrzOCENBB/RzhtofXoCKwEqlFZqSjEEd1g/9Jo9xNooygZlDT0Vk2oCMwN0
56cFy6+BjJnPiGH7fNegC7Dbs2kyXPwYPKv3mPLfdvbb5H9aWW3JzGrzqqScurVvut30cDna4gjM
SwQTgH2t5y+3u0pEKrL1wywFWPBdQMKyJH7+iEGeRA3xWOI5gjmIb3HgARrUE6Ugdg1Ja4pihkJP
aI0Af7UkieSY692Km0FfxG+vq32o7PjhaCtAvGpK7vE7fnjHp4ih2Jzv/bHvWIM1wNqjxp6n/ezy
NOvVFlL4AHeU+Vs5bm2FtI1iMxms389zIVYNrGEcSHP5fd0SyGAgtdkREOVe5cmOWtgOQT3lH3H7
50dbZLezZnMhPotNr2Q4T/+gA+RJlJP66N9VYXGjR6EHNAOlvOPfbz6q2qC4eLdIs5k91cbH09cs
iw/rsrfKxnyilLwC1X6zsgJLodm6YTzTGlwLkYW/fckVdFzNwrJcAgc5UKH7lhKfaN8f8B4BsQiP
iqX3AN7TgLzj/Mg2fB2qHpkWTYOFsvuI/vjKpKdQxBPDiteYOyivuqj2rvjKF9Ft3/YbeEdrpBtr
E7Hbth63EzIIqbmVhvE3Tn0Rw0y0W0YMIW5DwrElStzwiKI81EGR5JU8QAWUpje0DAy9W88CPqAN
eyclPIBZZmEl1ZiPo6ZtWBW5efIi/ZW4RkEJY8OK+/Vtj4F9nIV8Znhbkshhsk2PUyyCETX0Xrsk
OC2lVgG9ONxsTvTv57VGYCk64oRQusDf0/A45LnWRRiZiFMhoEw09hQ/Q0lc4GKmTZQEAqWnmXU/
skX/UMXb8RnTPBYFXt5GHSWM8l9YLgUxWobelzabtYW5raVIfa+jlTcSlIa141XrNfXiVjeiKaOT
iWbIQmsLRgtLmufCwUJGjX47O4jPR+4FMnPjrP8FogCbRmA9wyUCa/THMvRsGBBbD513QRWNTUQE
M7PUFh07GX4SRut9HjFbRJsOwAIBX3EsNeQBmLELDpx5/N5K/NalGZX+l3RHHPDrUX0oOJyvAaDB
ROIdH17o+G4Pl5pEklncu9wa2/yGuc009p0TSy78ZDV7Le3Tjdaj+AaD1X1imXtqLHt3D+HqdYjh
N/sTC3uMa2bHr2AbbTsuwVoAj6SPegao+KMdIWdduOgw1eNVbPcODGiFuvp1V7aSnnkd9aeZxDMA
BmkCiY6246SF9pW2PUxOcdUdvDgWOrS+eEEeSel65n8iZ+bApq1++rvSXkIGkATrpe1YNnbmeZ4y
C84yQw7FPAdVDq6WSbvYKJPXUbrMSCXLJGBtr97Z3VGNQL87NxaI/kxd/5VTOVBbQMa5mxcHKnlV
tOuI+ATbXasVPpiqrSWr5JarcIiKSD/bvI7giaowpmtM/zJ2j/vnXRA+YEowGTiVDmq+VsjN3d6t
TpYtDONeMK/h2jIs6wzMHi3PHQK+ytR+UHYqcEbSjPntaqpsMaB2BrIqDRXvN/ZtYP5EWd5tAkhc
W4PfKFS9kjqYa8YXPDZ1Ipw2LtkTrIyULf5J2k5KXY3bmx7rqUbEOfSCTiiqjJV/vXK+TK3soS3D
9XulHusYXXTsXVMs44unoXvg8o75CyrBeiCcYkS1A+A7gW9QuMcnEYMqS+DFGEH0iAtEicS34E7V
gRL2L6JEoCCcGYZFFijLOBAMxKaud7mI850VuI8CJ3LRsP1ok8/TeRMiIzQLgBP+Dksp7rL0adwr
iAuA+DHBiS0wnwq4WH4VkGT0JtSqZBH3DQVpmG1moPo0WcywEv9FWP4OEmcTbuhK9O6nbsStQ4h3
Fe2e/GXU/Msq1sxk9kNPe1jEziIZctJYv3W4QmlF2QsSLW1Ew0I/TYw3FYeQfOIna4s/mmzyPZUW
IQblMCrPs9Ov0OYsEmIvqjhnLuISD0Om5KHxpMR1ynlVk+BVgGctArNw3h19uUhHbknCVkDKVb63
89yZVXo5DuTEvQZo/jsypVJ37Zb66QTAVS4mQICeQEcQRD8Dl7A5UP5T1pwejJ1EI6fWkhwUi4vp
fxy0gVICdPPiEkAWyliLsdimmqaXBsS7WtEApaHhObYtjFuFYiEwkOxHIemTkN6/iYPIEQW5ENEb
WFutTLvkNw53khJGO74KgAvEjyIWXJDQkSrRyB4cj+9AMkP79uQLqZ94UvrtSLV2JBZT1v4GiwXH
MWs1FHn07zbK92sDPRPeXuwEr6/UxliPDJamulur2GQF+17duTSVwA40YODh72+VswkwB8CA5+dO
AfmDZSFScKr0O5rB8KrAh1hC2c82+McquhYWSmNJAtkh0SJ+CsIjJ+jx9Sku3WYp2dAgZxOFFCoh
+mUBGizUe3BB7AF2kKG/hl8IMEUxX35Eb36xbn03+85YMYq/e5XwaTFYd0iKFkrQDdoe1+fgQPmn
3tO17ckztqvYNaYqKT4U0gBgndT0ugVEfxUZ3mtKocWUhII94a9YnGFr0XFFIPhoLvd8OHi8hiV2
8Y5M6uxIONRB2hM78Cd6NcZzqq74cGmeCdGdcwfXMK1v61JSoSRYAa1OfJjQsHcTMrn+AbaztvwI
DMWhPG/ui4uiq/m3Obfr1NrtQE2V/CbLLWZdwgEXduM+K76RiZSuq5GOrC4JM7TTaT0PZJo4C6Cd
6YDQ74xGH6aR34euCkZHtrclOQqmHMF+94J8CTSK6yyY0FnlURsghLAdBvd4/UzDuVyxhcOUF5A/
bK99SxWycUrnbwpYvj450nTdo8kIm427JilomkvhjvPOrpTO89wKRdos1d9oWE3G3sqvqAz5r8af
orId/IJfqi44LQtqZ8c5raqP9kVick37nThXGi4lN3Qi59TxH2yCwcPG/XJSoNO1vhgu4hLr+CuM
2yfwMElIwFVYCUQMaoD78J9D83de6NsV37fbVRncLNC1NHf/LIqVMlOfSFlqYswmyOwnJuiCuZKe
jwr0qNBauzIelnp3kRLq0TVB3YJbcqRR0FeN+f8Ca6M12Oqh5Ag5sAX4DHmPtoh7lQfB+q7Pn29j
QE4udgxWE7SgniWKBUH08p2C32nfaRe97RM1RqTa23mS8uvMdFb6mt/Jo5yV0c/qJw3NuyLEB2On
W2TEuRl2OVbv4KlYdyjR7p12g6sYO5u3FCtWsango9KtC/m+cYy2FhnCvpUX1PqTxENHE8clSIPp
nMJHLfoeiiN3vZGVeoPSeahimuH2K2DUIBmQpE7uQqQK41AfegCJnk/FZf1nSuUkYnkC8J6obSTf
MAu8B3MjvWheQgXINa1amTupRByoxBoDkBxLm6yc8RobvTLyoBDG17JOhLM4cFf+hq7e+g65aOFL
WorA2veQT8ICVn7aT43oh6kPyYYTpQFRWDJN08cix7M7JFaEJ3C817xRbwGrJaKa0jy9yXA9Njgu
nDJTlvBXLu1pIA1vMd/OZs5GOwFlsd9XZXDbdFrMplHgoORlMfgplAZdZd9uURDy4dsbrvfDCfdS
EYSBVPwEnE6O9YYGGPiBilB8TdJz56mv0/94fN2nVDiyZKxpBcYVbTqvnBdow4OEuuRf9C8rJNiV
UClPZK+g/iEHSNs4nULfIy22vuXdaHop9zuXF3ByIzwabPbtj8mRtTWhgSihyEChMCCTECaDCZRq
0zOPS1MTJW1YM9mniXsMuo5Xuo128zuVLKz6g+dlytQVNo2UJMtgr8eXt3QkpXlzEki4ZiZR2ZLq
VbOBHFBBoZjZx3FSm3dSGfz8HWEbxc4MAdrd0jREHoBd79zOIcTZmmcfZIpcTUecZiNVEg4dT4S9
iMQI0hQigi0rP9Q8rWqZ8BJRaX7IozUbTXxD8pPlmRKX99/SYfcMcSnQz3g0sCz6otxDNd6Gegx7
+B5mqPsNeOE3awWMdPmKED/OhCWQ+G55CPwAsf5Oh3hsNZv2Pz6wZxgPcZqCWJeOvCguSrCDKjpE
E3wFxPwyRajwQSjdPKDgI/IS0BDzhJrRoGfHUg5v65WAAF8YDi1eLOYIfxvjxhNeVG2uxCyBeqkf
nwQdtQbyurWeIN12+pAfk9gkzWiVLYrqg8/q0/d6LkLJQ7n50gTu5elqO1w2FCysyvZTwRfzeJ8K
7dDWKYxk06/oOrUjkqq2Ye651jT7re5NSfJX+8NQ/fufR/svlDaC5Jeyt3+6zl7NS85OG0/+HBvV
2BxwnGhBpXvxkGOcEhTdm17pq53TRPG1fU4kAPXtPaF0IWjmylIEHGt33SrlWQlkrnNxhUBy10aQ
yc5kpoqOoIqZ3jQn9jxwBHPYcK0To8Zu/yRkZZZowmufKdS3W8BwTs30Xd9fwO1VvhmI2y9EVwtw
i8GrGfOHCc+VY9wwGw3LqmUurnY60HPcIUJF3P9JDO0iC2IgIqvuQ05+Gk3brpacP51QO+2TjSqm
gMqdLXCtp2DiYJVlijYQDOjmxB8CRo4B64gneJJvIVKoYgsMY3wEsECeVCnK52e/YKOWv1FJB1OM
a1Vm1S8FegI928xwBuyu2+FGRSm0caduCVS9Uao3u5x3YtGbs29Gsuq3p/2AwNT/5dQ3OoudaV9k
UP3htzgCaRPRnNx4562xBQDFGqoXbI2Mk+CQSOgSbDnsqRIoYty4I9VTXNOaceZgUGuZWKjBiXg+
XjrGjjAch4I/xCQXHuCC0noAHOEm8tr1JDxyabUViLHRuUwkzuAUla+GSYASw0XOatPwIcZV8R8q
/qGFO3tm1dOuI9+dmMAmffbcuMuHDl2BOAz6iK2TJW5cNbhQZzp2gLs1tdh/PG7G0rzVwGdXPmqI
J09ZANJW0CCrCtsOjQ8Q8wi3n2tqgU9pdT5vQIBKHqeWKhj/cyP4+k3ddzUDV9/+WZJHQlCYtjOO
iBG9iEGbLBelsva7g1OuGacrpZc6J5/wxWEQEyH1mzB+e3eOtLaR+OUzsM/C8A52Ibq2HQ4wQ9HY
x/6vMO1Vf/72fxfzu9RCCOoEJQDrD6V6RUkzvEh4jZhFKkYWPWLmehMFPybBMjGY8PZ5U+7Vs4HV
xCCt3t+xIcxTDI6FwMxGlsYvW0pzkxliVvrHux592hTpK4mG+upoVdN/AAz6QF2ETp3JAuIWwglu
JujJt2ew2JLTYAtUzNnIH+w/mDgi8p+V8udkVW3CcEI7UBlIo3fVGoblwD2F+q2CrEmzglyiX4Uz
g7tCAreG/DX5Sws7cba/0M0gOU1QN05RMTplKdVu7PG82SFNELcsJLxasF5c+bdji+OJbIjR+CSH
u4LnCkZq9oaPJXKtXAe661XcBCB3MGfdmma7rUEqrHBEmQWi2AGXWRymqikGlGodjiN3LN8x2scM
SOL7O912KMkWa4xK8u7e/Lulc2VB1aGFJftN1/2DDMOKlHxUEgq6EzZSXE+6eI4tmv0nqqKYKguR
xk2B/Xe5jRE+BBIZyPSiOKXGnli/YNATIkHNauZobArw6mrznAW6aa3eHGZKdLt6JJWSWh/HMIHo
e9qnsqQvwEtk3MKGN3vcNykHtPrUWyw/A/VRwA2aNbz3ZGo1eKEaG6YZ34o4kwunJ89/spU+nB+G
8kEnG+7Yj0lBcKFVWzHkqwdmhrnrDIOGsAOQRbNIBI60cgySO5jSZQP/ott6ykoQzdJ5secuTo9m
6+aT02tFMXuvK4sbSjfl9MLM7twya//gyRscTZ7KJOiqr+ya1xxzFio9X4030uSby+2op8EO/zsO
pmDbd2/PPduhkE9E/jfkQupUCRQq0Gl9dUNIoq9Iogm8hXbI62BAmOzYN9muy1DeabMW3rSteiut
+aTHT7kg5httnmAu+O8T5/xtC4wscgPcbEjJDUpEZaAKSRwFSMuEzx4pHDHA32MfFGT7IX/l9tDe
1lMxm6EZpbzTElovbg39tc5ypBGPrIrP/tw1I3Gdcwzo14ysiZ6ySxfp3su9EYUlJAwWu5o5LJMm
q2JWekuP4nhMqWczF8fR8V4hjgTeskG/uYX780Og10D5s/CpjBwqDKA3XphZf8QujGCCXyZMgEJs
4WAzSyWIvNYbsje8p4hH5Ue0xBVcNQfyOlW4OrcDKRb3Nf52pamrOGBhIqFAs3IjWJvlOnEJts52
u/4jLdys/MWIueqrusQjTToCpUybdsZiClo+MU9EuXbyXaxVCUl8rPGCAT+CKUSkoXAtIXvOKl0L
b2xWq52oyzzWNur4g3PoFlujnrgRFU+GmzXgjTInIquDHqco/C/GP29FaBOPK/VfT6Tnp7NJFbUA
YvuScllaV9W4BgRyDnbI1lP3IPNQAD/aH5yYwBGjn722S5TgpNiZXhvK/esD3XxWdQkkOUXIX7av
MOeTkM9SGdA7WOZXUcVbO0mh39m50M0MqzMHv1bdvCGpZRIkBsRIDDpNWTxkbeZooJeStZfWJFCm
2yHECSQetdJZjoyviGt9w2tVwNn1zmEG7eaAZAy5rW3aXSwl5vLkqLSHACA1EvPCSeMw0ooHJ7Gl
TAENJ3IcvAOjOP1HUeor1XB0QK8T1fhG2/aVM8HKX+ob2hBGj2aVxpEtfrLJDgrp9yFVC/LoRzsJ
ZTxglXLj1C3ioWZoirNaEcbqJG5zdpLUb+Oz3bwyFx6rJfk1LrP+HWjNi4UuFdIkKz96JHi0vxyP
t7PUG2Z3pUmfUYF61R/YGCY2XFZ0mFLUP+xl1NuN3y+9hyGWe2nN3vqHFNpp5f/h4XrDNulz4fXu
CyVXgIoBywHlYTpKB6q87v1DW51jnGz2tNbeLxhKrh3tChBIxGB+jqTsftBE2Ol09/2Xx8f9YI6D
TZgAoDe4P/cBbIqPLH2W6OeWU6/kufQczp6ak0T6GFb5cUfOBM4pIKBSV3P4pndgOb4VAajBHLwV
Gnwve7ZlitfmwxR4ilcq2xlHjDc5aQCtlId767wjlUCdSqksffn0Ou8TcnkAymmiRKIMoZlOeY1w
PIagqlbdoSvzbOa4BA1XmOKWasKrwG8i8608YA3rchIgMmJX93ql7AxSMrCKeZPizEbyoBbYtW3Z
psuLTvAJ7IDbGu1mPoes4uqoYazQpeREHuD1ib4MtvJqM/ekJ87hFpiv3tn3ws+gYRbFzwLNQxah
y3jS2tV8B7iIMPVLGBvVnun5dnqed6VJLIOJQH9O1w6yaY6IVjDY2jHGrG1q0ecUFTO/93XC257/
PESZEdBjOd9PhAeoiCS8Y2ZnijTeSNv1l6Fy+1v1aXnZvI0qdeH1ahvHzxkrynEWIWhEFG3s4hdJ
o/FLhWdytCwLlZDNVl6+7x95bKFlVOJxABMp4pivSe7zziithks3Cm4WaSQ+YEb+4PVkRhJxdx33
dIpp1o8t5qNJN5X5FbSnSRgThM/SXE9qFpTaajwSMRWW/4KN7UkRPwBvxe8uJbRKkNwgUeIshcD+
0QSU5ZtCZ/o1mYVwgRDmhxfWIWDagA1oSMbTxbtdrLWK9pKLJmuMBB5gpjb656ciTZbjVfUE0ZFx
pVaxCPubooi+uk2jcBbVUnRLehriEbgbUTsXs7FyxQHz+c2H8sbT4hRe38jPTgTTeVr5jF6geNXR
mxD6iu9HFaPWrE1cXcK/VRkT/JIdyWLKjghVO0+d8dNC2MQ75URdQNc1+JCDsbOISJgoJRjnjz3v
UDYwc6EYSFmhS2Tu00ow3E25asFteyiMaIn/wqnPikhiICZft49U8t+d9KpsB4rRU16nkb3ykb+G
SySENe7RcEO4FIPSz9nm04YOPEnRHPOA4fW+k0O4X0tOEMkV8a3hsg5tSg46z/5RNziyg2iUizI1
HU0StTZZ7+9JhQ5s+LYQs1fSkflfyHpR2enzF3S7vO0sMneSM0HiiouiRtK2R8T1W6jYMw+caZh5
64OvNSh3DVOso+opiLBAYii6NPxg5syyMeNIZ2EJUx2XFKavc6pVVA0tgEHuRStez8/SMDWo+BOo
sdtY8TiLXWdb2x4kMl40rDDkK3I2N+GVVzciLb9F1osh+pLiI9mtM05So193YWLKDOCZSTPrX67X
U8C72Od0Xe12t6XjKVMZFfGG/G3ajfJxZcnX/5UckUfJ5RzfBCyWa17TR+rGedBeVyWUE4E+eSHv
kkYaafREFF5B83AoxWx0mMZ/wT0H/Zmk+qxUGlMTbEye6aJ/tr7lQmh07oLZHEmUHsIlhq5Gmxgx
2GWRbDHMordm9uixfazTv4ciJ84Vum2zsm1uZCBCjBo9VVTcysDBmDqM3sH4wzqsNczCZZ1q/4kt
NFS9Bplddl20ISlW05ITS5AZvCTvvZ0XmbqqcbfO8/6ybhtAsPcNkGntjC7xEq7ptxym0ZaMja0S
e7NxNG0T3P2vZviNmjTuenHO/rF61yBZh2o/9l1Ch/I4HNnVRsQ1KT078n+MzLw/f72KgOFWb8J6
cAZYG3BI8B4dq9APqVpmyEKekikPIHpppZlBYvVm714IXiep7B2okpudiptXHXaFmNA+fJ4sLAXz
4yOIbo4VNhckR1gIwLkF7FTwSCJkA8apDLMtU+G7ZH79mCGUU+ImD9XXjW/U+wVQZDbZgLCnBCTb
X1TW9rzhTaY41eHeESEqlGrMWWE7UCL6DFBaJSFIYWvQ/KcQetjdYw/9AOrlL5wMpuT7LXVyEtOz
Ws6vr6HFODwgefUpf6plEGik586+wwoECNL5ebImnHrMuBgohgBC16++J4NIzuldk89zOq+23nJe
Kpgh5wgwjreU9uZA2oiBiwWvk+BpTZfj4+PXH86DB7hmVtkxL1eXyxUmyhvI96r7pbb1ftAepdMU
IZqlB5hxsRHBpRYdDh2LEBZ0UuRRJ+qhqSEfu0U/vMdCjBYU1lXNps29EIdRP/IQcM8j54FCSZvH
FTvVcKtka/JcL6LG6usqnpyIWn9P/nO8E7cfO/lWrbHGDm9ltq6g3G0Af0Lb1sra4xvVoZxcrG5E
ee6SOEsMceavR7HAMT/GLr14jk1n4n6bu9uO8Mq29wbRAMpvhFZ6sbmVHkujcsd2NBd8SyyfgxO/
AhyqXhIAGqTv3XfGDSkAbp6/WlfB10bCdn+G8U7nL/82yJ8pDcFtVthe4N39xdPS0YpSX5uv7wB2
9jDVoahM6VffaUaG2ZN3B1JZc+yvhRUHZDckNAIIEV3QXd+fYy+PGDGjv3BK8W2Uk50Iv5Td/jSs
ABqqjOjjTquFxJTiqIFQt7P29dQrhwPsSd71LzeKiObisC08wOvR5jD+TTw+T+XJwAV72g1zO4jy
VKnbfegL0tnF97rnKf8xOo2gUkvh4Y4yvd4RglN4k22n7GeALZsyGqeeF4qlIRjrBZGSrucQLWjV
5DztfIqIWBYt7jHuJpkDvjhWGF/dOvZ2kz8cBTPidkgc7R6JBJiSKGAmyswreBZ/ISfrYlNk8y7M
YtjzJFNB4stONHGpD4kQeeCkMkBI3temeA1tAdelwzzfy4GQXeYpvV5Ht2qbFHSfY2rcyAvXy9fq
8LecYmFfYtX3y6yMabWEXFcuBojHDhDJu2kuz+BVPGSAbgMMp5da3P+H0zN/mILj284biYWeo8L2
Ni0gUxrOUFY76vyuaxQOSbw6RMD7iZMazgANWaJa84hwzQgSdrpJktRYCLuCm5M8Yjd+XvJRcWnM
oopi4o86CFSIER+v/XUYf8RiOPCT+cMcIjRwyVyfgixeUdjYsAhpfk/YqU84aRk//RQzOFkYrc+3
2yTMG3YrfFa7UyCkQ+fVuwvXfdaGiVy6AQ0of/PTfMaVIDQ2jKmeWTsqFdqPzys8tff09gQH2+AY
/u7rXH3OJJwOZrrsfW39D39fy+ueSWSbtHrbX2EJNAflw9e3Whd1W3L7F5WyWliagmvjgC4dv8RY
EW1ue3kIMJOUBZxa3uKuANwkgv3ltHDdbT0sx06WDCDNrBpa6S+/QQRY4nGthQ6KgBFAa7cKnklF
Mq52FBA6m64g4b0QINOPyema5WLbZmV480XWZLZv6C9/ql8faEtYuJC85lUo9ZZotE9YnUqnS6RG
Xije0YDl5orP5mqagtZpeJL3eFTKnFid9hU1o7k9N9Z67F5DIhSs08mUYbLWfYKFlIK8bIKFn+E9
9mObigKj3RKfeYdHu7f0Za9CqlJcqjAqJB4W3ehP0KfnwT5vTCAa7TPj7kuYfNPQNs3Y1Zg6Ho4l
VCHKwKZq4GQPxMYw4WVKm5BoXzzomzI7CeFHwUYvxNagajtn3gS/tFp8fABhbZdHZPMKzNlKNN9W
DkPUy7UcYgnaQzG0dMUDJD9ujaSihjqyNqHRG2pON9Ef2YWKjj8MH3FPza7r5akQej4UbYEEEUvB
yRmVtHYPAJlgUWzhi/mKzEyc9N7FNG+BhgG1N8etf/I82TGfku500KIBGxck73zwyIjg5YXvQeHC
bIphsNmq9jS4BgR1RJ8JDjyDgbq6/ti9Soy4gSHdBGDlsMbxokc9ue6JKvJ7MAoullOGtpG/4C01
FqTRpffs8TU3wcvkKxFK7e8JzHFFWA9cikgkCTZLOv8dAV/EoObmnvmlHA8I6GkzABOFlSI3wxG5
zi+5jy5LPnweU3EWc8jYYesf+9Y0CUKzQqdIN01yzR/o3ilWP9EPyvyvrXnT//JXhjftFX9wmZMU
yl0syjoFbudSsUfWwJYxpcHcv4k4S+usTvDjDP6poMzRoA7r2Od+HkFoI5RYf4D+FV3MCunb5E2R
WQuvS8FaaedmOlCXnBu4DYSsIFxBubIz1s+QgBdaYiCp0CRydYVPchG+pqQrv3bj5yPe/UwfaGgW
Y8BQdoQCRPWr3bSuMp7l5hAoBL/yhk7P5c3DlDDHZi1GezJS9xrGhDA9g9wBTJZn9io4KdtVlMDh
CkK7YIalBQmgosklbyusSP0hHhewoGh12OKs03Wk+TQccOnVdlNvKsgTmlOF8r3ZGbRCni25RuvB
dv1sY/e7Eh7tUBYMQIL1EZEAAtaPhE0vy5I4024rk6+NB7xN5pnr39TvPlQ8aUx1s1tHvEbFIWh4
Kq+4CcDpPn0yfwpxYSANL0AoVKbSjy6uF5UGwPAACWc+eudYlsf4cJySMa65HRHl7Btu4WEXpq94
3SfrRELPsmeHKy9xQn4G/32i7cKbF8IK5Xy5dqtjMAo3y/sZ/Il9gNf7hvsR0TXD7eQP0/9A3bJF
PKqR/BylxOp+l1RRjsSFvfaiE3z5YvrxpjYlWth628C+N0xdH6Ww/QY9iH9pk0cRvBwVs+ENCyyw
f/9PxZREQJgNtBwKTWiyUeS1Eq1Q2M5qEgS/7wFFmkcShMSEiec++psDoW8FO4QkFbtps3dNfj/9
QX3Dz9xmq9J7/ilpp9bxbCkp6KNwB2pfEiTeFn+hdr6gp/FyLYniQW0hQI16reS5SUFum7AduHsb
z9ulVHMkguW3UP+IIwd9QBIi8BTGHBtH2ub524306brOIOl7LL3mqRG+8FO6fqqUTkRBr0VlFjyn
RUYfv1yQkFkZzU/TUbe8435TMpyl9+LZtgNoxEmdlspj7FzvLFoYlG0uM7DcivXrL8Bo9EBMo3bf
ZqmD4m38TJyc8tr//Qf1YKzCfKA/TYcKEUeFKacMTI6WQdw97t3x0ZYhTceHWR3JlKSJ2Ncw0Sk9
10nme8x0Yxf4PMcn8Tp9AOTITlZKxI38C4faf6Q6WA3L1R44KwM0XZcCUasJqYPB92d3e3CVQHT3
x8n8mFsoyTU75rWiqd4e5+qNxA4FliHoSFe9rJ1fmrofFCafKQ3CWwkwPmId8v1zp3CYQexrbKxY
AfxgsS8YOCnW58t4/3o2JrmXaZjHHjpfZ4Ti+w/UNM615iVJCOFoLcu4f7IiCpSjy3Yx8CH6EGXW
RiSy1meQ4ViWBNqXjbAcm0Bpz73JqijbVkQKk2AoKRZSPqTJVtM4Ac17cQgxWG9KXwl6Nun4H/oN
i4Mrk5QsNr30mokudteMcNWTeaFGhry1UarnneAKXY0VNaPbD9jD++9ycduuKwSHRjqBw7xnZsDZ
JonxD0UDX3Fih8bsTe19ixGTrEeYXNQjnn4vI4QuFF0z+MkJmoRku+/7+RCBAwrTz2idV+UhM2ue
6bD8VSQnmujUw21r4JKmxnUorbBqlieBlSY6Lh+OU7fZaal8PH9yO5hDs+CjonpX7uBZ0cb1DOrA
LCC2BEZd/kC0WxqHkY195/qpsEZK1uGBIq2CfSpxvtWTqCLD8dV37kAbkUU3lNyaDQZN7HbHciip
+x2ln+m48h2E8YQy0o/WfAsdF+9kK4omDViEtLisc0fu8AaVHpYoH3UsEgZM9pp2T+FBNQn8eu4q
Yj72P8/nkTnB7qUje4N90EiOHIN2NhnQSlJu4HCExJlDOn59hvZ2KnZJ/v2/uutv+HYeIL4FZXgR
8llFG91Tk+vONG52yQpz3pEI2sz7vrgs78Oc7Jkv6EzarFJcw8QPxldIvlDlETM5BWP4wxmYDfUN
j2Z7IxzoT9HK5EPVbFJuHq1VKaUFNjsOSKJB5fGQpUVO4bZC5iRu8lFbWBoIvl+x17fPAp04sqZS
nzWgdtMCrxg+dcIvYDi/Hu57PLsqWOBgw4WXEZPG4o+D3xDovj0ZuIueB9J1Kzcxo+ZiFvkFL9nP
sOSWGID0yJDJrG3StXKY5r3QsXpNhiZZGQx17328fWOar3fhgV4Dzjx2wSYLhIJV9Ab+faM4tygp
+jdjGluACZGxveZiUA1SvXuFqHvGlL3SDe4+oAajC4kot60UryYDhJVabOuqsq6WrtioWWVyc+ln
TUJ1mA0JTt01PDtouRGThqThtEybwp2PpnVyjitkZG1CEcZVQvtnBch0lxFh92U7sjFAw8IUOtYI
VqDUnKoSdLF0Br5cAP11G067qN42Uwqp0pIDk7CEtqLbRl9DHJhjoCptzSLO3KGq2DJBmI7zwZbS
hIx0pgIyipxXmSHzvi1avj7j27uBuJDFBvYilRunryJHoL+WzVpSz2hx5jkbBjlSc2Fp65R5TX0q
rPkeaaj8Z6mrylpoU7cHi1mItUyxnAoLFEyWa/egao8GzUjdmX/4Hf+S226U3e2qWqSKhIRzjSsp
Wz2KxlTaWCUZPIsErjKmL2r+3woprGrkEEq3eftBm55H9hLji9keNEhO+PEB4OvGk5x1kHa9Fwby
yZIXjyNj3KZrKaWCmB9nrYdy/sma252rrtIkdESEWOWAj0cCzQ8wiP/Le7lTT4LTjjAsDQzoRvQQ
Ov+JTWM9ogxLNd58hoyANIw1uN4fa6YmsAD7+SNGIpx2A/jPaSilgwlSMTYfbEPkGDB9oNy8kVz6
iALr5T5XTw+hKK+TcJmCoJKQf5NGvM+qYkB4JlgadkzgodGi0jTIkLw/mn4a3r96d1oXvQQyQxlN
TLRYMw97ppUF8UJek+B0AgyOj4YZLNnViMenwAzwk6D6CYXh8Kbl36caukhg52StvBd4pjMpaYgb
8Dw1uiDAzuoBOJAiO5zOrW8345KpaYGU5EmQ6qhNW8/6/aEZeaGCwKPWK2iQ3ABv72iG5ilRkFm0
YZ3xb0+FcxHkBB2j7s+y4w7HFbSv77dx9XufKzDtloQd7ud+uAY71/aNlEGnX4t+uhBNq9Dr3QZR
OuR7isRabk3N3UPpgoiPEa0XuzL0TYg1xWHOktgbQPULInOmq1cI1tt1Td5WqBCwQiw5G0hdFF0c
E/HRQR/gX5N24+rIo/lNWpBMQEhtK9H1reAP3OSbhAlF5TOLL4CfW6S49GcnhkzYO5foU26cKEvt
kK5v40Uj3Uww9rz6urd2OX5Yxugs2ScBifpOp6tavWP0mzCWkupp/CimHesy4168gqakul7XICTa
XoWwFOQkDej6ckG9pNWSKLAdvtQ3j3G5+R4HNFnY5VRgPer3DB79hx6pkFVn0WkIIwLtKI7rcN10
318p+OW5LlIOAvhbCphzui1Je31OdTBfPuVEj04rOCGo+JRr+htzYXqNhe7Tadhrt82Z5kw+l1C1
cY5RPPMYis3F9nsUa/ygkmWKRWb7vTnAvHAhRbA3G32Bq7nrD7VpMy6woU+Plod5I5haCR7Ra7q5
euM/6304FT0Mg++Ku75E4hzKSP4Jj5qo0RxvgVhgNMqCUmHkkzy0pnwUkEne2N0qrVWKxr4zt6Xv
nG1qW5ZumWqzh6hrxqyA+QlepnOghfiafndOy9/B9e/gESrmdjdrSKDyvmfHHbft0Hh9PMeDJG8d
hYCvZevx4QTAK84PJ32P8uClxOBBlZ4lKWlKfxSkQDxAne6Q/aWj8jKSYyfU1WBH+lu3jwVmWyJQ
xzFc9rpFA9qvvPQvYSEFRK50XXxNVr+n0uk/0beWNJhwy1u9ieNI7qKQ0ZK0T0R0jZiMSUlc3uWp
7/doobmpaGQ7Ffv9zmU7xq9ZAPFwBoaouBKBjYDi6ZLVmEibhLIMgqUoZ/6f16GD82Sm2CRSFWJM
CUcypjyNWA14T7wyG+dNtD6+Wzn0EJ81FHK87OvVdHTL+lO27d7QnABKIREBXAAmEHXtyHQXUC/3
JYKDFITeZxXMLMF/SvNoAYuMncfJxcE0Hm/J5VUKvhCBY3pWvSv4X+KvRi8ZYahvU4XQ66kpiz/L
00YXOKV+TdDWzw9828aiisea801ZtD2Mg1osMdHgNfju74jsfR1SZRjOtcX+ehXSuN4mIYgqTPMX
bjpOsKdTku9ibl08tJRFJKUKKfx7sPBCojd6qUuSqNmAUTAYyr/4IGm1+jKzJkDza8NUExj7Y0jz
uCBwZJ99RQ5jlcKiRLQgTlbyr7+wSP2gZq2d6woIk1RaKJUCYPg5xsBc+Vijq6BHmrJfWxeeGRHB
S2hrxDwTQiincJsTjCFU+/mbhCdLfocQj4SkBn0iXxRK/h6jK52ZJPW+01TFGBI3AsyUPqB7T4NE
pOh0IdBUWJkX+Wfrdp16u9+QNvixys6tyZoP5DFYPeR6lcLRvtl2pQ36Ubn68jzALpXRFyclE0C0
Pd/KfrPZs7dUk5+HRdyALRLLcsxuuJ1JcXPqWrwBd6GtLWpSMheNe0LnupFrNiwzEczg5LeLlubY
h7VTzDwbikYBC2r0vK1agYrpRCkJE2IPNFY5sBuE3ahAnNAvhccZ0kxYlmgAMXed4+9VBEhSnlLq
dN8mpwQLfKZ5Ol1zr0+jXofoyzqMBij3l5/+mpNrCG6TdvXRJgd/KpSNzo0Dl3U1rcYRozy2Vr/l
j+qo+KSx1BnvAht/RHX1aaTLTMTyDQzqhcoZLHD74Rf9yTHPtXAPoRLcy6W01BnyGnd9KNj+6AOg
BMvp7zPzA571MAiFVGOkBxq1uyp4MjPQv25bC17WdGl7Q+EuxZypJYsTSVyE6CwNKnTJjLOZ0cEu
iiJbk/OA2Vc7TfRWpyzkOMxz7oj4zqmrQi79J9360RS01HVM20KzWRUBMg8YezQ5GKf6AADTJjr5
TuqVLq9uJ2kLy2QxWJIH8EpYO++TkPyBx3rGbXU0VRhRKeJ+ZU5ad7ywvASXo1edELvXF7Utgtcj
+v0m6G6aeQtNw5o/LxpbIBNGpS1GWcuvrVKpU6B9Bt6LZmY+rUCu4MjcemUaduh/6AiA63M+Wbt8
G0RcGFi8mxsaJQCh98/lOAj6JNfpVxEXXKuGiYzjG/qo+0StVjz9DzTy8rAVAVLeuDoxwtOnfnxE
Wzrc4SIqftKtWYgyEntWSWj8xOOmYbdJZrnpfsufbCQPcS25bX9SYwDXHWNUujKiJRwURdOb4SBq
9mTIivgdM/q6wJpB8H4WkJopdHjTw2lgX2t1BwzSQTy15N6w8fDOUNJi+alHdPyOlRABy84Z92x+
yd4P1u9F/GpBIWnwWsnGC13y9HKNrilk+EqxuB9t/VJUpD6BuDuNTIlx3t5RI5Ao2Za+tAZOPrZq
C8aOFY1wWIT9RPyHvHMf7F7XaV4tDodSMs611VzKs5GnMhWbEbdU+lBO3H2r+cpAIItgN65OzNRR
V0Om8Qx8VtcIaT2X1oQ6gWkxqGtheC1HnwGkQrGfKdm04inpXjWhB/10eMB6+a1lQkuozD3o+mcK
gTSIIzXe8r6ma2BIScC9pXIIGQMfyWWyNFJoWyg+VEnaC1UAdYov7u8X3LezvDzbM0Cjyx3uYcLd
w0aO2og6ncmHzVCgmQW4uMXKHTE0XscE1q6fFNmdPPLa+Q+HcKyb4DgZxMcX2NWTsTBQHbNrJgO7
l4PaWH+eN9+jPJ2Ly7LxO72ZRfb5YhDZ+FUtYdkJpYoBfeVCu1eCiPQADxM5XdNmpiqVP1C2cuNN
38eS1qJAc0VUb3KTmYc2A2eAPpcmcdpEVfEJxsHU8G9vdPwUnMZL7oRtyoAfMn99wVDm7xom9UV6
7mS7mXvWDg9mNhgX/U4FcyESoLTwTBoa62+0y8qjtTM/YKc9xJzG7bt8RIrvo6Wf/h8A6l6FTzza
Liw+T7dXDqVic3ldkQl8wn+2RdlyTMQW1muNM1CUx/lnL11FMtzwZCs+km4aFZRo2DBgtyuexKE2
u442W2b/GMB5BDQwv/GVssAk6aR/6+u1xYqppLvJMQUca/c9RYtP4Kt84HmF/xaHdNGXQjHJq2mL
mUKI6kRj8qfwRGUkGzmhmsKYAfqkHkOJQUNB8NSjx7nLWA3/wZOsrXTarHqKDLNsB6z7EatJfGZg
Tu7lmfTuiax1Qg53OIZN01hdGo6Fbnxkg3sO9UG2W9d8N1MIc3FWNftZVDihB8Sono/K2tugpM8f
ZgdkVkJpmfP6gpZYbvBfkh9FAco+8i4d63QZUF2ugia2kq/SF7fI/ju9ftEYiA9PPlFfZJqIHcqo
7S0mB79OsmNPur+wecbsvSVU61nyvSfEZFIB92UeBCtepLwnONw9p9Y3Mh1gyiFi/5IMn04vHCLB
nAXZYueYA+NJz2dkzqsuZkp13JG7LC3cfxwqPEn8Rb67D7gOByXa5Lch/FgPvMqcg14C3V4aU+5L
/RDhD+2+PLpHQCQQAAnCf+BsYTMSNe9aUXc7hmAp3R2uYO+TjwSAeDf1X1x2uoLEsyyDQUW+oYpo
mLrOtKHQ4tTIO9qZY5ZaurVJrk/GhBtWmecM62IcGnBMIsMM95FJLjX1hazbc5H9LBAPVbb7OjGq
MJeKpVMNujr7y9MyKXrhIWPhKaMQcuwgMyi99r3UkbEF2TFPSvGRnnO+jCnuyQXRTKaPC/sjp2Ze
z2VSeVBRMd0szdD44B1azh3QWcwTmXdsxka45JgTU+LwdNVqOkJN5liNz7CZhOVBtuefmL5IAXwo
2h1PjXxrF5XLwdd9Aih/zgiOZ0DcGDO3ZXZgqqZgPkeEht8ISfpI2hGvCvvSBZ5pYE6GfPsFMaNu
mYiwPbd04Asc0BMwUsiGblv/g77ekwEPP2CDW57yRjT57AIcwzHHc5B6/58WxQstCEVi/WXmaqy8
iRE76pKaAwtBJIv4rPRjoC7hG0JY3LyerJxF6z2JuRGnnfhOzZJHT1heB7NCvy2n93n72MlnxwMn
kDe+iSn3AIUI6+IHunWqN3q+f6VeGrKqte49OSoikd23HnA8E76zNgI0xm8yXaGfBfWcCzT5DMgY
Is11Bx60xC9lU+HKZOolvdwgOcNoZWuLJTeLGoPiMX26+9GygsAI6WRBZQBFqAjfZUfCplxJqLXb
vbbEl8kLlvTV4k1h1voNZZj6UlLal1QnZshgv7GazWTE8+yfQpqqzG7yhyvxw15rMJp39k2OBzPX
BZvUtM9TwwAevDDU5ATdiaH+fUMbi7YB18Wz2cecFAsIvKr/ro7WlWjARItA3oGmwMjn6IzkD1Ks
/BHV8VZ9Z3XQivjQhkp5lnybp9508Qhff33mogznSJvtq1AVSeL9cipuNt2e+bqs7M3bzk4FeExg
Dx/RMsyah4hIWHAvEnssTvWaRJgsXHfXZH2OEeEqrDz92YoxacJPDrBHk8HnlejRVW7iUwPflfWX
kkntK/flS4Yh7/OlpbzSrEN9RuOdiUlhIgEpSGt1UG0Ev3vA6HLNfF5yLfs4NAzv/K8hFYtojJ6O
9KmnlZ/M2G6Brx93OgT8awD49xSgpf76Xa0PanFf+6IT9RbI8NbPBNI7+2yoTENyxK2mkxo00JLw
pQUGsjN/KbgEWOR0ArvyNJ2W3EDszn8v6jZEWTriLBCKxp1SY8LDkgD3iIWhTi082FmWkxQJ5Qfd
/7slDdhtHer0Df8WOamjN4tItZOUYmu1VWr3Xlz5aSQjr/MygxiwEN+CTLCrbih6T78z+j7ivfqC
fCASMp/sAlhsRYYW3hraBb9tI9QUSFqf7E0RerbSKTpK5x0P2E8InuVaB0COPjBnsaPCglP7HByg
IhN78ssH6hfaaL7TBrArVOsLcxZhh27ZCAmWB3s5ZSjmPjhNZwgz6nSzteOW/fyBp/iCvzdXhL6p
3EU27NLJ8iH2Ea67BMFc3UXqLkcxclqIb9maVv9T6e5fhbfFT5WOBBacam8xfsprOchtij8SOD9e
YF/BpVIMLLDoNpPpOdukcEVL2UJ4gECLMVlAPCBoSbnLjdhbHuKUonf8JzGPIE9fSQXiuxz5a84K
SEWKQsF0amo5M2vPqSnAIOQijhKFSZrz+6tmO5D6MftfkTKApdvjTTjowelvCLU1oNXDYUwQynJd
PN0O2Tt9lIv5h7KEhamh3A9tmlf+mVUDL/kxTSeZEPMFQQubM2WIPr0/P4xs/aJH9pm75q045QzQ
ZOEiDA74tVhKCo3cvCN+4d9Hrg0geOjT7Ym/3dh0O5l5KUKGGu0aCzMCejWrG8QhXeCa1vLmlY7o
5bFWpZFUdQK0t720vBO6O9d6JqrnlGOXt+3rVTTi4k/6ktCLnc0sgNKYaUqRSkUrmn3eTpOMgOx/
bKVzX6vw0zo9lXYeV/9vqRFdCyj48q2J305+WVCT60f4F8NbUCXTNUD5fzjPwnclMGL8ni3cG6lU
IYX8haYLOm2XaKGWf5bv1FmAbR4aN0zCgnmTTf89oBtXYRyl+V0xdDkjt3M7Q9H2dCRqAroXFP3E
90tJn7ZVMy+DNlAXQS0ENyuYNC4MXLiY5kZBuEno7m5hHz73NyoxtdL8Q99WKxMKisookDx6IIEc
tO000VFepcfyHaoQJT1r/DqeBhoesIHig93OfzHOxk+HJUyrf/VMIygC0CqDp/kXWLNxPTyFnWDo
n/amSvCaOQ0Fnur4V4VG1eX2ZfB883BKqIj9lKd2xLERc+v2WIbff6d4Hvz72PHGs9J4eQieQYk5
n4IuW8xTwaEUYdThWINc5sHjyykRP/1GbyvFGQ0gmwRr7DR8Pbzatn8oioK1X8FU+Axl5ng2osDK
0ftjD4lf81sSIvm+haKd1k7JfaYPSmA3TP+R+fMdUaQj6bFihUPYFHdVNxP8E6c0StSRWC2mMq0Y
veuQxRpeWNJadmCpruNa1Ghln8OLdfS6VD2jtDRKDMj7Kfori78FC3p/gQPjItt+PoLqX268lDQq
mWrEt7NAhMe4RJFxjWhjjsSTbA0ZA4dwDq5ywOesMBP5vxv9GBhJXp2NYK/Z7DqNMckrq4ui2oM/
qax79breJOcRVH0cT7+GCmqELYQbwrd/PiuDpmqqFCenhlfbF0t74v/jBZizCX7PCnAkkP0YNImY
zTLeJ/HLp0ykeYjAQ/DHhct4z8vgrQ3vVxwknFyYV2+wC60OFwcWbPZWVMz3qzwXbK3AQVUFPQov
BJEpd2G1CMnhH6axP4BdBC2b27Q+7ya9NJT2KVOAMdKygy2Rd2Ng67FJMo5qjOpssbKYmDpx/E+H
L5FfTvrgWIoNwQgDvQVU2WsAKNzQX1lf2/G6Eq5FAz8dIZhm043Lt2OUPhxtSBlOXEDJtY88zCoA
Z76UH2i7BEDj2/9611Gwllvr9UC9eAahYkI50yEmFPvhEF1qmpsLjzj/Jw0EtoYYWZkqBXunEzJ/
V8vA7kw6W6t6ycRVcWrPS9A7Wvo42J5+tmQnmWWsWC04PIrAbTGbj62a5bjk8mVnfouu1bwMe/Hb
PyfRBDDdUJYiBKE1r9IKXeeJ0T8n8uD9PO0XhGexMOWqyBip10kW7xT+MsRssycd+MaXQkHGfTJ2
mqkhCO0V1CM9zEljziiOzMYD0vXHg/rXRd5cjW3Xv1doAbsQE/7zEczg2pR+40XNZ514LIGVdbyZ
Zrlzn/9N2/GXMo27aPUQnz8/o3JFjssWhR+earmg+eRRP8KOmbGlC0AbW7Su3TDOeRgS+8BYaF13
bomuOypft1scsogLe6+DOhgOfU+DBlDDlZi3EKKMwmcVf+hPnSiG2JIn8DBEGWEdeP9M0VHOmu7H
vwfAIby+egtMZYoeiC/b8eaANQ//JRaEnY+aZ+Gx8qgC+Jikl8OvsXKFlzTODD6s1ZDMvwoLNROl
EHFoo+acPtGZTuQZLJdaecGD64Sdhrro+LTXuqic4D5Zf2fUkxCa11ru8Zce5nfkWuMm7LrN5kVe
orZKlZ5Y4HH2PBh5fByNLshbMPVtKnEgEoputf3Vm0lOAYo205rID3ovhAxOsqZImjTakVVe429s
Wo/Dm2q43uRRnmC+g9F4qxkEL7+pgryPxN79GLGVKA3zuO4UkJLI31Dw1s82hWN9VbNXw3zMmZiO
2cBhOYGRYSno7ayTstf2na39zI7HHHj1GuHhIbedED8AWDNQE6DMXel7ekxQEa7+lstq6rRrwkdc
X/B5Bzno03bYI50dD3iMdKU+Q+0rNcybqqBqbdRgCxQEEQ3FFfZhD09GQhbEZF0v3DXVsbrbjDPO
dr6VejckAW6C7ahjHiVD8o10mblH2zjc3rgieEarhiCjpsw5kWH8YoSZL9GdSdwUQjmDXA1eddnT
jKz2YFUPKxC3m7rv5Siwim/Vtf8lGf5h97ZaJADGtdWGDyRteBJW+cGAYRjaJSbtRejy+drpsjak
R7x9oW3acunRhCMPsBKHss036KgNvdXPDLH6Hm9UxmvoHopoOV3r58iQ8A/JfStyzbETny8REBp5
BsICKYfQSILQQ1Rl4WfFrFu+Qu1L0PFcaFeUu7+R5iongYenYx0gtQMJJa/xB2yVZjYJh47uaG9T
ht8FCe5cxmGAU70EFITWM8D7NOymAOFRbn3hlhBkdp6134BljRQl63gU4mLTHcWOs2uUgg9IYHQn
v/xqP5qqL/D0ypaqJTk8it1l6Ca7Upq26CwnzKBQRTkQKM85FieDXroMSnQIOYGzO7NtmV5gv+5L
Kn8qciwcImCLeWSSxs/CZEPW+4GV+sqf9xbw3NkM7Y1gCUc81K0tYBzzr4AMcs05sT9q0QlMaIBB
8YCF/eRL/nP0clAJms3dMrlJ3iw2sA6iKf5xON0Fz3vMbmMjeF/rEotgZj8w9kU3Pz8OOuJ92e6r
TFlVbUY4MAnz9SVKnjUSHw8udjKxPnymQbYsU3tiwd9auZ7tRCm2oLzUL969DowpWLld10kK4Yym
Dxuy+9aP1el5MtcID9zQCQwwVTrVmYlOPRcpduMb0uciKtUbEo/DXfLHVOAICEUSqW5HFjhZ1wrc
euJwb14QLgTtSkNrjKOvuXYtJcwstem3PXGRt9Qvk4Z+ZooP7Pp9JArslvc+zFCPcbKbCFhL+17W
6X+M3bJ1yt+ZGfeRvWTUYQZ0tJ/wdHK6QQxO0xYNpvcqiwSoIsXKday3vQfLEygvMRQ2695XTmqk
z3iCMg4hB+UOaDTGb8CETksEmS/+/Q2g66YqY7z+S5LWEUoFlKY6LhtbQwVEtIYMYfKVsFok7DAR
9w6hBp6V7dGr8hMPa+y/ia99hRo2vc9eAJ3N80gLtEDadBqTkJ7E9ddNmvLz+9CuIidXRfCyLX19
LIWlbp+O+bAtkDVnWtfWFhzniI+JmwwL2wTV63OAPtSy55gVDdOHOJUusoah/34tIv7W8aH2sK2v
u3rI237L5B+c4n2a/783O7Eeo/WWcrrGEPtglr/BWqkE/o+fxiZnBB355Q319/sm5vFBl/KaH/Sv
vh/E0nPY5msjaSVce7mkHYzK2p0VLq3ZNqk2VA9GzkpPDr7tEmE0v+ih3TNOTNfzeh3lrWZs7RMQ
LvgZAGWW/LhbxAhPuzovi66XMUUb5LX2e9zvHkzVIMrmJo2VaDM6zqdd7lUHnyRvL/yQZZiAmvlj
P4BoHFJff/12vilj4VPevY2ADwSXrBASGglQ2vuwj2vChnnyMsE3uTtBfzBzl5ZfPl61mXagb0E8
E5LXneJ2i+rINCzoz+NsfJzVjMqT4RvTzBwIzxLXwhYDjwwOa202UBTSkSGy79HKYfT03nM5/BOI
e4RuPaeQ71O6vYIy/4EiEgATLr6StL+mHKOKZh3iMwkfQ+YoKlKeam7rFX3sXrNRmrjwTeX3CgFk
5ntwcqo3lJfisQrq/NykqK1ZVfeRN1e0v9qigTPKxrD3X9KsmqPiVt5bxjZfh6AuKBwuyMgbDAjD
XC2lX6ROn7sITe17oplkaolhqbBpFw4Eu7CuFT4x4mC2vX2qZG7Hqccr5+dM//q9evVWAtuYIPPj
iQJfX4FHUQGxZz+ViHTaVDkab//n7n3xKWGNjaD+xyC3EZEGCUUGiiF+JsW0oWXXOStJkD88R8nf
SIgLKwOa9o9hL2WPxuiU9aRyTmcDLI48WAldcJPwiCua73RYMg430Nz1jAc/NRHgByOKFmE+PVwl
TmWZEDw1olQk8coEJpi9hmGtTR6RejgQ4swW+fHI5xo8ZvixV4C4XJEsL+35E5lJ85obBEsQfRMp
rw9d0CfspQhuOsD+dfskvtv4oJy9guA+RMc4A8SMauG9W3IIvJaqesbfvf19tJMh4Q3wptDb5htf
BQ7fSxrLw/yQvh/wPXOVGIEBjgkdZRy4bN6i8n9oQCEoA7Cb1j72rvh7oSblg5HggxxkgPpu7TQl
mk4JqSaI/ZHdldtjFosNZ+4B/7XsIgPuJI/zCbP3224MAr/F01MmOqVKjiff2jmVLdpg3QAxkuv3
997qseFzvydbj5S/4AmKAHrsNgMHSTjZ33/Or38QKKfHL9/U396C08akHxg4UNckh5OyVGUbEJSc
GD1jmpAX4MJnW8t18eN6uogYj/xwTeK/xrYfRcJ6gbPUtOetqzL67pEBJHqiYlsIk68uuKxhYmlG
6lpenPrLzteNj7Y+L3XQg7WU+MlnngZ1V3urHe340gZr+CpIoHviYS0IJru375dlR79CRqntqotJ
ZpwZhwRXDZdkzzlKHprIkRWQ1DZNU4UccjSohJKsex0HWhV6zPJjG7SJ6OEKASfTfyJR9Z0ZRo8X
mkC35YMuMRHuwEBIPnjoDiBVHt7LPw4bSbxuI/7N4zf+griJmgK9zw3blGOT7jK3DmWRkeBKG/CU
C2rpqoHMf37BbctksM88uJ7ZoH+cmF/vbo5dNRLThoJOM748fdr/0J7w8VyziDXWK8GqqtTJWGZY
tguiE7URrEiV1HdN2LhsLIeBS4DKxvbx61s9Wgq0aA6fZvjixJxibuxhoodwdSO0tY5eCV+kAd5v
PF8DJPn/8tE+s7NQv3l7D45MZavKF46f9BaHz8e6ssoHtFFbMJJ8+5/H7hTQaaIfWw3rKDYyhbAC
GufSawBR1iJNlOQO+dve5C4lVFFIsskI4Yi3NdJBtKFafwtd3YJJB88SsVXpa/2ZYAJiao6q+Upi
vLDpnw1ggm4dFYsjZHKSLroU+20rStU1iFiQgoREIWMMpuzGDSju7sAL8duVx7jJlfGWQdjq90Yi
ovSwBHzGP7llG7FDIsQ+bK+ki+j4uB+dTBMcwyo3FLGIlBCv+OGPX2ARPjLBd5CvVkl3loycDszr
S1WfuHuZV7P61I8CiLVw5lP58UddxmJ0YiIZF6CWuw0Q3v9mv9vPAo1prlRKWdVWRwMzK8X/spvv
HpT4zoOGLfBLIEmZxA9wu1K3IXOF4zpzpPZsfHkiF6zwopDmvglLbe/DwzC7gCcQ9nABfi2h2Vmu
qP/8eKD5fjdMIJFxz0qkmq4J2qf3upCFzd2b6dCsQj/zUV8XJLjYGZMl+YM+QNHQlpKoksOcqxbX
oQBXGTsG9YTUXaZdcs2IT35pvDQiRRXczyJsprk4dyALTI31WhnMPS4lyhDUkppqEOPjUg6gXsFN
IeAKv7DIKr9lV2pk37XSk7Igj0DrUU4TXJe5Nm3VP0xcNBvJ3Ht4JRtzPsjn5zcT4o1Dlp/Cy7k2
NcWovCuILwGg2daMXsFksBZ6Mypojm7biNSyTvn4sAqY6OAQF5RDC6VDjXuzzA57CHL2Fos3CBpk
AikrB5WlJT6yVv5Hp/gFCg/ZKFZyE0ujgzvWjpJu2rW9xOXqvdGlv2ASvVY8Mr3YeH2R3vftfdtC
PNupGxYZdtVeABY1YF5eXIbaJ0suCpCnqpsI2eNodYLtC63yZ0hHQrBzrq5COWw0oBJI3I7LGD8C
DdfMSRp2bE6VAVpMIwfZXzLZHuutDIKLTdSdoQbo/oxhRYUCeefb6prulEKknPPuNJelx0+Cp8eY
gzcvoKz+XwPxdfm52IWkFg/1NhjaNQLul1i6dFXF7j+YpjhHmFYhD2iajqWK7XpNC25cY56Oio+o
gDNuqXgvmEluRtMGSLTXGFOgsLQW1IttECiNWHVDAMm1f/c48jIOd7FTWp2910tJQBTupXcvmYeq
HHrI4Nkof6uU8qkzhnJaYrnBZstn4VG3m4roAx0Q9YfiYQ/KFuHDeffUmvHMLPKEQ9XfWxeo/iT2
8k+4nzvmg6W8yRrhJ7fYzn9Y8+wANLLkIvr3p9psqHqGoKxLo3gjlJZh9jReaPzTeLo3+Ac0ns/F
Gfnx0JW8xv8jTSz/AFfUwuVoVdMfyjxbbDPE9fDiFbjHEpQhLCsUHy+RMipp+4sOp3QTniqz4fWJ
uUxnPaZydv3z31/rz10/2x6TZBbPi6VejceZkdzPBgGXzM2Gb5U7Pm3KJ9vUCZtRkR/J7PVquBc8
CN5rhFhKfXVDdWbP6UMKR493ctjlXnjQ9GOa2Ow2IgiLyA4vVF8AUbajAumzQMN0+eBkwncrfpyS
AsNJjivqHwEhDy36yA0GiijQ3TkQuI2nQg9acbqwlyxHPYVY1wTkK36LinxiXKS9QXJ3eVjNY0MP
L7nNwdtDdd60q5YJOl1gcWSoX/9qkcUCLhw1gQK+e1T1GD54WtQtUKACyFLvty4SmtRrsLWzHSJk
LBblMm76Z8w4AIQGWpPPfH5MhCSECWqqwGdMAv1oDu3szkqkH2fKOpTY88pf0ERU46AII6GYF65z
YyV3iIkvmeyJl0bk5p8rkM2mV3jJeTbZSOO09f481eEp7rUp9TgwEWX5fJVIf7jxWVKALuXEd8g8
raLa29GUQbdSr0xLh8t65XX6OPvqyLxjXCPd/DEbap6pdAeGNEbJJToath9L2OTOpLwFiUK4u3EJ
4mgoGYO6edQ8b92atmitcWNLrqo6le7Qdh4l7FhPCO3bCS3xgqgOmFotUadHLF1Ai2+s5M8ChLpZ
h0mCMiOr8EZ2n5EDHlXkAfTLHIEKi41a2yrM6YvheMMMe8e6kMF/0ejRUFr1OcPv0O76yHACSJiz
rgwE0Xr2cmgLoFJvlCl/417Mru+ddy+FXRYV4uAvvgzSG/JF1gWZ2YewvBiQqONIgm6RidH0RqFv
XwtiUb6WCYHy8ZSWFRVCYljUlrpLg2VecnScda35jP1XXfIjvshDu/dSMjTcm/9a8iERWJCPbFWJ
ePJ5Obax+LiK+SQYnvD5JmSIJDFn0t23yHYQNJ24YfKQAvrkYwv6UQJYwvxyN9Yrg1j8v5zhQjeb
mLeqwiMtz2sIcRSS6O5dqHBy9OCC6XXMfz3uDw4okK+pKhsNK3UENqqvlXcPBvyxZO+puvbWucge
J3nM78Hzgk460ciO82yMjLTpqlFVytLHpUc3JuzX5oFBTtGi+VqX5FWh40mldeUPdj73LvHmAASW
4ZLw4Ic+n9YsFw6eIo0zsCycx80XUPWvPdxtIoz9bjPA4JSXv/Tk+3uUdoEQvf3zbpU2u3s4eJ13
mYmZumShY5kAcpBYBgXX2EW0qzcIKDnEzrCFcqsei8iSgq8ZWGBpOb+OufPcemd0aWFJGYy6jgRq
HpOWIZGP059oWjAfnx3R9kK9p2RVCC98UpJuVbY5JC1iyZdbULL+/ggzyx24Ku4HjTrjqwTPCvqh
dTY6HsY4LFKceAEoiZz6RLAM8v96vEdfctzLALxjv9WGcr0phC9t03/M+heCrs8PpiuqIebV2M4L
LfJ9xo8Klt7Z4Ch/lldhgKxLhDWwtQBfQ22HCLhDwdFY3AITpfZjXkI22q9T+yb818c/lUDCxaW1
6teP2ZhX9/hPno2xIYnPiKxLej7ZqaiiSMsjuDAraNri/vDYgLFmsMK7yGK+39K3B26mBZeDce6x
0hEYT0YcvE99L+6CYJoXBwpjclGn4y8hSxCRl+a7Y0ONSL1cfjEnPWBt4Ygac3rCcJk9jQZgDgA6
fQ/fn7FBvLAgAcH2PWsWpkBI6FLQMHvJ1HQInTAobNf2GHKs/7SQ0DQtxCKNuaIL5+d1zcGGwhtJ
PhzNQpWIfpJhNGdwvr6buTztY8AaYGuh6as6J9zxXa6PEw5k0oFCo7QY0ZAvZ4Vv9tEFe37clDAu
K2Dbiek41P0lBLhAyuvTuOgdxAfrADY8SuXxqBQAv+6DEhuBItxuz+8WizcEW6E1gdUOpBq+aXdt
vUIjIUL2oras45CF+h3KLaU3nDQ8jgDZ0kgCjcar5DG6f9qNbkg8cBMdECDEieQFvM8xsogdsYFG
kd+H18UBRbCeXGIj9ZhCzhgLoI04wS7BAkpIPcPm6I1xG+SBhEgeKWI1h0xzzOnuPHsL+UxGM1/b
0L7D76XxLnbiNclePS7/G3n4RAlOnCaxqXJ9rC8C+yGUC/M4wjvN1fVjtaTXk09vVTSbgxLNRGCL
idviUFxpf+rEwt08k2mCSmBqUgSp0pckWyOiTxUH3TkYQg05GjP0PU4yNyQqK1wTOHkMnSdjBOGt
jMv2hJgKVK2Gs/qj35D1Lvwrvj9luC+V6P1AlXnprDZ3tcUWkAZhJXMWK52tqYZR1a+TZELhhlA0
rmcALtmksGfrLVeRorinjL5R3UTBedxGRAokDmqq1+C9VAa03tePPSgk+0QC89qVMq3RrXsmRQ5e
xZLURpVQSF+JtjRR2ZYbKpG3K71Od9sJc4Hb81ShqRkvAVQwZ8jp3xfaCYSeC9TDKrb1/8gugGXf
4oadbg3tgpY9/nCCymNBsoYWrT3hPehOf1Jlo9fndwOcmSv0r/sHvnn9u6RVNNt4gts8706gqgpO
kuyYasiChi2aOZP0YwnGdnSj7VbFMg8Xu+86NYNtj7oy6pEggypnl+HBwBAAr0lSCKZ66lAt+qBh
WPTYmaMwJ0+yR3k56akjq545qtPZHQ5hOZ5qVlhnIFyl6tRJ4ukToBqn0aWqOU+G+aKJzmyR41KP
9wusDCBwIvadu8xKGPKa8njAJg8r2xQUNNh/8S3pIAkUaZjAF7yec98uWxXtmZ+PHCDCBpCAWBgr
W9oq/ShotoT0tMHGsm95bjTc+Rq7wjElhDBt7w3SYJFjfHtIYeqq/+YGqckq5RvbaLYPniiIbZx5
ymYqSzh+p2a4AQFs44vdu+Cz1pBr8r3SESs3I4IfeV/MRf9oiZTf7DdN3uxlvqz8LAHM2FBuCMjw
LgqRGkLnxWw95BRmN6K92s19E6FYLqJolFb82a8QP4wzElT+rDIzXdaQvCfwcXO8r2mAadcw6IUw
377hTbfKXXI3QnYO3fE8o46QFGCbu1wa0XOItTtwuSU5Ka0QGMGX17aLHaQbjB0xalnh1uUzFGKA
QDm4OsF5TS2buf1s8KB4zOCie9NDk2G2SE92iOXblpn8IO//482ZYY0tMRDYpUX+TFyNFf8fPLMg
xyJcaG0FZrAKUN3oj/gNKdqtB8uS9+LSZJFpqsvi8VA0y8/7uapL+o/92vFTUxDMt8KA3vT/XWdM
rc0GnOxZg2ZnWUT29fyJ+X947coXWIYIWF81RmJmM/uN3SwUdtaRWc7yPLKHacAQm8IHwbXBlnfz
hhSyWM8n4Y6CxS9uyZJortqlePr/5wPayDUtdffuhfFb1QLAHNkLH2F8Mt9KgPPoj+X88hWWS4R6
lplA2TNHuTnTyShH307p+KN/mP6plFhQlMFwO5+djq+upq7NELKcQakChk0yc8SrM6Cc++RFIdUJ
yhDW3w+3SqyiiRmT6ZVu48PFVHLZFdaviRqL0ayCuBg4Ya/x8A9uQ27XqyOhHPW/MmClTSSDkX9o
PsmZsg9ukDdncsh8Dx8ZhJxl165EXPlYESAIWC/ms4mxssWimiVkg5jLqoULD85HmTSszZ+b5dxK
j4jv3NOnC/xXjvKJl9Y807S7fE1EfykfNMh23N4rEA4hnxhO/jG7N3zwhzrbMPFHWFZdyNPKdupy
1UoEmppSwIBLcmuwf79MeatCwWW1i5vbUiSkLM3JaJuv1M4kZZpCzFoFv5NntmEbk3W1qzfO9sxa
McHbOPfY9N/0YJ/eVraHLb6/kYWbhIm0SmeoPcS3BSlhrbOuXBzGy8h8kA4yXzwu2K8YVHgLk4ug
yGX43ih7rK5ncRrswWTIKUPeRLlvWbSIJ0NcpwPMrizSBArFOfLgIUbYcvaj4ufHZor6N6woFADR
IKUKo+0GZ2KFtgUdn6nCGUzrahapP45FNQ4wTakG05k63ifsC09RVV2MiPB+KpeIheLrPbWf0HT3
gnEmadw4V/1p08Jj88XpCrfwrxDOpx44OLr6fLOn9pvcQJelIU79nfY5jypFKddbzjzH8Zyy0w42
T6pQmMcs1AtGGSWjkI7vflY/CrEGpYoN1DKRucjcwEAC/hNh2AWXu2NrkatYH8/yrOYeKudzG4cV
AyrV9EAdoGFSHXxq45ODkj1YH+Ol3xwK+7zLCF2jS1Mcr7hFVGHmyA86tU9VhahiLmb5C+lHXwXK
ytiqzFQ/+9Fd0+fVzSLperHtxfPz/WgzCowfLQhsKUkLg17ZD4F4zCpTvrtfnF6d/M8vl9/eK5YQ
kACs+bpHOHuhDH3ne/PzZKKteww4CSMiXjpMqKNczYzLM7PYJ6VrDWjpnNzNR/XtepxnU2c9bP8R
iY5HjkCobsVohUtz3eWUHk3GHwb3OGieFRn2Y0wRVXMZmWMnG2otILGphbY+ZhVP21PTBdsoRBEk
/LqxA0LMgjJWg+6v11/xjpRp5E0UD1sucO3PzskQ4BOtAu0Yq9QPFHtiNDq32kMWCqkC4j3/mPh0
P40dZ0YHnZi4TWOH4Ep69DSpF7e820+KaLk2nMeE0sl8rRoIPEB6MRUDfR7TdHiJ1JKVKUpKT7hl
x7uFk/fkl+a/izxngE9VUz3nNpMKz2ZDNJeC/TyHG/wZj5T/XB2NWQWVbkXdREhM+YqdyFsZ3PCx
ebbcalTC4B/Wj96Y62GxYX33SjLYwuQnJRY658SIt7G90Z1q2/AqW6dxioGn0Xc+XtLPMdVQw4n+
d65Nmv+hNndZaGKZmatjo/WbM1jOP424MvfBdUbGjCqYar3EAKY1YS9RBaOSr57zImS3mJ32gH0b
vT76HlvENUYUQdBW6ZW2ElIWbliHbheg77lqSrVKQ3hpd2aF4Z3Dir8aV+UjECRRpIDGGWOre7ye
rrCpD/ENG216fsa0jT2siujK1+CSMve5O0pMu5HzkgrZgCwPCBiPxVxONxCj8HhLuIqGf3BownMk
s9ctIbo8Lo1HJhyiS8lvj6FFBWCG3x7VMD6HXH4w/ltXkC//IMNeAS7LxwfTxGY2/Dun+xocNAl9
rnavlWe7KVyrHmUd8oDRFrE6U5m7ztRC5c+hCVuUjcpgbajgXw7bFWFr1i1DFOOZn5nOlf3Mggzf
P6raZc+cNlfH2ZhBfVzE6TR4rW6HfiigWrVv+KXilMoJbX/+W2WmwWGuICH0y6HqvrKJ5kKn1Yqd
vBseFIn5mb4GV3KHO8ckdHzguxddjSRrTdf2A2j2FRCT7ZpfMeIkOgaLc6ba8QobxdybCzuEP4RI
REX/yh1+YWgjYjUbqeoKW7rBCy3zM4L6yxDsLKv0PA1unVEI6PK34mP7psQXUqZbUcvJtu4PiGei
a9LGZKJf7Bhihc0OlSTmOc7qmedaAX5dmxtD+FzP5sKZWLAeEFIKo9UNgFdVlY+lo8a1wB0wRs+4
60uL+07tqyFBwbjYi7sEbZiImRarJqSok1+fXUt174k+gRKh5KnYHZ8OTMa8uVH4KcJ1rxSuUNZ1
sfUmIb0neswFMaN3kpmOCAORqNo4zZP2znp8Fe6t8Mq2th+dk3Q40zU3ifVMDm4AKJK7ShO1Lacr
ZXj79zSMciGilvLocivIIfbpBQGoC3ja7YZ4fzrxF8985sBaKUxE6N7zHSuCt4020ZoQnN51Wupk
WeHtAOUCJDfdkQWgzh7CYqC3a1p7pJi1Sne9Z5OsR/HqyJuTgQRirU93v2HD0gbJ9lmwm/p+efF1
3+t6n8Etb1Gc/FHM4xfDWyUQjtIRpKFocLeUbLNo+5CR1qZLUPBGodZeTgrH/SkJPNRe0xeTm2LY
PPLKPGbrC9NWlPoQ5+dYh35Yc0T9Cxwq3xI9jNAgD7PNCC61IhPecTw0iq1yVHOT5Psb9WQHbZS/
XpXcrSV1tcZ0e60G2zCmbcjyzwEGV9O046M6r5zdqHkxC3nH7F0XpgMHGe5WBE3TieFt0zJznYd/
jeZn8fbcEqa64mmVdLoGRSLrNwQJUZFNW4RGJmap55h84sTZ+7QrNtc4MFi/u0s3NJspPP3glSdz
sXKCkQtwteT7/svpNlBSDZ3H2NmUMhnM3n7+YBgcfTPxqUzYt0RiJQ6KpZSCBmGx9LAKiZF1nw8L
GhvwZgyPFvS+MziUfROzfeygImqPoW2sqngzQswCdWKzX3E1reDh66+4EhUmnQac1QDrcCI0s8FO
cc14Yww/ApJu9B7O+hVfz7fY82gOSPv1FlkfFG6zf65Ats+fuNuKCnIuOdcTzWksXi2gPOZbL5e1
HLSxZimxw8mtaGablmxcXXTpLEdkZWaJTTf4Gn3037Byxu9xyiG3HcjmY402uz2Lixbac5CjWul/
zwJBWYMW1g/CG1mR1sQbDo4ceeKiYKAVLqrlCLvmVgFiTa0WzDabhoU8I76bp98NGk4RvTncOy9v
llbnmMdeE4GvrWDdXfogJZw5uxnjRxM2Vyvuj5GC3HJ86qd/Zi2on0QcDZBVznDdu5nU0UlnFa5M
8bgat0ROMjXx2FQnAhcDFNXkgjsxqcoflvKYRXhIpEUZPvGzX70KwxuBKHk6HODNnf7xiJGz+DKQ
w0mO46V8Xxwl6wzZXFn6+s0nAP3RqpYaJLT3jqvVq3B1ZcafmYe5zFsTixsMNRRgvh3lu3+wyEVt
y0OiQuZ4tHn54CwLpdGBlhHfIyG9f4YzJ1kyChZl5t3/Q3/m02/xaOoVVQTqPcSOGeGzG/UB9iOz
VC6m3WVPbduQtfGV1Wu6jUTzrI7d0Zx5DHdRje8rzkkN6FCW4K1wsENWqp83tHvBNVkB5bDvow2j
ksSKKqD6crvxUEMCBhgEbfQvNGC8F+bgj73Ge07r9XEydGdwobHvfe+vejakMsjEZe9QOfzeJO7o
sIrmKkH+5Sie8QUWYkRP6teiqc78CbXY8iqBgY2kVGIDAvex89MJYsskPnSei4mpn4e/XO+xdhHM
aha+25CV6f6OK6aL7TWWasbsrNqpvk0PmNzlxD/YvlN1idK0TstwfhRB2tBss5SN3v10nFSMhJXf
/SI85tEDgdAmfqfvGyG4Hwito69G0wKQy/l8f/GKz9XfOJ8gpR+fTTYiRIo7OAkPLPWRB7MoXfL7
n6etkQmkOyBqz91e1k8YNf2ZWOjxxspttidy9zEBu349Gb/RcOAfqD8k+S84vpiTwwGiAZnGrrJ3
uiKstKq+dVtfgIyBxTMMNcRBZUxln8EH0OlaxicRy/bIwV6RjsWlJpkIY6xd+phprXb9aVCN6gl6
SC1eaMNCEKQEYfOFXmn9/h5rUDmoqGH2WqRDsdzSmJqZKA/c1gg0CdCn0pLKtyyHf4viB78ZJLgT
cs/uhm62OlN/by+cQ/dfdTERYBNId4lx1yDekilD6ocDRxGEXQz9/kI/e3hFcqcgRVbxu45mZonk
KizjepFN6bNPRW6uwShQ1Ett8B+jNJhXmq5zdD0ShR64CAOzqkczpHFDwmFg+8fTDRHFjlSzPo6M
6OUEAKn3u/arazXAYjkCX+LgKC4Ak45nMbyhOmBSq/balQcxate0p03CO+AHDKBsyEb3gQuOjbT6
D+KGt29j7j5JWg+SaoabEFrdmOMPNOq1E+KLN0HA0tEVvCopLHkZJwbMB/thhSEREnjhTVeoA36S
4Zu3vXgLGAEJ2sanhq5Fh5/p1hBaHwj3i1+S6yE/7kTH3OsM8MIcV+3R4ZkOxWDUH7mhHZntnY7r
8Uxc18d206vGrbfGxhiS58aXZz4oraXPPt1M+z5AXk4ANfukrmHg5YQJPzG+lanR/CLFrMSDYO8P
Ysjp0XSoKTMETmP90rTrwl7MQ5kmAu62ywp/zbVCkbUxh/TETISrLn/O7gpuTtcy1oxmWPFTqkX2
6l2DYfzuetbbrsJYZJ4jls6cJb7FwBc3zX3Au64z2iZvbVlEOXRSMl/ci92mz7fWGb4EvooVl7j4
eSalwc5pDv2C+PkEdy8DQAl5QtVSajpu5Kj3PJq1vt1X2gY26eEHRSrWAfV9Ni0Qw2hKaEDO02Bc
wPHQkdZmUAufYhohdgRe7b7eoGO05CxwIIokEWALY0aI9LadyMikLkDK2gxRjKR80Tp1bG8QQO24
akKJJ+bmY4KuJ8ugb6zBfPs7C4M6YYqjt3VdwAzPwrmhCP2FRfCeLub0E/HI4QHN15iSE3hSc5kZ
iH8x3pfLtZY2nxhmxqwULRHyLROFR2t+eVs0eyZcbwYpnjPkgwiXDvFEGS5O+3OXJ3qoc/B/jchI
2T4XMc4cCr5FfCfcQln/jiyCcgd5Dl/OJYAiVv50q9m8pmAhIlgwQw8u5zPOoKzqIO8K0+CEJaqg
SbYr+/B822CZuCMzKjB9CDBSqrNCs9SsC/EPHw5qdPFH2rEj2aUosJ8x/k9yplbu0t7w2UHw/Q6E
1tweelw0fuYmf2IjKRj5x9yY3QwKMUfDR8Og+xI30kgeTPquLEj2PNzMpBGuq7TSp1aDMjZm4mQs
jc5yPho9ZnuIgjBncucdfpCQIHJq7G5S1c/EZOzYLXrrN4FQv2Cw08z+XHvTGv43s7I9Cydy6Wfw
2wvmOG6dk0u/jITkIlfWgMhR135e72PjOZbPk7BWFBkDQT9M5DEga3GaZ2DIp+TBoIqyTDs6drcy
mUgJfZKtGSSMxyxs2XCc4LDKkvo5WAdRqEM8Fq7lS4mRg7gEwQgHYmGF7tYC9KpmKeYP6S0dR7qd
+tGYPPMrDsUyUX7gJtFcaugecUg8zmI6o1bLaefl0Ic1BHClpOy1vO7NDGf5yqmORtYgzt8AOOmS
Ywk7R+EBpxWFHRSw+6S9cxzht076gewA0qh6w11A2vuThubt2lqkyLd1ixHGxY4Vo5F/dy/K0mY4
VdYZZUJ7uzdBXqcz9ImhCas/8flRBBR1rGiw4K3gDTiPzULrWF/Jf2S6+ErtF5ry32Zl443zeP/r
Xu7/ALYdlueIxq2jHvmAQwnymQc7QVNcqIW1ChkydVyvv6/9TvB0DxApY/1FNeUBby9/qN+MNhwr
H/o55CxCtqP/UoXJ5C6BJURDEHL7aEbhoevIpNKLtBhGp0+fEcbbGaln6Ogs+gwvO6GWYIIOXSSJ
aQJeIfZnzBvvlG47m/pPQu9IP/UI+lpAC+3J9bpy9Clpmnm2OqLgHJs+xO8iw1PgCx1l0oVJxGnm
cChyAqVanbd17cxAMtONoKeQ3g7nfqtOsXR1nAqeKyn/H60BU8+YR2v3PhgZEPglwawFvMSwhVuB
5+/BnVW52uYAt8P63vrQxEHPIzvchD7ta2eWvogZPCmPIGizd4VO3WoSyERibKpX7yoJp43SwCME
YAcmlbsWZrGPivrEyKwqISXpHGiGaoTizqVo+F2AGa4JgcqgSxZ9C5JPBHFvoXTTXSDSMlAIEho/
7c8S9/fINuCmsiR/dCA6wi8/chLkEh/zxhRLbasagpsRDIawi7O5t8P17nwd3w0Ym4o50tvqFTWO
V8TbMHRo8F95T+d2hoa4HJSQKKmZxIZ2bnAntF/PFMT8vV2E6nFpMeRWKn+lHoH1fwP7kWkMPy/3
poMBKn0JXKKsR0oR5jnVYVmKxCD4pbCOd2KjXV8/lzBo8JFpw3DABbxYARGX4lXQtiSO3F9HQTUQ
19RIZeRVwkNKSrvCpQkeXHQl2TntgKzQyPqhuCm1GMSqNCiqMxjlGcHbRqLUfvQezQLSXLwacXHS
OzHl/aTjmBeq/kJmS9mH2N69E52N6Ouhx/XO/YlxloB1cER2VNveMlEWRzI6Bc+vTfT3vX7/fXsW
A1AurBDCkammQY7wAmujTljkwfJCXToAo2P1g/S3ZYC+59n/EtgccKds4PZVTF7Ztcf1qZYK52wr
HxcZ03E3fuQ9l9T+R8iVk8trIwMuAOEk7I9cacpvS2hPJs9xdKXybbL6SUsO2S6cLe1CgeJHx+xx
24yAOdh5/ljf28hyLxSFs2+wold5gMAxQBuo2xb/8pViPGZV+kGs8Kb2bviRJrISEzA1V4gAvnif
zPZddpWbSDodQSsPKglge7+KPKR9ckzcgWO7oAWHk4tRLHMaC2eM8ZX4Nx/zrXbo1t3yLswoa6Ti
25ckooAQBRKXuZN27KRiMrRl4L8ux8df83IvwRPCDy6URxIlBaKvjFD3FVI5vxNTrdUeSr4b9Mvx
WRc0ge2QLAJTLakDiM7KyQCtolc1MdSsxoBKmFnM/EVzK1ZegNjSNsp8orqxnKhFR5Cz06wnSfzY
8AwRq4cJxk3NJKKBdzUaDD7cYBw7LPheQGh/fT/2Ki37KnIaJ09Kk+kimceHtirU23lowQshL1b/
9gzwLHuFp1XC+TgBa9Dl2VYf81d78ewIDuSKH+1klkPxx18SsaSXRNNz8bKIfPVwAQqsKYBskR+k
ZxfJyZbCPZDu6/+1QJFbzuiuB/kNDcMyBu2syjB0VRw8CgqGDPL91biXUp4JlhN4wMLYDptBi37u
L/qVHU2n6eSUR6KBoAL1LB0CiXTScmPUKA8Bg1F+dLx+2DrDjWYLrbYqHL4Z5Qblojx9o/Wk37tB
1HuOeZx5Yue9D+DMxAY77MkEpEg5p6chqa6Tq38PUW0XyJHmKhHHguyPJHbzAporfAW3nuQBUorS
R8Kv/Bo/LY9qU2F8yd0GR/AB+PZ0KSWYcZXphswRpslNqAaBD7Q8Yh3DSsw0GIGNy5AX9Wl+zJFw
SBpxAJfzOt8+XPAqxFwnK7svAciEbU2p0RcCC5pLy43yoA8avWyIWWIWSwvpoa6uclERXldRHe66
k8ibv+kUEWUt0B2lHgKTQOoQoOjuaciiGHGRzDM2qFf11R/iqljewp2FtOsracvS6jCrXiBz3B4e
lMGYaDB8Gmvha136/K5F8pnM7ye/8Fv1RCAssgVv/4iLLf3SCzqYK6cyGviI70xR9WwgVd6FDS6d
IxubP4d8gMTiYfVgmJqkWRdIWkLOX1NCPeWn///FkFwsV8aaaSZsoHyQ9OGqTJRsPfVm0mvvwp0N
DArImMgPZY6px0KfPOfXlzSEBmaa9lpf9nocj2GEiA23IbMGgrBmviE4vVs8Wea5ZiRWD2VLWMWC
Ka+nkKs11bzKKajxbXwb2XaEUUq/MfIf/c9Zmf5D3NtVlirZX0X2SsRRK36MNL1vmkRz6RxaHJiJ
2Iwp0TL34VTxa8pRaJNeNLKzyZi5UzHjcLkU75AGviw81MspvU5fRI7b7IoU2ZoRj0bs6xyXwsdD
2WvqPYeFP7G19KLhVvMcX+e8Mf1CdBA+6vpxfqFV9iM+PIUgyG0/eX51gqc9X7QLj/+m86VWmReH
6P7IOYvFKPxDZI43A5E3Wbzdkj7F3NsWoYR7P9B777uNQ2mVa289ITqMXPdPQ2b3R2yPIRjyMxxZ
dvDjwPJkxti8/WbydA7CuXWgqQ0lVQ+x4J8iJmuwE3z7z3EvGGmOJhXPeds60Yy/j7a4IdVFdhsa
wFI7uGrS8Go3NCZCa43Ne49cTHBMeRsNEe0D0rYS9Fou+sTobS1jjBpv9WcgdcFoUkGBq6PpG/69
jsdT1JMz88ydy34++KDUp7qKqyo219igdVcbKQ6PUcLcS2ogpb/vgpMgb3Ow2r39siCIsmTufqRt
+ucECxjBveCQ8mJkRnTR40lKL5Siq+ml3bK2NEl/Me/oT4+aawR4fhsBVEhNE6wsnBZM8guyzZDG
wF+ClgaUbJ1BYzXStg2iK1OmUBe62ZqP00fvcFdSEVkTifyr1CDuwCsl6mUYYiP8H2AZckbxEcxJ
KvekYPOMDHpFHMG86tVQ5+PiK0NP+t8q5DfVNwAER87HhfLUK8Evw5+2pm2w0A/8wuN7GecZa9fd
Xq++0zdoB9e4INcYt2rNh+4VcpmO50BfhTrHT+2JnPGK7+TwrKtwIqiK/LxeS7kM8m/H5qAa9EN5
GnTarOWvBre53IP1WMxAOhSMmEDoX3GC69IcxpXYU58RnQr9lLNhfBSEbWU8kKsqoRjI20rUS0/l
6QEbQj1ioeuchlkYndsbbM8onyMfkVcbdp3iUlvpvLyt/BtNcGLRufMaAwFQE0HpTLikJtfaBgr2
3jAszXpD/Hg2no+niM9TYCBTdH12Iq8S23Gz5KBtplbzOpVFbZGLXfYF4yReCytw1CMmqFhJJtw6
4eMFH+R6Auhpz0bdJgw6+pmNqwI6xL+lCsvzNFCyaX2fydqruTz1V8L1+qWw9OGmpl9Zb7hoUcog
93gDh1CF0kJMPiX3qMJO46QDyn3jHAZCoocgezdwGddi2Y7kOIuN4icHuH8rHqKgjUKmUTmjw+rS
eqaU0NarB3YdzqexJCgQCvony9oZ/Dd9sqNE3G7uRjF4Tvk7+nI1KL0iqHCfD63Yp2p553fQ5ktH
eVX/kuVOj1fJ0Vcz+v4VNrOW/PLJfQoUDyoSuUm5ZT7YhPCsDos58RNBJjl/a0HWK8psd3rxJ5W8
dBNFYvrIqgoGMnSU8oPOT/TfiefK5n90EpuwyqNy06q9jxh5vwda+R8/r6y93QvwrfYPhAq3c1d9
3PZh7tdLbvGYR/UuVHb1ADKfxXqO9dPHzrGy3KTbA9ympUpP38YlwAFY1ionwcKdg8RljwI28rao
DDCJ+8CcSFCQqaw03zJ/BWpGnXASO20sFYw9I2X6Yb0s0kXGOthoIBWpkzeqUemaeGg7zlHkW7S+
MLU7N3FUwojAS7t1nUkyYMo2+Z5HRByNo4Li8pK3izOOyYZwCkOWVb9WpSeRVBdUxRaWkIU64KX3
aOHxNYO2oTsqtGLuVGtV3F+cThp7SwI4RtIFOep2EOI0KpNbW0OgUznpEn2lpTpWc31momH08Jwt
sFEfSMZ8QX2Prsc7DyGyGAGn+/Fnq5IX8VZ4MWbmfooJLnLU6nInbFdcZ26VXe0iFCXnRva2oxTU
+CrtRwKEPo/fgdpiShtt9bPlUDtb9+REMwysTLaqxpt8EGxHlgIlXW/DbPOa38Zl90GjwNgxR4a1
FLsed3CqZKxoB71+vS8VOg7Uj2fnOlifY5m+mLkddD1d65PG9bWcGZHbSQ+dYgCj/SrKQ5Z+1NIT
cSlHy9WSuaKyzNHN6ImjM32XI97WzrbjYFPpAzyUandxWEEvNVHmkvpkpw7HdzRkIp1OAQRmAOM9
defRobjVZpw29a0L+jgRNJxp8LMKBsHJMiaXSDgF2mco9A8Y+tYWeXb1vz4U5lu05ex8jInpXbp5
7WzNBYNlGq66PVRJqJW84kzM/faR9Caogg5TRZNoUzjFd1gM3HoE0afQQuEfRYbJCdaD1eH+ATQ0
4dZ9A1hvkW1khIyaLuXRGegCIjp6elMGhmPqazq9l95ciSH9YbEpTAgj5gz3bVKb1fxPZP/zsJKt
xONDal+LvM0Y61KEzNbZNpSRdFUj47vk9GNvf3STJVB2Rxdsj2Ct9wms9et/3NyXzWbIOV0E7r/1
G2FpAsJ5KT66TpB+TpHkfGyQ1ko0Jcchk3+8UXAWm8r/Mr7S6MYdHsxRiYQ1y0vz9ZRZxRAZrIw2
t5fA3c5fGHg3J0B0Qi/KDk9r0ZdxM2Z/QHxdJ1gyUzTjpx9vzOVRVT+Ca+62ZEB/oy6F5tlC/sY2
cE/ggeENKA6ETHBX3FMzxmPfX7xQ/kHyF7IYUaj4WGH/qC2NLrk1d7IvCjZ1n+Db8wA7nsSU6Blq
TIzEFIZhwe4PxUPUMJiRbOzzfMyg26EaefF22/Zz3FAN2Nzvfx7TrI9mknfCAzSeixrbWK/73y7Q
LNEImKADDyuMtyuUHhFxMIPCUaJ/MHEEIL4t/E9LrrjE7Hi2NWMjsoUfDlvBbarl053NlgjQ3zca
lObd4s2u6S/8POLc593xDyiip2VGNJEc8MQyIiSCzrhiwc1VJk2PtUWPJIGkzfXWkd2rDgQClJ4n
R1FvemnWcwZWvnQP6Ns6WPiUDVXVBhp5nYg+kP9xYIO+Mn8+iVP6ZtsuvGMie9uqPk1q+WH+xu7E
DyTgI0+ZRsgnb2ga/p7mlsJ+zL0OMqYiAdiz5DhC2pd+kOijHdEVCtWeIa6VmKN3Cnlp46NVBeuz
yS7aa4hrWy+d54IywYZOhgx25C20S3bOIfnhkPesvq2nld2ZGWITJEEu6pYAzqAaZhvn2PLNmctk
HNjsAQcv0ooF92BAGP//+MZUwSoPkZUOnTP1NP/XXESyhXeVDuzgG0+vGiPHqk0F3AhvxFDpHWMs
ZhZccZZDXw0is6sSqQcEjPQUdOHMWzUNEMakB1U6abq9opAs/t5a9TpD+xo4gBD2aoV96gw7T9n/
xk4hf9/EhANZeor96T2sgFwmYuj9JAuf44IKOO9yuulk2de6trk5Eok2poXg+C3o0Js4P7rGGse5
4gBSJrCmIoad1yJuu0IZbjy5ZYGSSMjYMmk6vvMnHQYOPNbRj4lqNrxKzfPZEdGKfP5OzZkdPkYB
HbUgyXulOv8cBMqewcE+8U/nJh6HAtCABUrsslfi0D1132IPXx6MCNa2FqucH6r6439HzEodjEeH
GpZeFEgLnhfXVbQwAdzhZ/JCWs7BoxIGx3L4X8/eZP5i5qQQIkjona9zTNEooVRMpsXpLIgKint8
yvwDdc/7+8C+1F/kDHKG6ywHqDStY5PA0aljSjMbMqDiVRnk5i+h+4pV7EAwnBuK2ejEO4Q8lK31
A9U9CbSDNw97g1UJrdWy8yjm17y9DPVZefiJy0Kv2EX+sevs7iCp/bCTmlVaezY9oy87oBAX3aaG
DJsZsq8sTTSi/j1gQH+Bf0m7fgM6GScQKQe7CiyxsIA68fLVwytt77+d2d5MYl+JxnrOTTOkD0br
7oAb2PJOMYnN3QqALXE65jHwB13UoxVuTxw7HcYn56ZF7WpGWDEd9UpI8HdYSZyEQgcWLzSehxPG
a37sMz47TGkZloiUdeD7I0EraFgy4UeDymXwGXtPYnAS8nWSpC5GyDG9zPMbNakaJTlsgKTmDlYV
GWF0oUBQWojHL4iHBFXnviPBFvm+u9QormaDxkm+hHTZS9qubXB0LUnXexX6bKPxg/fGQSCYxJPT
NiHTdJjAee5mySzVfcncisGt2VH17IOUrvoqiOhByAsFHMF+tiYOY5AzcS3CgstsJZhl9OGawA/y
uKdEl4nN5v4Vcr/27WpbO/qXXdyBftuNfYr7B2t4frOhcTFkl8vjgGEfggFT3oAgpUaVX/ujhG1n
2j7xMS9jejSAlElOoQS/YqGPMfpIe/M6wSmh0i2ps02Zc5x2siS8JQ7uKrOWiJYjfaBlG2F5Y1Fe
m1w5NKYUDpga58Mpw9Lde9CwwPIxfSyTd+1oNQOfX/CUAxnk8rolktFDSgM2wYeqZ52TMZRdxZ1c
EjHxXYbfaJvY5lOqxU306hKPjq4mIaT7uyT5klx3G3gYEBhV2ejnCrj6POm+TvG35CzlD+crDz7Z
NrQ5Km0NyQ/7lNoLVR3S+SOSY1x0d2ceEo9FDZm9r5KHjMy7hRW/e/7gmQfDKhMh/y3iQhyj/UdB
dqAa4nKlBdzbJDI7Ks2iY9Kt3UjZLErYJsl+KD5Q+KWROEGosXjuaE2L91TKgN+KB5ziHpeZ+UJe
NNUoH7t5XUKU53iBxgQ66BZF8QYi9nDa/deonbk9AZNa8j9hIFYCU2ydFKrdCTA3y0pysQpB7rJc
kZlXd2UAYAKGkATZj12cBjj9sG5WJrat8zQgHb2mDKzEvlfpOybZ19H1+OT9jwt5Xzo+rXbZfR1d
KKqz/Cny4InNQiGFss1uaYy1Sc9O7Xjc69iZXAYTU1DWbOzVyo+E8ccvRtFqP+avYX4Z/kktLG6A
sdvrRxGdVtlpkYFbzHC9Rum6BWi09WSTqC9fvZB1hF/SzfTclMP8t0s2a++bT3u4adBFrODr1lp9
Z7W3Ay7POp0TgLxOY3UY7GxjIbAQF0nqgIaxKl2VyFZ58iPYWO0d/RFzIzXwUsrcLmmJqJx4nhEr
Y9XJeMUFInv2Hhz83iR6B4xr2UNjfWSB5H7GcgfO12sBrO7lDZHt+Qj/Zj3MGrDwNkk9ePKjYZDV
1jNAkwyQqywjKUwnU8a15bHenmAOEWSeApaoWu/xMtowEDTQ0v5MYDSpYwqF4UFGgugycEM4d6Jp
xISfdUlFjLn+cjbxiK1tofz2bmxqF6cwSTbDrqmXAfsYyqs43n7hU6rgkcmGbDjNRD6SMmrIc9ds
3m6KfO0OURyYVXJvf7coR8+76wEZh6JIC0tigl1zoFgt2+IMWwfdJqNBIKmziNaxD6q3xR+S8X/1
Gwut/AyDwbW6e3LvL/hTf8IdXKq3/2oIjLvJNvx8/uRe7aHc+hcmp6hmtW9WmmJj0Op+ADoPfnrg
Qzh0+022oFBjlYaxcnHtjHmuhLmfIYYxHjixy8ov2UmK9J4+I2SUBeEudYTbijd/pIOu+JvqCbtW
lB94W4NowhCrP0N4kaWKxEe/yRfZSBRTOiAQhRAJxl+BEe/Jh6OPYAlcPx8xao97QjkWvvO3gLm2
Wh7/JNqsEEdqrW111hYQILp9KYduQvvh0qRs9AF5JioeFfDmY2U1ju9BJ+Uvq/TCTD8Yd05NeFh9
xePC0KmMoudFlaAf6lYwnBpWnUu9yoQpekJfQ1A3aKhy+0VD439BrFnpfyJV9SGCMkFEK7Bd+2XZ
yOdJxX/jSUNfQK2jGYJH/d7fmfGmm06J1iBb7evkRwBsa9oho0zUjNUDqjTEbtZtMNNLaF1KFKFh
ddB5OtgtmOVKkyqYe3EuKokqNeaPZ9wHJsiefs+Y2PPpEMuloS2pEf6X/6YGXDOqKRpa+KD6tkRd
bQ0I6ZT2v0M1dUr4etg75zIfMAJWdeImtw2R5cFPhQRMmVahoB+WV5gUyLnKZfu1hEZN3b7ztKK3
4owzogBuq26sPNh0t5X4EiknwNJ6CXuc3rYUDke0KBGsGU42chZ6sapfaYJQEb6Fy74dGfebFP5u
QSmTau75cs2s6zQmt6j9IkehCY8nhtsahaoTRhQfQHIMJpy8+Q5j/n4FsooO/BvDyKZAYhEAwGjn
D/GF7bMoHPuyRLb/0GkJ1MGP0d1razQwDxs1zvMs99TCp4u4i0fCnB2wFZGYGI1xQmiQ13cTOZL3
nBsjUqMIthMNr2kAigXxeUNkANvJvFFu6X7hcqDE2gq4K5W16ZpvdgqBKQeehE5YUNFf4jwZ3ulj
TjvKgkeDFy5CzIHQAiyYTsAPMD0vkg9RmDO5QdRMvGd6Y+49xjiKkyLJtGWbK+6FMXcfE5kYkuPS
ERt5zB0GkbT+WoEXIuFzH5A0pBg3vfSpYqIgY5Crv/JTwtOrCLzo8xHDBVxTS8JlnnoPAdbbe+Sg
qU4LGkZK4ekY4HC71gs17nt6k9nvGhlCj1tfzX+Nd0wdgqr3ue8zL87uYRI11iAxNWwigdhE4gPF
yZ2bOTd0iGMoNKfE74CcHWr3oQfQIRwF+gGCP/slshC3PKx0pVjOyTLW9CN3m5y8BBh/meDkICmU
o1V998hgVCIU2p4KFDld/8bWw2WoKD9lpuJho121Dnp19wRHIzWUKFiH5vO6qowd1sgNUPpprBDJ
2QNZ90qiUayqNxtFGKflXrVap6NWw6zJ5NISDK6nbUKs86GbP+SX6S/ZNFCpuNFgnEyR0Iyh7yAZ
Dmj9hoGasu/vSFAb3OpGtbCpC3Tnjm2Cbi1XGQUpQTifKVifc5xaWgOEnKMVxvn21YkxZeNdEqiZ
NQleCZqlRrpK1zwaGKTxpVS7gLbdYGM2AqhVlXW5k/uL2n/j7KR9+1cbYXp+01/1Y4gWRrLJuyz3
JvBJ0dzZpXhpuMLQkCZ4IaSoZ8Vun0uMCQZF099DI6R4Ss2P9JRfyf2Q2rz1hu3qM+p2zstxUVtV
wxBt5FDqW/1fzM17Ii0dlguqaDHn56v8Hbsb1OkgIxefgKSN4UQbQ8Ta1CV57Kv+D/TKvp0A9FCN
YOuU/ECzGKjb0KQ24fOnT0ozsZUk0GTR7R364cUxNPBpni+MLgiq1B+invvWwWQNaE0+Fbs7Eaiz
7yLps2Yf6UYmw/8rf9VL7pGktoWU1MJQmtJzM70Js2/gYQhNuMKqDcYJj75X1YBK+ogMKswM05cC
fhZVqW0917r5YiFOpOfrn/K/18cFZERWT6aJcKI5gKzMfbDjzKhT2S8MeagggUN6Q4Mv2LinQ1Ex
CyST/YqGvruNntnlvXIrfHsgFeFczpmDC/JgpqCC/KvG+0+5NPnwvYSJDyqPDP7ytjiewfPcgedz
fT0AoyuBPnhEmoYUpKmCToapM2EMHpdnks6229mYY7JfpyH8kgjT7XTvyeuq5ZkzE+ArVUkmAPmS
iVVgQxdZADEEX4LLiXm9TrphUXl8VPghpcmgA6g6I9oJuaLz/61vxwAdzK5GCXZgUUT2GvDFIXzM
VnONVNHlJCSxbPAMAoVe8A55nPnN2T9FdUybNgK7O/jTlvgIYSS2JWZAYZUYx+f74to4Cm5LS+8O
s4p0VmG4b8FHQBvGvEfzqsMeYXbdu+NsXcsAuMi86FFBN3J7DLthnzPo6CoXEVa6bCFSMRnOXYpQ
pdQVDW11ZAY5Kwi32x3+TgdGCVugBBcxnll8i5GFlZf4KrjrcuQAKsdpoaGh6eHzGfgdfX+UxknL
RHAg3NWKxQtf1UrSohsYEEVT9m8pWpdbwftoux7wAVcVZ/0xdLsndV8ONYV9szYMEJp03NoKpYoM
gJWT0uloMUdR2DrhOR3U/W6jwPaEdeYiN/M7ohoNcMA2Xe3/uJFaBf1blUNhknj2oAiajx6fVrh3
2nSFBPZEJPbRgxgI5n3pAmSTrYvvTKhNKYYznnFjOkz8koQ2HM+AN55FR4bGassKsmEVbFOrUm8i
4NXPxJiUfGBvBv69cnAO+UyOHww2pU8GtvXjQp1zb/UVVFnTZm6ke9xdp9/HRL8nH3W9C+cosIJd
I4fDj6J1a3Bk8kELFT/bUciYxUBG9mxwwvA2Uu22q/g2h9LuJHjL4Y7JLnE1NXZJJN9CFCb/C4iA
ciWTFvsHnRQUY4i6ThASAo+Lg1KxhVJvCkvsjpOGI8KvQ0QXmIXN3LKmXUx2BjbInR817a9I2c16
zYMefhlmSyzAcwh2J/kWJtqViCVr60F3TqeBxVg6eSvuRNT8xRURAT2HC7OzEtQCpqmvXfQILFqq
kd8miEoY5r7kvfDQFNy1sHMVvp8P+9XWg1acYBo80M+da/HjtSaF2kj4KlS5RsJdrCvFjgunuSy1
ok8qViuh2XmSJ7aoi3Ou98RgLj1yTesrLmSK3OiVt5yl2lDngPWgzvh8bsMiOFgVVF6NzwntYaAw
njwSVSRaj079v9gjkCuqvl/IdYBLW3nrTZ+euMtNRFyTiUnndWEHd4BsVGBmCi40SVpb77GmJzWZ
iHXOXA276WYIp3ep4Zd4/YKFNPKryvQp6ShV5eW/rl8oJG07o4UQEqjczfoKxB762MjX+w9SKCvC
IQBzv/YgfdFW1clBKg//kX2quHoNtaI2Js3njs8057SuECow1dmsJswoRJYNv6X7SRt6xXf4UYDC
rGT4UqUELu2T+e1wniUXzSnRKxzZLcgwz3wXksyIIqaazmRd2SWECfcZM9enum4ugwjvUIrfNDoX
s/0I66mCFYpCGaN+8XWAmwtcYCZMD72RxiK91MtTcQMYvS1XGys0YlNkbL+iZw5EkpF4aznlda6J
OGFAts3tn7pGs4I7dGUfnDAWFhRsM1dtd4LBTV2VVgZpjfO2ciutHjlCwBJl9Q/F9u8zmZlsJ5Tq
BvybKll+0oZmGdCYDbfVWOvPHNm4g09R/4orboHt10L0W24vBjoQL2+4s9e7TFBGmuZEZzrNRkCx
QUhjXtozHb2rodKvS025glQ2MjYuonx0SlZNM3ivePHVey3Bjnue96CHl5TdoogHV6jLpdZf75AY
Jm5ni6uFatgk3/VsQwHIrdUJlBI+Vz/La3cb5ADId5bo0aEAtVyONwl4wS9JGjjD8V46EASGyvjU
aO8rV6/tcuZFq24CVYk0yHDyBUwIQc2pWeWmBNcvy8i2IBZH0ASLv3bQA2an/Q7ZxslqvZ3gTzT8
4m7K3dIFQP606Qz21Md45p9xoFLSv2EKKYoFJ3C0tmQVeCbcy/gcd9F0//Xm/AXInGUFmTafnAKu
SizEa7FZIbbVSMAYmY42HrgdUdSYeD2v0Pj97n1z8FHhsy3Zc8QvGZIIMI16oPnBnWJCMunYrLXb
dWoTl9aWNQ+IRx1n4ZJYuvZ3XIfz0KfMxctcNU2DiHmSzlsH8HER5V66HXfIhgCOdwW+NGaUW217
S2+uM1XO+vt8vxbM/54mkTmFHf3MliDBvwpWRuTtT3N2ROYRzr5wLv7Dhi8UxtG6szgq5uE8muHV
qbt8bASyAVYAuCgO8Y9HgfxF1Ldh8kKHkaQPNuChFDywMSsPYLhPUZKZ/JB+APRfc/6XCXpQJdGo
iRhu09dT4L4Kzb3L/IoxSfi+rAJC78ildSN/ccd6+/kviYHh+u874EoO8OlEP/VIiiDyQNaYj4Kt
owtMWSELWpvFPFcTMk47iv/zMjGxJILDHLuRLeETD6dpslE4W41O9MYeV0uJOm2bcuH8sL4tIEJ2
pvxFceSWgGtTAVCjmwIcUOwHhhTu/YtSwKPbdZ+D++ekV+NnAqjpwT56LQ62oldXyD4i1ODY6IQ3
xuwFE7PbAxRrgSv6pScdO5drA9N2+9xVazPH2Fb+1P4PkdyBjGDAMkwV2jWxm8yNsuNw0eKVoIUs
D27/TlEvPN3bmu75I2fzB9hhwXSjXv/gqTHsXfl2Y3bPcR5I6CFp7xnWyVKlwcjqZ++l043qJ6K2
B10Qb2Po8T73XC0m7jaSzO2rsbvrdas3wk7mnW9/mXeZcvIo9mHcTMwCThDRS3EyOAm+6yv9w1Y7
lKyeRfVkLSwkq+i1xu8soZim4lywqfd/6aa0s0fObZmMyFOoiFdk0Os63Gr77Ut6fEfwK9+DcRAa
wwhw8+/hCNor4oxdtlPiTtkyLsdAQgGAlx0vxAPFspV8jf0YX4L+tfEpuw+GFzliivs4fMRqUxun
PiZArTnYMBj9woV5Yg4KuYX3axQr5mxATykA2fjB5Cj2Av0L41IFcAoc4XhyE4u1H9sb7vj/SZfd
ifRpwirPV5H/Pm+l6744rneNNRbqQfnbkaFTXxi+VU8a7nxnMWzQG+rOKIx7/oc+hqUZ55QPa6o9
2PnHrHEZpDG8UxjFZDAYWNWAG2SVS3NOQJ9WIxziyy0QknozWQJygtSQrRjQADJLHRwCQ1UGoxpo
63eA9xkjUfvrc7HjMbPip1gkDvYaQMIX2z3OZNm83ebf9nnbB4KoyKdb03FKNMgEMEDDlNVbRPXG
VPS8E+Xx50Nel6V9/aQu/1cM5sp8/wf2pIpEpeVUIxZLmBT0739r6BtEJU1trO+7FGePRAamKoeI
fpwy6P44PBcR8iUsq8JeD8ZynUXbYy5L2+4cxIopX/NpD4OTjFvypB9/ByypIyb5KFIsZh4sNEr6
Fev541aDWLgPKQgzZjwAyr1hBaw444BRgyx7BFo+rscfB1EzegV1pih8zZ2qh7dTI2HuChCJez68
YASmQegKUnQQ7LIUi0HrEkkgg0hqeX1/Ce+nVlJci/5PneR2Sixo9Fo8ltvjhpjbieX29VDzOla0
5rQxU2t/3xoH8NBbe46iYdfavpKmV9CdwQsatul1mLX0IKdm6OUhyIB+VlwhNvmpvEHDvzMiEtC1
PLWSbY9BK54x4aPGAwJ37z13C8G22DDQoQe4uT6RQgFK/0H6fEVGWrsQLQLLWq66UG4dt8msNAOD
MgEyJkrjUOvv0LlR9CFYqKdZcWynykZsgZYgA5PGKQs5xGb3OL3Wh4pGauzf1vIgXRjVqZQaRYpd
ItHJp8SyUQ/wEpZkzhJ/G80TGjeKoyMgRTC1Bbhb98lUxkjlecupIt6be4mgIqN3ifmVmLsAnRx5
MFgJtEMYqp+6z6ZsYueCy/eMzjxwKMR5Iy/+9DDrEcvje9mjY34hbPrgz4CyG8yDPGHKUBZTsqMB
rK5Wt+TmKBalB240wybwfGDavLSW2a9XSHxzY7BJd1jn6u9Tgy3QJ1oUE6iXTNdRE3VIsddNUgiN
zCyWwXxvGVJtC8y9kFsTFx/6iwE8mYhxW3m4Gx7fJvR38+USxIQpCW1KYc6bnZHrmcRV9JDKY9JE
YMa+bQjtUmyDr4ABYinb2rowZyWAya+YeZcI2PB4PtdHxCrNGaaOy48LbWr7s1KOq/7O0FFcw69A
GsbyCY4y4ztoCVoPaIeubUyGwINUphj1MSSAuIbz9psh/TCqjQRyF73QLd8M72mqQA2NE+0lhmmm
xLAy9e3X7QPE3U8u+CjixB0ddtQszOL8p0KEBceos1XXTNvZNqka/CcQMUl/PzzuG13IAudczYcP
3dw6eN3fs4vD+Ni58B4/9fGS9yCmHVpkXnDeY8kFBdeSZiliJpbbCE0CcsoxC7V98s/2DTa+s3An
Jh8lf1EEJVztWY0cKCxqwKB+jILsn1esprtX9iy1lQ6vPVMQ633ENV4XR2bG8W/ZbTuvCHKm/cyx
4yH8KuX4G7MxUFcujNamIVSYNDkuc0fXtKHsMO7zg22Gg5BxrFuPQabSqs+wpdDLK96WYm3zv2hI
7KoT2Fiv0fZBoa6n/j7Jcr7wv1z98ue69eKOeJd5wjSFqncX1rflHpxfDtI0O2b+z/CkoGZR1ACx
XDToQHNaz3Q59kV7rMwGpit6EpN6vF0Hldo6LPXCG3M6rANINuuop0aiI4WZoVCCpHJRLvf3mcJL
h9neayqALWDqZV2JnUPr1v66RM/DV3C62NOhqegZnEIDfD5lwJm/ZYvZIdBSau1fyIqAETbOOBK+
Xpxny48pXzw73jCx7jN8dzYjCL0LE9zfqbn9qM4BxofAebOU9htV5qkZ7r9HFcZ+jDlXMGdHNsYd
0hmR9njLFXtDB1DRiRIMS0gcdxlB1oCUWjBPYM0RAGG10Nn7KBsya7bfrsqg62vnoYOYvfJzmO5I
0N+QZmGMxyv5KM3yUVkG4VjyVEyO3L2ao/uON3L5vSCPTZM5e6/O94EIrzOCQi0tiaXcQ03YTmIj
2MdH61gp1nNPatbdHDflAMrfbTfT0kgufRdWMh0DtGdsn/yxMJ+vRteyQa/YBV9aWZc56TZ7/Uxj
tyYufQxYEFuKSitxDzFN7nPHWeC3K2hLwAzNzm3QNT7cnIblHLnPjrgyiqBlED++8zQiIsE2rMc2
IuAMVOv2K2dnCY9bEwFJOezG5FV3CITlShD/I8evPSL+2lvs6+T90OrQg0yIgaFczRqPxnK1LFE1
n2niiIq7gwHtAElkwsMSZVl4ZdfnWZREmT/n4MOMSwBiSjzTmzVHH3ZNv3c6ePV7JOMJ3XoF2/UV
f65Jm6XvHq99AyXoDhe/jF59hUgzCcIQlMRArDfJvbWtdf0uLTc1UeF8m3E128JjQ7z5+fohYPqj
0GMH5vchYlTPg5QKDeGQEMHIAqZDiSRb2E1DR+92Js8qbY5zfUYJz+e3yrxp5ThIahQZ6C/N4mB5
7D+5Ht+v65/1RNmvlv+GKLD48ig5bB4nu5CyW+t8B152AscyvlvROJzMnfLYLObwq8+102IjLvU8
BxQYrkNv5vR51fCgO3eBrrNhgUCauZMqqmT7dht3qDnjrm5dNTXkxAicGQ0Y1ZV+2dUHA2jKsX80
qhY5bZnEDj9VcGCFdxRHkzzyiG6cN39fWjHnrDo0ojJ2QgIe+JkEN/JMAeCJz4d8hMjJ4seNBCr4
DuCPugRZam390i/TZF2EiBKoicQPPjQ6RH2ODbb8vYunoBryso80nFcKpeCtzLEL1ar7oDLMJlR1
g/4wcIje9FkK4qXT7V3ahvfao69nk5VKutjgPNAi/QPQpqIiR0Ogi9RprW4aecM0zUbRiAvtmrFr
YQNNLuqySeESDoCvUPxLCKcSfd/vu2+rRZZaBekPujqPVuEygyfC4AvNLgF3LMG8GfompQ3epbgS
K7mCFmEi/gy9eIHDitiDsKJclBVcGWfS6ovggKCdfNlBioPkfHiZGW7ruX1QLbIEIOftBfJbj6y5
LMEpmT9ftwiQIOYh7T/Mx28lbt4zk5P9xc9skO1Z79A1ylhKM/XiZFfNVILlYIzuruI2QmKtSlb/
6MWF47gEtkYEq/dWrBCXh5bESiDFrfd68+v/qGCaXi6/OGPFPNXTiaUQW5Ox8z8VSNIiB9DyDfrD
NjQZOqUlwsEq3kLHUVLzjy8EBaCIA1eWIGMIA/LIT8pNodJAgIPYu7uP8TD+nF3/GmUoTDd1vbbF
HAP9Bhr/i2aH7iV9LiiurD0DDPPkmVx8sfz17xazg6G6Yx072aq+7v+Eb0lAN/nA+HnTDFIhQnmj
1IDF8Lz/zofcOpDOm6GoifInkEOgWrrvqwf7NHyxaefzH4bpIU34qPOGezB+M3W+z9X884lrgPlC
8OlydaFklfGOGIH5lN3PazaTpWcQMYGW1qQ8m3rQKXOki/6UVuH4ZhgljngcjuZkuu2po7aiyjt5
3oglwz8VIhjA49G4vf5G42ViJjjNg9mF31bGB7sl8ZBQ3AZn3j7ufp7CsR3fiYsZFOgDQEi/MjlX
GZOFn9rTQpxRGlA9ag2FK/WnZK2eupXQlP6yFMYLT7rFC11kcyS+jLvtuZt8CNr/OM15JjbqPAOw
jJ955B4uSsT6e1nLmnu+wuUdiBy6rGe6rTXYffEOraGWho91hiSTndhDlTynG5BwOVWgtrV7R+et
wY4CVPcubDFD9FyeZZ099a8S/QB7Rug7aVbRreQorWIo/zXr3sAufkXNPxCnsUJJzRhx6L5eNQJf
Z69xM19wY9RaARcybWF26Qm3e81yqA/2Qn1KUM8whQLcChXX4IUyHutCfgD3JwlNCdk0EZSee3vF
AJN+zqHcPf9zjjdb9zX51cNh0YTApbyzuhKTbo25dIBdxxg20T37nUIkrjt5X1znLMzFyP4+TqXH
WpLm9tfGFKmIGRvUHQ7/4E/GeS4fDKe1F8fsqc3knbzZ7i0cbwbdUDF53OUo6sumZjjhRvLTA0qB
Yd8zZIpKoQupSGNhdvFbGQ1F3dT+fKcMmjOnHwp3DbxXiy0E4QIZoosxdxZMOUdSQibhrjp/iSrn
hYvgH4+tXzdh2rfkn1XYRj8csSzl+phEWLDumnYfUiumA7JSiSPs9BPk6IU65CNgobvIHovdBm+N
0lJioQrOFxKsAT1NdM4htWIudPX3SS8yNW2GvuzKxLXIFDam9oEkse/+tUo9VNXIlL9zJB37aP0f
draL2iifJGohmsFqmYR7ywaTTcN8Ko/Jn3pxy8pZH/wqq72BKchLCtOrVth2fHy6hHinLryd7Sqx
FYrAIiLRCX26NNO3yNpbBFwZidEBGaIm6WSoxrswfS//WJphSs9OcE11oIrd9Sa7UbZ+Vx5imZTy
Upcx+pPjM2tXL0m2ZEYW5e+NekvVwGaMQLFIpHlbvDmQxApRe9L6y7uh0QmPP1aSlYwlAJCd2r4r
x0G6i6yzefU7IbZ1oY3LKbochm5VReSurtktbFYOKlCNX+BwVcdGW1bq/Q1SlRidAUtoujBtoHtS
a4wbRHYM9bQrmzVaDL4B6HuEm+9B5nPoHVMAgQFMaeqbmRE9atcZx27EN0oy+SHYTrNn4DYe1DxB
mYVxQslXNxueLlENAI//YNz01ORylFTq+rRQMiADZlfEppq4wXr1Nq9jpimdyhybiMWqho0onDIL
ZtQpmquXDpcxZwkg8Dlx18GXN6YKmIlTvTtEILBPd6JUxM9GxgB95BDfI5sto6vAXzsxZoITtDeS
ir/GHX/Ldtp/4W9xVye6m5DBOtB46mEEeB+tXjEmBnYym/bxOdnbElpdeml4nlSP8Ajn/KqOeOVJ
L4AWDaLaGj90VDtGf9iOllXJTyhWBD07IPZMT2B+6hQpyFiK7pmWx2muMS7GdonndMO106FE1/VF
DU8T6nqc6ti/c32Ns8LUqtnlYGeNYA9yXUOWXuPMenkL2Gdmkub/lGYhrDNymBpOPPYSF4dx9aD5
XqsNj8tUqJVBpaTq1JbQqdd6iN+yY3S1347lLgWWbMfANDEtzLb1snc8S7h7KC0OdezsDm0XaVo2
aC41GHW+1AzhCekBUaJ+Q9Lu+FquHSnTtx4sn1oHGI16GaMcrCbKRaoP3kqq/1/9wxly9iBecJh3
kcd2kujJ3i/2uWe/EErEHoA/zKIVl6yRFZgs5iAnCivkSjSQqt+wMx8WK6m4P6l+z0YGMWfBO2Gm
x/DPXzgevF7PZGMoHKZr8ExTXyOn8IVCYv80TdnHv7PzMuC3+xAqhtlqmwJoswloE6G7PzqcSx5v
4z7tQC4Hy9EhYN6xbcDH/z94pyhG71c/r+60FZRxKmf+WHZi7VvTSZhnG6zoSkMK239/u2UOBPAc
Vo+BB0e6BibMH8d5gD6GyGQD6CPJtpyk3kpivVM8jyTgFookgMxniK/il2XQctFSnwmXyyOFpWr2
x1dmW99dHKn63cjkaOEUJjtr7C/SK8SOECdRptAZvcn8IsUR0jq6uDPH1kW813Yd1t8LyLMUwU9f
UZuXDfz8vig2Zg9okNksdweO5nanzX/v/9/hL8QKcZuXdLDigLYokLhUoo+jhsqy9jdaAoWc0Bj1
/Clb6GrG/8P3CixUI45x6K9cCg+HWdjjHTrcAZpOcqWAHM/LudxDo/FmKyOJvSeElBudYTm2Yphj
TyNf2IdwQil5Cd46NYcwO/EIy3Z8qiv79bAlxp9Of2v+AaIbpXprddYxN/EctHqk+WQAwxp1nX5U
anty/TlDOGtpgEwvBKKjWMTEYQVMr8/bHodY+EnJjdPuo1Oj03pLbkr4Gvmpo9eYuiAsT8v3iC0S
GNpDzMjpCG3IBvPf4gaTBEjBcuvE5u+DCCHYmyCTG21djl+lKLI6peslRWO+U6j6V7OdrsHavcmJ
5cCfV8gxCI7ErXA9j9dwBn9bkTGV0S3Q7glsXp9mCpXhfoE16YGru6EtP4ImkLdSrPevx4uGjrTF
r0fKu/LEBpHOwNr9tIZTL9O3NSabPh5Vd9fv/QmT5OeX52tkLmGQtbOmM5UVmfh4UjPMI+nU4LmB
EA/xnF+eEErm9yhplOv2rHKY8KUsQHP1qUdPYB6AqbT7NYHuKqmvgXPPRfkTP9xPHZ42isU7MqRf
lVzpbgOMQvoSGcSFhTPg1zvb4wx3V3+GCw6WU2HaUGxguqy8lMaZ+VPWMif+rWrlphLdL8I/cLhg
mZl95s9wCn2hsk1yPPx5GsYnskQU2N5seQGSSrKYJqN6SlLWngbxJFYoWDhFOVnmK6NHRyKozZxI
M2lXuV6nFcFTMwK2QbPoqsy2bF90jiE4tF5p8FClomSSWoaQoLnXxdgXY0L3gdqnktdQ/kQhg3Ba
kArppcESmTwUlGJR2MrhRicf02ZtjuoPD7hVL348ob2SWUKd6jWKi0Zue37rcxZOvsg97XOAcTSJ
YaX9a44uwZOalaH/wSSIbI4xOVRtKe6w5qjXd4HEAS9c25AzUl5iRacPFjHczk8lBfCeX7qAFktJ
3PjZxaosEpblwf237Ahy+EvA01Ti+XYQhMFmbOSrucRHnuZ/dIj8HHwHfTytDiIW9VkT01YrQPEt
JfgIH+hyhrQBfwgfAoOAl/yav3OI2PZpJdPj/EYxzci/Re9EYxZ5RxScYUPriHeSQ2zZB0BxJkss
RdRvuVfh9HQh3UJa1hwza7AdBTFNSz2+F1a1mGoO+RzdHcINL8hZeBNoy++LVuluiwTWePRBhF/6
qKcnhebqStDlvuiMWdlPjUEbBHHRRKYeBeJnHXBeY6fiRGnUfoZnSPEs+cgz1DHFi3w18jZNBbzl
3v9T26FGzJylbucTWW6zMa2NsAa/aDWaTLW5aKCBaURjVQj3v62TmzwLkL+5Rpn6Q2AXXqCX6/Wv
hiB8EGI3NU203A71mfkTSHeb4J0i09Gw1oYGCDzT3pkN0kM4HkbEJwBrK1ho+mJ4QQBXYajr+Tk7
cPWQY3Kq3ab5krPwouG4jaqf9W0vCrKK6MuUaBFPDB1vdvlLDGt7FdBzeK9PV1sgwxlo1mnhUCD0
XqqPbkJKvow7FnqYSqzWcUowCOxKIBJpChF3Ji9OEEpczQa9297NCLjsVVEriqtnr7aug2wFhnx7
adLMQvKOqE9sSckCvRog6AQS1Fmu6bn+2Be3/yF8s2hzmU6C5zZXHjckLuEL1G5+55Jwd4N3Ifed
G4s8d9V32Q5CwJOBzch/Aeu7GxH2KXrM7gsnnEEon/QGxdyq2cUEPy0cr2OXQTYg+mR/x4rFB+DO
PURogyyT5CNWEUddJLAIClqvnkHZmJRz5gq+FusIslGOzXjBOQyndsK0jmTrnE+qjyucv5JHrt6r
DxYebRgoSkDF4Jc/IpXyrJTfK5U4ZCkCGkGZWiANYcjw8b5Vgpjy/r4MVZ62/eFqsHcRiyUI6FpQ
h3Ks8KZGDWAbSW4Sh2Ej1LT/lW94eSe764HpvKPx85q5BFW03dWFVyVkKOgXhFLbDQobR5PlyPeV
1bZoxHb+slPe7Nd5Onj0Kh/jBWcWYRXop5alisxwKyOOKjEACjGdK75uY8PnjXfI0loFIi3490eF
012eVUiPm22TyNIHkgKO/tyWf76xYT4UNWSK8WQc95vY+QbOHy6uUzxpTI9Zu55urhqFChpUUfCk
2uPf0hflWMn2SN3+lahv9P1bGgJUfBzukz2NztRE9VuOmALp9/x0lMFEXajGET/UtiMZ0xfaB25x
WIKlR00AGAZbEEaBVW4nAEudl9VlTu8fk3vyJrEdBwbi+OE3Hn6TpINNrS36Q9bzdak96XuCIuXq
SLNEmu79cot0abEaS/8XZV53QR/5v8tehJOmq0WzVepPA25Goqm1oLX6ywfhxfwc5PwX4vdTTrH5
WzaleH2idyQxJYwcDp2+/2f84LGlF9uWOmB+AvtrJaR25emq08L/W2C0lT6QdlGG9kcok2MXKnoM
LnEa7aSAEd4vEv28u0JTGt3vSyl5ecyaD/mNF858XxkmZXUqOLyHv8cPBvl5vbXGTx7k5MimPSTj
XmKmeNfCKcuxA9wn2zEwdnCqX+bNhug59eRZqm5GxOLwKWbSk+NwY2Z8mqEPY0dKDe7qdRS/W6PN
UFXvHLRwLLSp74+8my4xp4ZjEvG1/XnnRKop6eBY2TJ8uW48da4yV37AqqjZlW0P9EMjgwMyazi8
xE6JxCZECHrKqA6ZEp1YoZUmjrVH5TnsEV7G5G9EkBPVy6fkAY42HOkmK3Y/Ausxp8bqXcfRxhQC
tEQnsQ3p/0UJpar/GPH8V/zwxah8LQ6C5vUSXCfo2nPZ9LfQ68GS8323RpX+xzboTNNJPwFd8Q9s
KcBXW+nxgY6n06gCBot5xElH0+7b+ORoeE+ODotqn1ShxqMJ3jmWtWBj7kJR5v8QpfdVPfTM2prp
XDilHq8pDIjiQOT1Wf0+h+ZpQUvv3zBbXTK4fR9S2K0Igg1x3s+jRN8qxOwTWxL4+5l66MFY1oEz
dLeHIXWJCmxY0t6OWQOW+WxwPxkD3fbanlNoPkqtbZvXayjY3jMFFhv2/2k5BIPrauhDSD+w1tA4
0G7/WDHxm9fPnoExDZpSk3tPVEJ/smpvG0eNW1qcJf25E/o2V29KmJZphmoGVIbmd+Xn00763lQz
lwk4r9EXlvID1Fvzt1Og84fsmpnm7CVRftU6UGzfCWWINhbW2uDnu96qbURDXgbvZQjge+NblzKZ
kWuF0Bb4GTkPDgK0V3cXMNMNOqBEoLsMUxSNroX6V2nT/0AxEgQn3EcZmzkJzk046DAbhAzf2lBf
7y+S5TeHM+Kk4vNnCh4oIZG+GAllKcQtIsKvQ6YmEHl79nQcfoMcSjp++t+qsmDTkn7Hj6qaF+H0
koF2owoUNEpW5x9k4hHJ/9r8nwJFfdsl1wlgtAYlzEW9LnOkRpCaZQJdrR+6CjYDLz6M+Kld3hNu
lIjO9UxeMBO6KZAkRMdH6sitYfUM5Xbu+cGUhvigQLkIB8qOPMRCnlDdJucyx0f9mJaQeTPahkCX
q0+Xf6WWSEGmK62SVJeBljQtlzbumlWDSF02ntZMYTziSbh3GYCikuWEUgUvWx09HJG4gmr0FX0D
Z09C3moNRPlpuoptHQpFSbaUKdcTRFjjnxL9Fby4/QD+1asKFyQsrIsxngBFp2g+gYKvjGWbYswV
wU6/DJQhR8FJmifeju3osBFQQ2DiDUTXfje8cd7eSxk1b6pNyF8t2dBCSBRqIEto1OlE6httG111
200TxMnZfPFZ+rSpt3tbBZGO6ZKOmR2dDppjUCObDWS4cusMy8NEXmKOwxhY1E3gvG+hEBv1Ch6N
vDmPJ5ro0Nv3C6GPCqpBr2b7GvyRRSY2OE62azvB8uRB6goofNh/5nMKBpY0QaL4Co7YjCTyDCTC
UxmcN6K/6R7lzKpzXzuv+EouygRPLlv4dWUl6Ks5qGQL3ej1YcBl4h4/RwaHJRVjc7LWB6vs3Lvp
GpQWD16gAyKfiiOYB0dUdpCduHryDjKPv38YhxjsbemHUII/iuDGvKsfbtOIbsQv7HPMyYerYCjJ
+uMCjN8Rx/CQWq/AsRFJ82Z/OfeV332//ng6/KQsfkOXbaethMhCafIBmEgUX6YHCs9x3ZwHR7bo
vGiu3CGO3dcr/G/c7/ad5UinNybR1rDTkaVIsHcEb1zn71EG4IJIyfNK9b/pNhDsa2CbnT1WFWRf
1pnKp4e0lZwuZXRIaeJZNIYBmlNdMx8cb0fXL1hMg/+Wf+zjeGY9WM0z27p92bfDbKn2s9DOo7Bi
ExR2DF7YbP0yYc4A9EfcLJ8Cz47ZOwYIf5o9cf63McvqHJ09LxTz3PGV1BC7VZ8bvJrGQZkVMRwM
nd8OuNW6tmHhVrg0CEKlpi+trXbdqbAEaR4vpZP5AUsr7IABKUyZ1rtMVuoLtrYaV05HmOWJ4iK9
aMRe8VDKVSabAGXGAlWTv37nRWXtbEDDP0qJIPW5igtRF0NPTxpEeJhYN6hpwYWs7twmELjbZQZM
yrzP9R1OXjRG2hmIlKQ7UiQV4GWOPoIP9Y9pJ1fKeNu+QwXe3akDrDXsBy+AyWvVX40EZX2NXs0u
YD1r1pCM9dKtEcSMiFjvwoc+PJdXNXrSyccaSeM7LF5ebCqjxDoXjjNE5FsMGaxXXCULDm6eTbZY
pJIEdn550ZGa4hDV8TwejdnK3NEX3+c1xaJFnxU4M0oVakqodFqQ0J0IYgRjA7Bb6Kpl3GrDJf9I
1fCv01zfF9SgKxU/DZvlAs/EHqQqPpj++7e2IrBg0HGvJy1Gw6Z8UdCU7hVzUm7zG9LJB9rQOw+S
7nzoi8pV2JSilnaOMLSwrpDMQCkJqoHyuooV3Ubbbgxiscrpz3b9LG+nbx4EuCPcYSOLStdFadgn
vULA5k+ruVB8LsG/XzTvpV9E/ICdaFJCo+CFxLPCP1Hbe8WEPqfJ00i81zknmhL1iTcV3qH12hTc
UCTtk/LaIOfKkvB50HlqqmZhRZBTOylwwIfsFyFV3EoG4OF4zimXpRjwnrMJBHQ2VhB1GDE6E9ba
BfWRU4ASZEquSjKoNA4jqSO+KiupyZsFDB0VP6katSvTPS+N+IarhLN1j476z0WQchLJ+i/ZhyBR
J4yBevykQeJgTzaAoxrh86RIhh8iJse3ehUhHTvn96h5pZ2gYOl+O/iP+Ws5iSCFbx1TOTVaS4Gh
YEUJNohLrUSPV8GXNFgjMsNd6XHreLoilaE+riBYeX0Q9nPTqMwk2V7SGsCRWwkmI2xhBKeKx4Hp
gJN+WAcvGkHYmwPUtaHmhFKsVMEf6RTP6WFQrvGt6UEmMwBbKHu3PWbpW9LKySfuf+wh0DNT+rh2
5lT2nZswkQrZRAsawjbNMCp+9R9nnNY4WRUggX5Xa7W2Yq/RxPkvZyXfi9furAxXf1b3Ic87sN1K
vJ5L+A7Y63Qt5CAadiJb6POl6tN5ha1Mz4mNBMttQlkJ2XFV8oYWGgEomPnSXauDuwwvqodDXkEt
R0FeSFp3hWI3RGLWt+nLd6ctLEkREHeYmFgzZp/StenfKzvhBblG7rx46M5Ye3x6W0A//0mcaQhG
8/jBx9I8PpgfGV42iucgjNVYYGMzuX2OSGan2KWuSqAXZFqsxfRSzJbUCUG/oDWODbkNwMisq+FY
taZYf+V3MH5MXKsVHp3XU6zBmf7gX+bZW8zhLwgeDX544vy7If/nlf0z/XSqUkdZZVzkjLqX3CQW
YBXu+r574sM6Ej2IqKKzYBosSxnUy2Cj2ltpe4qjtYYx/+Ev5oPtHTopz5QRf6XZbb864qJz+1Qe
ZcZRYZi75mv19lUaqxmk+fRGlQyrOpMKOFT9fOhc5TVN4UsAcBgt0k/u0mDn2KaYTduw9H+ZlIni
vHUnXbF/BI/D2/+Utqov1MreJ/g80FzRQStrj83x90/sDYieykBLedOXcKAWSRJC37E4d8RGbqHC
i6jkxn3hDxcncP4X/sE6d8nHORoXIfsPCF89h9NMHACbzdDCpQrI5JXlTwA+lfBiELTWJ/gDZQP4
8FL71jvenhBEDjoktnvIwmozVrIlAnYmMyPDgDwix4U/ufjhBkrIRKmalA7b5yI2mMOYIo9YUjpe
5Gb7jzghOPy4adMOatE83MzxWTnRWR9tl5l8c+rSl20RF2LGjAZlL6V6uSfJx+X2LW3wyxkjj1+v
tZKaHfF9M0cIcQhqyyThMvieKkXakq9pd/gm6qJVc6FQ4xvcRGfH60ePjDO61XpaCJhcBo/bo/g0
PhTR9rvU0anbL0tq5/Y2yoSLBuIeqTAlfbn6oDiHaHUODryeEOvdMrpesb09OTHDw+aqAciLpzlE
sLdQiTj97EaC9XQUzaozYA1NldwGlhI9JD9HiS/B9JJxhQqiKSDDwzhyyhw9KFDHBQIvUryay91N
Q8LaRI+s3Xmso2QWa4JwDXq/l4/rl4sCyludOGGE0hmkBQSPNxktaC7q75nV6W8kMxUI48uJBaux
TexOiGYXPnyOIA2uU7EMly1oaOhUpMDon1dS+RCQFx8lF4+Vxa04PdPnqc83utMVMxxq1N9Qnwsa
zfvUp0/35P/71FWSEPiqKYVTmXepJbA88ZmfMsEBEFIROHrr1ogoJlRB9GHHzOe4Qf8QAqmrnKbp
gQ5IVD8HcnRjdZ15tnk+j/SSdNusccf7UPWLzkE0j+oLOhfFmcrLYu1TC0/JTfNKlLHW7Q4Nz26M
XE555hVJx4qLhIO7mkidAA3xerm4suVtbPjPsjZ/hm4B5Ptfh7kgOX1uZJQWwgMdySCDk9GCsV4p
AsOcB7HGvvytCcFh1/M/YXRAbNni37GOq3uHGB0h1/9HMVYlU9YqP78fqef9npRSbhS3/RzvbXxU
LAHWkCEm98nZmngzYnQfl7FhFi0/+A1aVvxBGbXxWzav+0GVPjibbdtbkVJz+mIephU4djrQsq8u
D7BnDOzqLt/2nYuh/Efk7hSdnW9qMFYs40GXBY5eEU92sa4yLDrItr2n5Ga6tQoxNQZmWj/2hWCO
Nd50xDuD754GoWNrNgbiDFgHj8lPc4KIRRtXRKvvETX0sl2q2EChSfsoBE3qQSBsS5clNCIJ44Rf
qCTpiG5XP03uMX1SDkZ/TbPc+AsiK9VYVtHzhYGUYr5w3vDrhY7pnPwZWM3Gad8QWYPPJvPudU4A
KpTgZ0+au3D164oKiqtDu3/Nf3Zc42Sc3RNRHnkm2beg/L2I3Tb0OfRg8NlD+ZLS06Mvy+T37VCC
zopRfQUpjUlbH4qzsoBeDbsqETJZyduHHr+c0AefnvebN3snR78D1/CSMvTW6nbEBLo0rZ8yyerf
l+Ztj/pG18bcGVvPqw3gCI3V8gJZ259bsYy364BqD5d8nX15iO/8Rz2fV9e5/Fi0KsGF+X0N3rer
pGJyzCDomvVQFrXs+3vPHDrutX7Rbgf6JZwFdGd2QeLlg9ozmVbuw7DaHpMInpYI1XBpD5pr/Z0C
92pFDqBIaOE+RQ6MFPYF3EKj9TX9fQ1pBbX4o8g8kMWrD3PAycwBFbfA9eTE0K3KElXRZBFNNqif
bL1qWNLHUJcz6mbDAy1w/c7zy3erjuU+aDqqZGHw/e0men2w/6khtax2mrgjH/Sn77o1HboWgb8f
achBbrJ4fpyVwUWcgEQH8+4cHYjOfIflXOkS+PJkSBN0h91RbvPmDGBOa9VQ5emGXhW99Eun0E/K
FS01+KtQUSu72WYZSacOA2RA8DSXlq+eeQe+TsBq9nX7jdCFTpDY4YOADFC9o6+KEVQszCDKAr5R
+jhGoE/bWp4kugt7MMfe4USEf5UgHLph8q/VT2CtKfPDdscX3KnHK48N1orXGSIxtZbTp2GcKzfs
H82AwqJwCrdqTuCjbhwHsiDyCZuN/A763aaiY1brVr/i+85VGk2Zpg5BQuPZpyUzKO8kIHkCCeeY
P56ZTUZdIYzbcIGjMCEzMKEiu7jLNiw6+J+WGcIoiTJSF9ji+R83DjvidFpOGvTbCbJrWScjFAJh
HPq4a6LMOiBa66hORchIWHqur+GexgsSRVGe2bGzxcM2zbABOue4C8fw4In6mIqk1UC3pXtmjFnr
EeOXf96FvW0qg9RJ8YTvFEP2LU6dSJ8PZ6vEtVZKlg5p7AU2qPa/hiniI5sGZi0j1I5gjrST8ngP
zKK+uOK7X4ZOUSVWu81mc/9Or/oLy8V0s/KSsoMYt7NSXE3VT0DkO3iGbeOiiGxXfc2+8w4N0Xyx
Oo4wMTI3WZU+OSt8SEM41JBfFfmpJ7fhhfnw3IzFqzLbLEdumDcefMlXZkerVD7uPNVkgVI1f6zk
aq4ZKn5IU64CSX1wvm78cEMt7ThlLTmkzqsE7MCuR6XkoXsPluwV6OaCPkiexlYU9oXGVTzwJcDH
ee0AZrB5f+ObujdnUuX0XnGJzm8LdezZ5TNnZGHKYS9mGY+9QmDa0k7Ui/MUjtcjgLvty5wnc9hn
1D3rNaIIjQ7rsrkCNM9lGvLZw4qLYEGQMMwVnCXDQNOOniMi7NeFK5KxxvjUXkksSgxz8ruAJ4bu
1jIjXu/bo1yuEWLhYNM9ZPR0psAqQccJxCTwERZR0Bo8A/2VjW9gRIHVSuoSLzWbk2VYt079KklU
I86DKJRVQZ56ruspP6aTOrtNWVy/y16AIPJYZ7f6Bvp47cI8zgfu28EUhLkGfWbkcIO9eeiFSrdm
cweEmUfAGsDoOV+Kb7lMLRyLlGZ6Svg2jrauhT1XFlqY+nRR49Wp0S2NUeLiC8snhZT0vBJYOwR2
n+50B6affkQ76puuJA3xCO7ev+qDCVrUVncZwVoPKQ+GXltfMvTmhjntt9liI/3FidHAQ5Vv41Hm
cC7en+40cLAF8lpbsrH43seYL9B5c3zjcfEwbXHkLs7FGYbAaa5nVBgPRRIt1iX0ctKoIVnWdGSM
gCqqzZ26URfzsLI7wWe7q9Z2/I2KQn06SLko6Adcb/MuDz11eR9AKzZEtIKC6Sn8k7+kO/OQYKOe
SM4XGwroNGGXk42sdbWvFL5yyc4O/WfOa/O6lVQFdCAZPJOJ+sBzZX/aqFpuTA5r+DoH0uO1UyU8
NrtrZoQpgCjynD5mK8a59OY6Ixsa8veCFjVNszbIWTw4j7RaZ2RhUH5Z9vdQJrJBk4cjOOpDBZN8
SqIxtuI9yeikuIUcnypTtQaUl06wCNDWSj2qwWPJtC1vua67JluyrZL+SQ7J/sTO/j7+XLO3QWzm
oUk4U/To+LsN66JV+jLhvWN4zTE0mHc8HtXiYX/R1/4YKbxiID1VtKFaUxDqn3OwMl38+D5vUP5c
IlwZBI9/hckQDDHvHlAnDDvriH3nw2MByIkjX/1F8oxZqLqF3D7XTRAhfPKtx51UZ+Y0h/H6cADI
MkOT332Ix0rN2B2UAYhyFCq9tNfXamTeNq06AGpjBswjXsg7VgakuFb4Ag0y533F38EedMEXi+z8
RGq5pcshhBHamw53Pt98aSB7QxbH99oA3uV4NqSgK6nzUDa5A4X13ri91xbOCdCkoxp3ssOtoDiy
xcxkvuowNg0XgI/1Yaj+5RYah4QMmGHXIZ9A0/OhlttqXPxHgJAdkgyGJIsMf8unPxJlHtljijuQ
FCjJk8wZON+7DpvQpvqX9Az6aqd6VRELRE1HvI2CRvKd26PtS4JqCFAm063doseR/NVw5uX5YlrG
awybeXmWIR9geYU7yPFooANenOWGAWW+gnUfz1jljaswyzJullvT6jqZXgxjINWQIfAMZv4yimEx
M34NAE+4o+SXzcQeQuNcKs3SdTlwB6IpZQfJdiuC+mlGFUw/KEb/HAphD4w3csP0z+GCqIlzP8rG
pvNXk3G3RFM1wigdIbF2jH66y0CvZnB7SQpBkiXT8GdMaxlO64BG9H7gaD1Lf6n21UAXlIuhH4j0
DcbpIHutkGpRkKEagh5vcRoftdA1lfWnlHLRAWZDZWsqhneeBU1pzrDQWHcrz22y/dWL+SNav1QP
idnoS7vDEi++1rUprPUmm1xzyLarlDOwZ533sthaKeE2QD/FpsY/tG5tAR5otEAIjfipr+sqvfmh
Q+8FqXctBD0jzKbTa5Baaj+dzKFiDQNLU1bru9hOvaq/r5zTpmZZeZEAxzlM8OUOAXuvVxwF3mzB
WViPe7G+MTxal3dC0f1U0vvVvPAvqLzrUWsxjoupd7EgylmUyMIvaVYfhJsPwQd5JL+g2fUoVpvw
eRte9/DCUlU7uLBvKsTe5CrR235aPkLFVWhYPLnstmTexTfRoN+DDEQz4xivTvMXEIBiwWk55270
tbsHaz/AsdNsUqx5bZB4C61mJYrEUG35qbE69bKhNGLYYZjhRhiT086/CH1dk4A24wvycuH0FdY5
fK9JOGT6Y4Ta+i4PNmv6c+fZh61hTlYVL8T/9jU4gVbvP7CDoSlBIX2v5vwn5PFlOiZTuad0OU57
Hu/kz8RStuPTd+IiAkEC+x14xEz0WSz8EAtIveUtJdnuWJBthIxYXLHeV5gkCsCHhP33QiwhNt49
OPy3c7iqPtXm5cjFguGWvoCm9D76ShRt4Xv/hgffU6Xd8lVU2T8wHQvvGI8UdvInNU9906qikYo/
Jq58RS8JlNCXXUU+cQYcR5s4ZlWXclaUpZ9ueqvQNpk8N4K3dcXa6l3j9Ab2pryB5I3Fk5o3CIYA
SczJjz2Egr1GIIHOv9Tj4kA2Yxoj0Toba2LTchYUH4RspvEx0bjZEIc++tQVqjBcoNyB6CfqYLXC
kH2xN3vbMHtss4l8LTZYk1Oyg/ksFv/m6g5Q/hPV6qSWwt5kqzFV6e4sX+YcwHpTp+d/T6cmLK/z
VElktnVGOmkpTRaeBm3P/UAyYgyLTpMLojHc0QN9rmX2YcbIZspfnsCQMkno9aP3h0sLwQ6vlJuv
jIU0jjjglufVGySUFPb+z3P9ktk9ySFVodVQioW1L8owKm0Y1FE+az9awea/9l9jslynR2GuuA8t
2UrND+WXiO8jTGSC+tt0Z76labn6BkPLdP856T7jmDh27acaM2cv/xo3NkB9ZaLgELI0eoSbzyPj
hTGPr56HdesikCqtFVcl413K1NPmMgs02swW3inuYt1/Tj1pSj5tEe4L968e0aFqRafYKEUaHErs
wkwMLYPNh/VsrZgQ6hx+3BWlC93aITpYFr57xiu19apCsT3ecPelzJXJ00KmZ92BESpnkExEbSMT
CCZlbVX4J/QxUx9D1DQD3l+izRXEVxnb3pcTB8sIBwZCk9vMnVQbkqcdRpgC5ZmrmdUG2riY21Cl
sDktt3pzufl/iXvWT017oa6xVHJD76frnoMhCTcY9yLpGtcovc+V5ZNz5ZI4EePvEPZkdSHDmoOq
Nq0WBvd1ucW+FvFdAxEW+jLRPuI2DS6jypNFACWXNOLVwnUKFJGKjRCy3UtdsCIFGO7xSfEf+pO0
+TXDuG1UUiPAuY1LF7PdlJBmJJWBXxARTw5xaca4f1gvdtutBvOlf90GxOYWFbP4bzDQBIza19Jk
gkbuNC/VBDUgGvD77kOnLrpma0v8HLWtBiHdZqj5jOf3rFWcWxsV1vl0dla4sbf5/k2DnYw+/fYb
88d3ZT7WYstv7oKMcTzG6F8Q8kvZ1kJQHje8F9bb/Hk/Gk48S2CjxqPJZrfflJKRuyW1kClbQRTO
uCpaEOSkcjpK/krOPJQpHiJTuN3npxUv/L8685rtkBNNBvtPLL75nj9hGSGo99ftFKwmc3NURqPs
HA9Jyj87D5pzyEX7A3s9zW4l5On96fVgiYH/TE51v/Z6hc5kbPz6z4xvAPDBRt0U/9wrSlh1dlMi
4LNw6cWxb+nXVcBvdANCQdkjfuN/S454/aMLyIAIUWiexBcsUsT/B/2GwPf+RAs7yNXO7FaAV/bB
nas1iyRbx/w4op1m1xeM88eAT//Vdk6AQJn++3oQ34rUUfbqMji+ZTvIZLnkB8+itVGGgIf8AOV3
o2OBfvA6mqK/vQeqqItCpEmzgL4S2hhDPGO8lpbFqJousIvm70TiwON9XOzzUwiB4dXKXAIbs3GU
ZOHQAR3q/UiPkaToCtl9QuFqgGGHZab1sZy+kqZNIjr9dNp61orc8OdXdLV6cfwtQZQA68GGioiN
3C5BIXw+zVIGRnM10yfULkgOHoe4FlGbcpFGzM5t6kiB8i7xBaDbxl3LiesHyrLgjoNmDqyWX88E
tdvnaCWt5ORpufnG5fNHcT9aMOfHjhyJy++F5LFeWocSnJfMqJoSf6Osn0Qg2hrnTwjN2tCJwqy7
bkPdVZeHye/3XF0F3M9er/r4E3r1ccrVuQFUDiBanjWoyIEGeIxVXd0OKAbefNiq9wJWsWrVYkC0
qjN6rTVHGrtX86kARmSmTW1WGdRIZ/kkdg17lEiRTlV/qB0GuYMmS8wkSaBk4y3hbYBQs9diRghS
jdLH7/HVG8niIXibpJZn7lrTnN3b+VIp+UXsimnfx/D2oaO3mfpAwMctjLfQkZERBpmlnUehT8s/
1A2RMLkuW9+LRYTBpgvGDD9KsZ4zb0Br7hF2Da6t8e7sflsAwCDb+sfJm2b6hRfAAGuRF82f+OsD
1VLzz+t0AMFiRLDZWUUXzvoXLUlRbY49FpqHAQwWg3CyW3Vj8XhKq9MTm803Tc7yxxQl8frEGShh
GvlcI9WgZN2sS6XUO1Gef3kvDb1+9BVfZSmR8CTKps+wC5Vmdk4Oo6MS1fPZ1nzrI89dPqSrwAvd
GesaC8moArXG1f+D66gsM9X87gExpvIk+lLi4zKXX6qHkS0zcfimcSzhnf3t92KXOw4z/3+zQjid
Rewjilioc31HDn0e1VhfzTBplL+gcuWvkY8DK3v6c8tcIGe/4uy7mHRWpX6ACglHvcfyI5IX7X0k
VZBLmle4OHBjPa0+KdQCtfangFrg51UdHpggOh3f5/RK+eS4vbcqRr9jF4UV7gv0+KZGKgQLPz8b
dhZ10ftyNdzeGQNfIw6ZHM/1YO/zaHoPgZeb10pwUHCdckT4ZtA0UnQsRHFicUCy24f1nbJbEYyM
qnrSpGXVHupcCvSHu80lTe/EkSA+CPHuU+rVfajLkWPaie10AbsMvcPDY5PpNtK6o3hhvOi5Jc6n
UyTog6I927/DKyDROQp9EHsrRhWkEwUHmp2ymB3dzI1jBaxGGIm/LfL1X3PCaRDTk51KEj+Kuar3
xkvs6R2kElGFJYoQ31PV/etMKYXf1z4/0arFnF9MWu100h9awuldmtqHLQJecBtHpvW1/GiEYaUf
My0Fu50XbKH4u9Qmb0Rm2feQAvyvu8uY652t9XVj0zSc6Up2oUCq1u/51LGs0V1NSa10Uewr4eSy
feS+QWLDe9yUfpxxeGRmrQirOC5ZPbE8064Ja/eQN795aj933XB99cwCBid0O9MMZidSaGEQVmJL
ATt0QHNZgBp6rjPf4UnUXvU0QEjQS1a2ry9fGmwGPVbi6VqbKbxJ7Mr+8u9Z/EUqVhp3R11rD3R4
QQHthdbb8mTR7oj6ZaXqlbZmveLUW+7H4BVwaF3eS2AsMn1bCYkYsRm95rir/kV5scLK8zmLxNXD
PnAUxMBZgDcqgbdOucAA6j3sle1WWNLuGnZLpZ6iR2XaLTHmAYJOAacZjcjpQmIwmtbWuypfjLYM
JVzFoIbDgxYFbAVKFp9y46xj325wEM9fyKghucjYikcn7dFZUsxiuLtPPtW6C745AiOdFF1e37h+
f6ZX1kZRxXo1vUoNsfFKegMpJ8Br4qNf3Oetef7bDOdnE8khrADqFIQke3kYiyl9AU8CrzvMgmae
QIEDkXw6lSjfzBgS4yrIPAs3duAEEyi9UDfdsuUztdHgmNflIgM6xc3bPf8DDit6nAP2zbfDlubG
tWgxiDdiRYifkR6ocqS+sFlgHL5Pv2MRUs1MJyXMeIBj/O32nYwgcpzP75E8dsNvaZ/9GPU1AZPI
ekj5BiyDjpMkbnYZg/0Ks1u5hnuGkFJQap+H9q3e4NPds5H+G1k3ZZST774bsHoHp1iiYHuCwSOC
Kvvppkq1azSr2xxlixmIVdUzFQuG07uZA9636NsOn5UW8dvV9wXoyYnJvAmvbQnNqa1kW9QBt/P+
UqUwlFH+LODC1kSfoEdAHu/93ewfc2k/rFMiuidkAqU/EfIhJlC10Boh3QYU0JLhJbfZWLPfZQWM
qHS78DmkxF22Op3hiowlz+KaDdmYMU4sGEAGK2VJ4NPi1ZS6/4w+5m9Pz5tNHaR3X1p2rkk3FbYI
zUXA5EtBKXlkQJWtwwNNzOhy7jV2FyUi4lYE5U1q5dBRtPFjBlz3GK54MASp6ebkrCzbsgKtEXjb
cdEg8iSyCXhbhGUSX1KZtFjfwE15aTcRoesOheAV/w0NYQsOwmrnoW0ChHUQUkgWjjp0xFyub1YC
E7ENHdyLsTnDG73MHbTghmqJUY9wK4mPduW6Nb5sreltTw+9bEKYtL5H8lWBZVwn6Gc/eKPK1s7l
Qdzlp0Ega5FtiQ+saSGgDD7yNEt8tLxHjWSzo4wCpDGQSwRJYkJVk/wBxAaXbLrtAmtAK9TzaAwL
UI+JGm7lDU5uC7bqXohVXgTmtdqIgxrElNo9DLZarUPaSGkAvnTnlPUiZdm03MjNNQj8VNR65uL0
PMEyddr48J64H8mB+JKA6cpjzbkvbnsI3kbiGCHSCBRTpRek/ZB1TLTxs+3dRRg0E8kUrm98gk/H
8ehFKFv/8ZrblU+m474Z2kMx9Sm9XYAdgEXW04Bq1QrdaC0b8Q4W+ko2fTKPTWR8DSG7bppeucZs
+qivmzFHF6G5BA638q1eQ47FYZHan+nQvk5UDSSPw5kmzRzmpYUNA5fcjV5lAebTxO1+lFQG1wit
xqgbp5EunvDD2y+wPsR73DbQVzxZsZdXbKlPJbOH0eyTIQxU2Tatd2jm1khsUOJGYgfwb1yZiT6u
Yv8mFLavWYs7/9xrsAN+EokQnPjFMu77QnJZnMFHMAnx9keYuT0MVNPCQCPvwTOk0yUCq7SdgL/P
eOicUElCpXQr7OpKvkqklYNhr8vfJspzxClE+iAd9xYNEWwYFHfKal/k9aKyulw7ykimOIXa0UDs
RQIsbIFXU0NXdhUyL3h8S/nRZADsH32HzNTCJxt8VpJ3gvc6IpxYTv6SX2tUKURPSICuBhGGq0Ip
IRvlIuFjuVHUJODEp6h4rOs3xBLk50QgmbuRRgXVW/oKtUyT6zS4kficpAoA1tSxdT4v05nqrQeq
/kCf19ZK/G3lBlZKTm1M8E+Ox/m5FBSO/NcACYCmdcwLkLwJVadQyPYgbchzNpdnY0nDqVgwpNXx
0F9opyFVer0vbr5OjAgL8qMUh2NkCTMRsTXTGf6qf+mccFlJPkP5DUUQa5sJlp2MeyKoR6kItNY/
HoYC12I9LOnoL7or64Ga9ej33OxqjfSSbRFAYPe/vyo/i//wdzUc3xY8SviJUTZhQteqwLRtsVKX
qGNhAkOQQa2g74gszUcq5N4DniJnRijE4HoX1bobOQwqrhO7hPg7O9nsOYQUQ7xJpdGmICfIH+OY
58R8wHmxt7eJA4TysIFR9dBjEZ+biSX1UQqDUiZqsz+R1YRjzJbyWjuPgdBR8Pq8QGDUN01WBvYa
4zDkvev8aho2C1Im1sHoA2uSimU4VvjfluhOOKgcdU1MnBhZZ+DN98zPTN0pYNLcUhUTG9sqDmFU
Jo5xCpzUuXsYZDxZkJCkRK/x5eSVG31KS+AdWOsU7bHGPK2Zaw3mMlkYbfgEJBXh0m38eCSs/vU9
G/C++BruTlFdb5Z53YP5eL/j9jfZtq+9eyR2xI9H/OGV5ubXyedGQoTnilIukb4Rxkqn7aluReSb
ITVeEOoovruSC4UR3RtyFieYwYSQwZQaJExrr87eZfKtBpsX0VsXxNBKlgxspnmOQYDMdPSRvYju
qTw3/gJ3mI1cNTo4qXR9+fJSklsXIpU6MU1n0j8L0KteLp3UWgZdygtCY5OvXkiROdJUXIUuz2Md
aVfvtRge9wSKt69QnI2BSYXylMklWvAKWsidZDXPDD5QUYYyD3Pq5wXkEiBhzOgVpZCZkgBCKepZ
3pVFUjSyRXLNRIa1C5neI/SE+N67JKTH9Q6As3cNzfejsm1ne8EG0Rzs8AZ2uxjAHM4CyGHtk9Ck
ju/pHrdFBxkZ8PpdvU3YtiRTKeB8x1PNhG2LOeJn2tf5kYHRNWbk590a52zwd7W1t8m9jIXfLGQx
Jq+vbD/p2w4TZcYCFCdYL3WkY/HCpg1Ep7dDX020nM3tsZ4ab0M7vLFjel1QAdZn5RuKVsCgfTwd
PvqK2DhmNAVGT4KMnLwjLY6bNcDwo+SYD+0pcNd3Pc3efHYbezYG4GAwy1VB8rWWdZaX8PX4iKTy
X2Zzac1ai/t9Ce7GdQg8N33fBFZvEI/S8D+qSBKa0i2aukTgdYdagqLO+YONfDCUSs0qxpySNGUZ
oBFco/uy8+xILpbkEdHQacyDndVywIb5bvWDnvz3aCZG3DRdSDg59rwfmKzyE+hSpkzYgm7FxTRr
Mu81ZB7iRzMtN9tw+unMcVPr5186V4HPY4w0KeG9SQ9H1eb7ZbtxtOX6ILzlhAht0IvIY4yDeFqR
JHFuxPFhjgL8qInRhRhw4uzJJVC6XMefYxjw66xdE920T1j1v/Lvkhe8ZATtAUpel7RReJytx+0m
kfmMLvoqe2GsZryhCsMmSygcRWwoRkVD49gXJdVF3JByeSfrY8LcST/X5l0rxooo53Wx0QovlGqW
GtbgjujmaiVWLiCc3egAPArK2lLPNyrRD7eOUTPhmRnXDbnWn9XnzSo/MWr+KpbzmxHCvNdOspOk
LNbdpZw31TiUpa+Q4DgUPcLDMIoMT14dqMnEMGe1e8NlUDW2tTNVdRiBmGR3kAwDFjsglbZQIfk6
tbFQPS4+bVavjjhyEPlsRwlTMu0lLJDIOcX4VRNuThBQFT5ResokhVqZCWP3nlk4E5YDsP2FLwRf
lBnOmlZ5mOWbSZZlT3jjvM/7nR1xar6kiCsTRTs1OmpBz5h2/t4Hmd+72ANbxyOEdU9wVuIAy3g3
fjZJawPtndsav64kP2TARkLC9SOidtxZnpYJJ4rEAc3MbJdRXPjuJO6xS2YcI6440n45qwhaVwtw
xnYD+TwE/rTO83ZY18r6CAzw5Kcuz6u6gXNi243CS+bCqYGbm9UwiEJtO5ehzIiggZAwBwTMM4OA
vaOXptkqdIDO/N4g3X1F24dXyo1yX+l/xMqTDuxP0nnrCeBokTgP0pheOaqPVrKiCC6GYcKoQwm7
YTN7q9GR07vLGk0pMBX+H27odFw9oI/f7qGH8326LXR8UKrjuAyJPh7rE3PDKEyMKAhiKwiAzWZh
SfmHbUxZUOpiVAqZxx/pnpWsQLQNnNZ31OHb2ou+v/NF4ZTeLOiHefDZSlWDRCYFse/CUNN4aObT
GtGYlTQa+Jou45uihscLacuyqIdbkv771sOz/hXo9XPSacnW8BcL769xAjaOfb8254z9iYEpnQBL
sZuk8+bPdbp64RjUe6uY2A21J1xPh6wUNRv/JNvlwQOF1vl+Ocyby+6buMiFlnsbavRyymWKX04+
kdk0vYGulFUq57NGq8yzhusEWmn4tZ9Bu1xeUvDj918d5DTYoMvQTqg0763uVay/A3w16znJwt1L
Y5rqa8VKhnfJrGh9/dZzvx3HbKrsnmoCMY0DyPPKZXU3ptnHSwXodY7/BorvXBtDZZBetmmv0cjU
rlUpJpQ84oQhNNDhBCvDKIrQLrwye7+ZpX+Cge9hfKdWkOE6V6BCUgNqWog7BEkAZgCfejmhRj/5
kSmRk57PSl7TArl8ZS6V4sl8gDTfbP0EuTiN+OXBGCWJmg3CydIVVG7pf9DrAPyYavu77PzNfnPo
cQYCm0FEjDrwGJFEd65xMv78jrwoOysySj1izvPYI1LnL6FM9o0ZlPKx/tVxt+qbvxxaK126YM9p
tyv35JEeY9b/Xt6toNOOxnaoXYMjD0fdyh+nBE0p5LiZthn+Mk+Sx+H59EXlHdar9VN+H341nnEg
Fcd4lUuJC4jGIFaxksaQn03M7qZgzVOiDQTWPs2dF2lkKSxRw2wvvLrV2eElRJJXEKVWMGlUN4Hn
qKPDsdh/X3KHvhePuRCFa3GoOh7zy73TxyCZZxM5XzHtJ4H69g7a+W8su5szM/zoti/8X7BGkKJO
2bgC5izK6tesQrL0RIl9nBZSc9BZLshQMH3rxdY/HkCUfwDHLYrxuQbSUJPedqqopruf4PBZD4Zv
gMYZVipiOKN3uN2QmvP10bVKFgKsezH7cuEb9WBF2L6vsSRnKfJC3kWAPlS9oHQFFfIspEYtJpwr
RkUxedhqF4sKIVSFa5ROaT2SHibk6JqeVXuU7WS+RMGAeiVEyX7Wca5FXmzqi30JqrQvZaaFqjsw
O/YFX3eFPuKnSOnOajXkRLLORDhkjgBr+CjslMYnqM1/3hwUKrW5lJh3mtsvc5fNPg2piFPLjeaW
Q7ye43cSxFGKmQ609y40RMhQbNTEFBaXr5xEg4188ShZhk4njU4VgCOdWy4HvhiQOJSk5z9yKaBV
kYl6tKBlDY5mDLEDa1pHyvLAZCMXTesthHm6TOGCF2IWvyDYNgm9TKWVdFaS2b0E4kEYH0qY61Ci
I+RT5oyVTZO6XIb1VhzcZ1NIVtfd+Xw+EYieXDyOcP7BI5HZSo0ysx7GaqmCmH68dUZZYvveJbA4
hShdGaoNFStAZfLgorWVqbcThcdrHNkf70SW4js4JwAdgAKNB6K30nz08FqxbzQ7vxhBAQHg1/Z7
bpl34N6zl8fjV1JLtkKWRrY/JIfysh/xYiJ3Eu31FPjvL6Qeb4XfnkdSKDYZb2T4tEjNaYVg6IHy
Utr/mlKqxOKy4SYrzPXCZaoY7x7sU86OMp0oGR+lf3zBKNn2xm0YsnxRGhNXq7J2EWZXr+7kVkN6
5dQoQR9XsFVrfLFOQolJ66dmX6ziMOc8rCDYgK14EyvTDy6aPgCA6bT4fDZb6y4F40tu2xSAiyrT
zN2NKgGkAJ9EfY6lQ+qtjcNdg5k6KWG5cDAGAebBBFEvC87iKW0FvyjVOWHLdD8UfCO2iLOgZtIS
lsYLsO7IFkLwQ+ioGU+aUncgcmnKe/IIjbck3CURjAJXl/F5Gwb57uTJ35+C01ApATJjxHOuZt/r
h00RinuZPTJeaGTHUKCAjeAaZw/7X/HUN9wOKmK+7NqNDjd/N3aVJtMatfJlAFZbvl2N2UBO4xOt
5OKjYr64GhGcoLQhPCrxM9yJ95A0CF3NU/VOIYR3kRXs0Mr+Y+VhflsWs/j9ocKuA482qPGY2DkA
CSEa4kJwcxBdnnfn889zWTyK6WKQyJKZVNZ37hrhjKaMaB//JBiM8JGjGC+DJEHfzkBw9HzRSKiY
9msOKF9siRzu18Aaj3jehOLu6pCg3Ovn72pyucNW1bjJAoYQHxOugl0kqMpJEsEjVGqpw+Wa6F5z
DFdemPyjS7h5GDiiXeR3RSX37X9N7E16m7Ph/UhQMd/p/ASxWbciECoNKhExuKh62DXDaM1qY7D2
kLgPAVDxfLP88xCNNBP7UQADIPJTld+kXLryPtShlT9wn6MHGDTPSSb889rV5tqpeaUVuOJ9x4aT
3V9qRZoDTukUI0/CxnpSHTF0ZygF5wMLgYNZmYis94x/yEcS6aDbvQ7fPXzHT596mKTszeJ+Nhtf
X4WxEchkf9w9myE6Sk/jiS1UhuegIwXeTloqU7K+ldx9PmXgymMbzluZ+eE6BB+Q/IUsnoOQyV3j
V60ffGc4rK44f4GKxWzqcWu8aF7UC1TCfzo/kQksCl5HpXpXQ2QAfL7c0Z2AI94PPcASPnmEmsia
/Q8HBN85h8Hqb07eJtpKsvkBcCLUj83ZiHGVazebwBhL43yo8JpzlI7/d86vHlOC4FcE0O2UhIyD
gXY2VcrGldmbnPMAb/zco7PAzutkqcDDm5FsYLBLRV2GY1hQhguYD3EFGzSmpRSi4CKmL/lW+gCx
ZIT/lSMmBXBQKEWsy4UXuc27HNFQDGuQ3WzZ+p9q/FLUoPzZAVndMEPcsxw7/E+XAW0TRQDrRyOX
MbHpF/m3v8tdcJLdPjIhtDQUN7l1TojHIAVEkiQCPzweDgRsQTedqgj8ewy/+enGsrReWQxyh0+z
KTdJuOk/lXzQXGXX4Bb3+C08w3xdwS8YczWTDUP1wDsc0i64NXiJ0A/s9hkkyE3XwHOmywSWskVR
8JRcDm1pmAQkKxpA8gSkK268sqPgz4taWhPAKTGi9L6Rr4jZhe5RgQVVPbBQwm0BYrBlIJu1DPHQ
JUJL4AK5hv4gEK1WBovdezirtDnTz8l72Gupd4O8CWAVBUhnADxGX+LzWiasYsoOmZjyS70uq2U5
44uGQapWrEii7EYyS+cUXZFSlfgFdbjbL9+Tjs2Gg6H2dPUifDpnvZjTNgcrv6qGoGECsK4gIdkJ
OefZ/cvOJsfhvvTdTsmIVHhlYg1/cRSN7ZUVCPX+ZLDi/cUdUWpV7RgyI2EBFBdYYQJkwORjLJ1E
y9oiyCFGxzCDZEdP7yXj1d3d/TImWqXb1MuUP8bgSvcjpUOE7NzkAnt1ZblibevKgd4HEbXcxdWa
upFqW5MkOA7svb8x5ZoQWzLbmZqAoQcZ5kPQ5VsS9W+pUZ6NKwxOLEfNIyaGH1SNjCAh69CpyibZ
uPRzUqZT7DszX1VhC7HYS4Jy3zkVEMrd54ETeaPp4s68ORcApM4lGz3qbWpCHzixnQvmY9RBBGSz
CurvwErVBcRIiG3qJjyQ21MPYDEnoQG7yLHARlKdte/7Rei1hE4WLVLgNSxobeg73k1m57dJQZMp
FPom16sGSDNONdW7UP4hDQCXDKKep7fJUQCQaN9WTjU3QXTHybUIy6IDCQ8LKMohAfzuwIZo2xVM
Q6tzDecLSenykWWuwp50vEyfDg5Br8sCUR1ErNPnZKc67byHPVs8OqGiNIrJntGRjbPtYLefzNrt
W0c007e3btCOlm5nYrJA9VMmPBfiZzzRFELDOgQDL1QOGmXPS4XGIY8bWqgUILtcjSc0yHoeVUZu
EILP7tnh6Qr3UXxQpcVvV5+p1ZQGvKNeEGvTQr9QIZcHT2JtZ+ZoKxu53YfyQLwqIKEDm4BIbtBP
nB0IBz2eNmyLinlYIn2ghCtS7b9ndZcNjU8sx6j0F2zl5lq/bQQdnHPNXBnPaU+kSY9fUKyaTlku
hRMyNpEblbGxhmWvCBkPXZkH99dv4Qrizq9z26lKu/wDLV1dhhmqx7vEj/yQ4dSV+7kNkLIZfuCE
AOunUwwlBl5EGaqdEIIa3wsCNkMh3sbevWQIlAG7gCvts4Y+hk3rgbpGdQ0BXTdyTPVr5SP1daqW
NeJKa1/398YOlV0yNE93/CswFK2m+QukNvsib/7YEr7wYcyV/w6MKJg3wXmYLSFyROzRQKPE2Lkh
xz9sZ9iarmK/glPdgekjyQf+LY5YcOpH4EFaGsCGExLZvTxxlYv2ZnlyRBcUq9idB3q8Cqq7PKw2
6YlJRLNLZhVFnBBDXZANSqv6dNLVNDl2hgVsKZLq9daLZV78aa4cbW0quTnQzpaxuiw3sUhjB8rz
55koHfFDdM/7ES78ROdk7V7xHMnuFdVA5+fqQIU301R9svwduWvw5j4EOJvxf2MlXFjiA/TY6ttE
aWKzwzOVk7f2Kb6I2E8+P4uB7UD3iFmxO3LzEuHgjMOOwATt0ClZpVFpat6cLEi2Qvph1Hz1qf0U
txmqx0e0vyZbVyzUAiUwMU21hZM5AHme+IC6PozUUNnXQydkZTrsQUWTzDdS/wyjwH/kvUc945OU
YuElgEAiirTEcN6Kg2pQvVlkhkpUKqC8jtb3DCrK0ZiMcMpPPS7kzoLASdU534jAVUdZFshEkGcK
Q1RLGCjWWmjts8CecdwL2HXWeqAMPFPT7agDhwuMHQLHUx3tWMLd83CSYOFRDRUC0ub+miciBh9A
FD/RR+ZmuaKp+78+CsC7QTu0B1T3TnPZdt+yz20Bf/72Km8ZCkLyXHZ50BCloHqoYjaawJyNgF65
0RaViTm9qUNwqH34NngdXlbqSZNYFiK/O22nxxtYYl+fQzhgc4DnYsU25f7E1vxMIzsjxs2sxn3C
NypgPkJ/uB5lu8K53AKpVNeamBVnpCaa0AacqIc4gNX+joIJLFWcAWdcw9zcjTdBIOBkKlM74zXM
KUwu5nJIpjHCwRyqOB27eYPMIt2hR4UlJAmVzPXU8oYx4YXbJlg+FiBK56W+oUy4AusL0UImAhPU
9apOpwqgWgndcvx1T6eE1sawSStq44rBNifqOMKGdqfM8zjGKZeqk1Jwnuw5eNWuunJmXtm/jKAg
AUYQTQ24NaWvJkFo5yOb8jgvpCWEc8mOGbkuZFca5sQV2rlGQc62y3YYcOyrCaLPyL/Dsey1pG9Y
mrC4drg6T1rqeQD4g5IdCvLY2klZZHLOX8xX7I3PcHfZAIjQi8tZlLdz4w3YC3ltODOwl9ymm0vq
IZIa6IWUECqWAVnJMB2T9t10btPwjTyIZdsSkBS56xtnFT6SRkJH4FcX4leYMjNrGtgf/7rDsrd2
5Hdr8UaEC2JvoNTS2R/yhYOSiKY4jnKp36CFwAI5luB6h1wlSIYLD5FU2isejLvHdQxWC86dLuDW
sAj42dftdljoUWrQmHzqYN5YW+cOKkq7j1PUOiwPjUyB79hJPWCtlxpESRJCjclOFlXEFz12WTNR
WDyV3OUyW73hHlpgR+qza+38ocZm8AwACyYc2xpLByLkWArRIICnwQq1tp4ezNdrPLIDxt7KmpTk
arWndkFiFVjFW1Fj0OZn8CLFE68KvPkXIkhs1Iftm7Rauf3GTNq9eL4fIB3cRuVmUv5+wde5YBCO
wPCzGUNgGubRjbnpuyjRiNF5MqJ7niqB0wn69IecmJmqiO8PrhPWydPiTc7fkP19osKdTvyEDS4t
G0825PmJ/6jwAcX4Nu2OfHx2qHPF9/HuMe02GEzB5Yk7PforNQZuDhWTG1qNFp9xAIA0M9xQe0Fc
gTICert5rGRdFIw/KwiOBaumfC55TOhKBC6K3A+O/Fir4rSmCRTYeGehpLsx8yhXGbsp7i3IS/xz
OP2dhBha0IaPM/ZA6olZv5fILmeUE6LmFUdsstvFnpvgAgqyR7X+I1biIYmiKOqV+MH5zmKUQc4/
228JJABC9hmtnNVePDtaxlg9Av1UeGjwT+EUOsdn9j83C6Z4ZL3usoDBTjzAGitOOb+9QYsWkcVW
3oAo98PMCZAvsQQ5wg2TmH8MeP8Qgf61jZMnGSim4vsAY3Vs1h/kKieuq7+GiQs+1XeaX4hOrsCl
LFfQNXZXBmliwBjteQFXF68aJmf32Zs6Fgc1cAeg2LifCuK02HIuSLf7BrHaRS5SfEYwazvbilqv
n4vmgVSkQwuw2IJOlCRTNinXAon4LGC3YLRMNFXZdmjYdPY4mzFF83LdGF0fHnjVuXBpMdv8h5vZ
DXkm+H9ittCzTV81CZ/PjS7ENWDoewLYKMdIUhNv8b4Lla5WeMIAJZH+gGZ6VrrUZQmTeprWcLNJ
Q7t72up241V77cDUJAhnm8/oiVa9dgEPxGyorf6TQRSLTJ9mGAY5w6Gq86ioCR6Fm7IuRsAyMSbx
doFGjaya0fcumIl5VG+Y/6PgkwIhAs2ERphgpIadcqsHyqrm2KPrlPX8c8eOhXN+FGRW1X02xlza
cJ5QovLrzCZ06ZGp4yThSqZsb1zJnmyypqG8GALUOKpp3KO1VUoNK1RoLlYr5Z6mrU8ER92o2CLz
ouD25oEy2izI8l5kcL0xQJaZ1rNs4oglgLoScqyV68s+OUIY6DW/auxHjo+vIK4Nc/27wZEakmMI
k9rrym5Zzm8oGh+rR0iCzCDqbtULPNU/48sR2R6AmYcMhJnD9ZSIuqz/vtQeBbfglK2lyVXIOVH7
W3WpVIZtW5s4zhXi2o30lsblAfU5xbRkRv+VqTqgNYHOEuI2K9BQGL1gwb+GWrL4B9bWBAgfRMlG
lSjERl8QqG1WWcsTA1ahT0NQwjWUpQw82LQZhTZZcYhfN0d/qoTiC9627Q9Nz1WE54SIFNduyw2l
dzJNPmkiV9DzkeNS4CA8hJ8C5o16YIE8FekRZUQtvNoxs4aVmvpOodt0Tgyh1nbb2L2j3cKWf53e
Vec1436atGR4mopini/zkuhINqJHRWGJf3H9YN/1+W9kXdFiNSq6iBTowdSUYPWb38XgR5X0sKmx
9XFn14Ei8eIekeEx59W3WMyp6eBw32VWxOn/78ijpGsc01SgkZ4uSwP6e8FIQ2vFWIwqRQswkE8C
VcgMG+n9uqtxXtf6T6ImJmNtwxuLjZNZ4U9IrWhvjoqDsBijp0M9u7X2xvw8ICeWhKivNjs+B9sL
0r6MH/tT4jV8N2kCBXNAHOLNnWGH+IMpYuFB4AXOXOsQLKYeXYpB7RtvskshC594R2cQNkGuv6SW
JptOriuLkwI4J2DYZrnQkn1PSR1b+oF2df9/Mj6Fu8k3j3JqYcpaiZnmNiKIBajYdD9G0svGfgpG
DV16FIGUbXvwOxfl1e4TYUSXmQ0YUSlz8UkoX6n9QUMDvxZ/0d/GmyFJacOcQv60Kf60k0xplEhj
7S/vrCbV86Bqk4Hi9un+8NrZupHlGWmLxnFUfQ9maR34QS7wrZsS2J5a/wrYQMCI29LWmGmDeIjp
06CqUyCZLJD3o3Df9z+XvBZim4dxNuwNQJSQs6FX0aoXVegnbiJJwdHx4PU77IIwDYbx2+QFudaZ
DIOd3pVfOw2LcsOM/e9L2RZzui7RB5eA/87V0c7CeYiFozxSQO/S3CKE8rB5My49oWXiGMlDlQj7
IfmGl52qxqOQIXdLCFOKKy8RGR4JFtMALd0c59fbdmxAFS+Mnp0KGILBmOtxlA4LH4+Qvr3ESPiC
OvL7gcQW3JJMolO/S327spUPeyrZjzU3qZotV1VLt5orlX/RX7NLaSPRpsDG1U+n/QskHHVJbLPg
BjRTp7P+ASUSj7LQeX26nF402S62vokVEr29sMLI/xViCGUjF4zh1G85SuW+qBWQO3BPs4EIu86O
9/ZIDRU/NF1kL3DhmPRUeTSTV4S+FTP6V3RMJ30egJKQDcLqniDy5cXniTSkniyi4YOcVFrYb/ep
UBetE5FgiKiFf/Pv8hyzqbyd3DVYIiszV0jipEarw8ZevfIv2poU7mVjMTnRLIahjh+hnJigxla5
C0KLBk0vWO0u3DESz3axjzvU9wav3KhxX4CElpuL/2X56O6aYmTiq4itzrVI4VGzRCytSnme+VOW
ULTwJ/zWVA4sTMBzxaDRxtud/dau9BwzGCgxBixCKU7/49PAiyRiVqRcb5sk8VLx9kOF6EmsJM+6
j2npOnLSxU3nw1H068w3oJlsVTMgD77NDESTBDuWONvKI2kuDsQFvEKjpJtxWBzajfCArzjGUsgd
bZI7UBmSwKJgGgkJPNgGsdBfGT1uFO1V34pEJkt2wAav63m2n0KEJIJDQfRQ3y94HuRJUtaXaqt2
4lI5/MzDxppoq/SDI3cZ0aXAqquYAJWZc0uM9/P/grC3WPAJ8plxWcDYtQWooHXXKEIpf1wdb6bN
QZc0GhiXIdHSEQhdx9Xu67/lnHQkFGgjcZZAJVBY4fd2btuYOfyNp2IYI6vwjsfa9DclGpZbNY2e
OdKdGL2wtqFqVlQU5k8D+xY8aYsHu3N5TSRaMj7DP4iymyij/0fGihOda01ecByB+B5S3BWtzm/N
HzVKmmmlkYlODh8qtFYbaKykV6fPq9vbjei6yB7poy9NYcilquBg5mCP/Q+YohMHi6EXLvGq4o9K
c5d/ixGPBZLEQQrkwZCpuUJYIgbOAvxBTNWcCgWKV7jeeeoWvlMvMUoKhmEtwVsqUeJ5rQQ/MdjX
Y4xqzmK76pxFyqm7nSFXHJOuQ4rKawznNkcs4R7irmOSVD2smoye7Ba+nGyVw+2RMDUTWHdZesxf
SRUWt7fabMcajm2QGnr7UdARjKQqNZdGP/8l32XcP67W8QX5aIf4owGquShaCTIbQsbZB6TzGaiG
b7f5bpcfPRCd+SxgxL45fCaEK7Mhn8qJNOiE2524VsLP33fuTaKV+D6Qo8Gnxge4MHeEfKwycVt2
Yz7Zg8OtuBSo+peWrd9CKwD4Mdo+4VwgcV2jeJTXfdv0x5WYELBXSjpSqeKO80XQyN2KipIpU0jg
qx4iCu+1B68pOIqKcrbKM1dWiYTV/ooyeu1oPBv7Y6l1o72KUu4Xh6kMSd8cxleplQ2lGKnC17C8
gpzaoCA6Ixe65l5+5F2HD/DKrGGigcK2AmW/mqucV7uvBLKpN8hMIvVTmJn6KgJUPKDXwlRdJ3DF
pWNJufrqwtlYM4PccDjJwXlsxTszeXlwZosLHXw3UWFM15hbJllDDXJZ644c1ykIzyMM0Rai1/0P
9FHeCaxXGVlNo8BXNEYLbhdDtHIankYrFfXzW6G7DT4h/DySf54lhfzvVhsApX5lYFuLsLpDXQ8E
Y5eYM0n5tbTMiuVZp50y15iwegu4ve06A4RazDVmenq7dx5vCWEYtokDk1UeQTfbH72NSBeQplHI
6Ry6REreOKj/DL7jkKXsoIoCzZnN5aw0uDFY9wyG9gR34isH5RKzOtIL7A0FbepEAOUcn5fhyMY+
qOjQAv5m3AVLXqjg/EH0xzIpd5b+v0zjYStzwkTBol8/PxcTg6KLZyXVXlGVn88Qp6u3phW+qzbZ
HsihZRFtK/3PDyk0/mz70kUtkbXYYYO19INFHvdgF2ZeD39C5+BjOs0zZFrBXLsF3WckPJpcK0++
pDB0UJmU+ddCmvp4f4JT3CpR94acXLAyLg3p5M02zyKr966UBSITqZQS2FBjVARDg1DyhRkSI/Li
COUpj8X+PgsIHiiX4ut3D/0nSJlxrAiOO0fDz70g+caIsKOt8BmBYT5i750FJUZ5Ol8sBUeDCvg9
xOCeR7sId7rwg6RIINxI/24HsTC4Yran1FFekhAp/1BVv185nRlkE8Ti55uRoecDfZOrNrp1RZPV
PsJsWlWbX8fploh+M67efFhlxv6umkN5xA2URHHh9qqH7nDXXl0CjQ9HZF6ihI1pV/9Nb3BGnIwn
vNI5M/9Q1tUTlC52/p7mneD2IV+c09fCBqPT54dgtkVYgkIEIcBCk1st+d17hrC0zzWSqA3hNYJ1
vhiv7HnRduJNVGAVHxbYu9bsFmmqGuY8sq8YzE75b1OJKTg9ro2R+acpbFpvN3/KIA3Ng3c+/OsJ
/Wk4epcKrafd1xF6Ni5pCRuwJeX/dOSzZnZrmSFAuVl6NBy5TSTqH1O84adBb3ZAkAyt6kXqGtH+
95u/5IFlmkgTAHHa+W0WlqGt3VUao/QGLv5F9uRVdWKrh8rMt3+3wmLtmYyTNLRn/KK11nGmR84b
h1t7C59u73VkvkJvsJcrgd8FR+pXfwVJmGbE2gE871quuCMkJiBYfUga7FYevJenE8hT8FZLIooX
J5uDiczPbjyp1TJ0kv1dp2UB9el2zNMM1Bwmqgr8q+PM8rYT03OdD2JkO/pptEf1y7+gMEbXMlaO
wOdSpwMB6dDEW8XTfonXquo4zGgdIcuDXWtScXz/GAALTJGHp99T5rKO1bmhBEXPkQVd92HWIEtJ
pMXFWGbB/+t0eLM8uPU8EAgckBYDxuA6Ik5E5E0jLaon14ppLHVr5xaNAnozBlQTPUHbwwvKEB0m
vdNaGgF7AosvdWvTCCQdb/BX+erYWqVcVZuolH4nEv09jQkTMRQnE6gpN1Ea9unMK3lIXWsPlvA2
96K8b0+NH5trbqr/QeN+TwWj50oAVAa9HPYl6KwuMIy0XYORjgYRtVfUdn+6MMv/PEKGQ12yqDvI
6GdwdaOTctxdJpff8oj0GGmv5kPODHX6nhPns9zHQ9sCx/wr6oJOIBWWVRnlEFY1w/PgoGiCn4g8
quN7ZtOk9UZyXR8zwiMVIxQnz+3TILKNxIgVnikwOR8CT4MwsUb23HdXHPceyQYf3GpTPnQCxP89
3ccONPNVmv3c/aRwjF7Vv/4ToTp20Xa0zmLJ6/8jCZUVOqdDbsuJMvwEN3uW7kJ7QgiU0iyKOqRx
lvts4pBk7A37cSsfT33JYx25FkTbQicXq7alk1HzmZRnMFxFuCih2pvQZoLSWF+9fyzK8ZPAaiUj
D0ai07E0CcYsgKXIbc/CtJwGZ7zQwXQoe8ULby3zkoeHGY5XetrNdcEzHktEjMTubl3Gxect4lf8
o/XOyOeAoJ3kE7kJUSs64kiQAa1CgJVZY4IZAcjKKHjjcsTeiuDDBPPb2MlfB2DMv7MWB7mcJGSN
WuaXqzMfcLhOA6JDswtrZFtUV5hMYf0uwh+JuMIq5wAH25su9pjS5RQYj+dtl4I0TmKxu56f0/6D
0cIXF5Vss36j2tX1EpUu2bcmFnnQ7FzoghVgUD69IO6w4yYRggMBSzE/TtqjPAjApTsPONpEYJc8
u08dO04M4gJnbfbp4SOBY0903rPm1RCxpWoSussHCDwNk/0ncignTd6E4rrm/vEFte6h+wuyd+tE
wlPClv0Xc9o7Z98cr1wjyyUFZooYXkPSeAfT7fdVjkS0ZiAeGYUlBje1sQ9Nv9i+8p47AM3spjM4
5GUbDleh840cBvti8myB4s1BQH/NjkPqkE89+ravZ1HJbXxbTmjycJqHCAoWs2kidpVS8CyWfZaZ
kgvblVRqLXdFfAxaWp/fCoqx2yjEmIHPfpbhyhVelMkWQrAtjbTzGnbYHA3ZjenorDs2ATNtyCW8
N1/m+f2jF9VGlkGMFAOAkE0vvupcs/t0oAmK3XlCJnRlBMcCUV87pB6+0rQ7mBny/e49vya9FPEM
3XYBd/tCu2gzpEkkFfCaFXUEJOkIwJlJyZ5sRizpuJmQw/urNBlMOvRN/kKZdBn8ey1/HE2f/V3j
4qha4qMA7x+4hNY4ZodaHl8NUmcI3h1JiwqGWU3kAzopEXzOtFi10t2IWIW2whj0FiJ/PCaY6tBQ
P0PjTBVhlozyvI85RNUdMRdygnC9vM7fNCZYtDIjxkxMhYr2qSsmXR/7Zc5wJgC+5xUQ3vqrdkXU
5iEbkasED8uDwUcJTmSfNJLNG60+zZwHHI8XOHVEA8e7RwM9wWu6hsqNpzHINXyCDf1eUpcflAog
a98Xk7MlXYO4bW7RFtiW0IJiY/da0nYfUPOK+KSJhoOwa5Sq4Xas01TsU6faZiC+MP8FJoLTZ7jq
s1dD1t2+UZwvxy+vWS/K89hBTNlkB7cG2xwUE+z7e3bQNlUsb1K5M74P1AdieQrLDeQTAKVryIsL
fW+9DPCV9hgb0uUHc9lUMLe+jy2BUD3eMuooIAhI4+7MLfu3MtDESrHMyXBwDsc5KYOdHzDOgGDF
MZvVptmylIvHT/PlITUcQZsRlmbFE8xYPuPbD/nb6IknyPEcZabRwVTF9/ohJ6AC38t4P6WYjIo6
NZbFrOQ6YYDG5l1y0Sl9eJbk40VazdzTUSKH9cHYUunXdRodDDnEWxernHIFePHYuDSIcEyE5rpI
3CQDkWyHVxjTTeZbJ3w+QeaXi+02L+wMAKUalARtQSpM9CMOlsu2WZTOpaBfH4Btf+nkgu9mTqIT
U1nc99btGXWjHGiG0k0v+xyZz6HsFJiR/7Zhh9B+eBjyiclVYD/+unyiy7T7e1eppXA9z34niayG
unPzjdgKf+tZ80xb6s7eP4wZLTSbnrhykIOejsQW+scxWQSCOeJ+PrAHBV63AyZnWtnIkuwGuikN
H0ogEwbmSUeokqzvHYl5ldkojCVmX+4fnJDE0lCHFSfjL/V71tJTxvAFuxjRrNYCStfPvo2h7eOA
VD1JD81s6lt5rh8O251KkNn40GbktMGJ45d4Mi95sL1NykPi6FSi1eY2NfnuRomMQLNEsNO3MMDT
np8XjrC/njX3UM847zc4RjLoO9A0gPBOeiIe21bwswIMGTejP9lKb5a5cKoOS7QYMyF1vhZiPThW
AWepNzzaN0LoNd/x+q7ZKO4KlkxtHGpWOnfz0rZ1J/3Qz3Bllk39UuQGjV8ypWBnaHYtslYux+zd
vxrELgs17dLhRn7P1beklTkmSm46wsSmJ2QeObMbkW3Y2W+/1rHGp9MA53BLfUNTHpwANmmlIQmW
LDlQ70oQsLO21l0Oe0q5BJlVDF607oTMHSUmMTzU8mkTGglsAXQNggKo7+lFpzv45TVaNd9yrM2b
sYrVT/LKU0e1EDzMGITTG2hvE27/5KD23au33ICNfI0BY3eWk448zJGRY7ONccUswOjFkP/btuVb
XH1BNZlpNuU+GNyFF8g5uZzja2V+BUvQIq5SRooCF6i/BU5Qi4lHe9BqH0M/jlZpor4cCo5qym7K
7YuIzqKlNmDz5NuRthgLsNWVyYcV/MwgGJhyr/sz13iKiGJTS3NFVzPNu6DeC1CsA+u5rPFQfkoH
mzlqTxFgtQTRsO9JSuIarVeJpMXiCHwujxxrrYw75iMc/Y/wLZNsH9bEouBxa3/rp/G3xl+MWWsN
MStuhHahobB6VvAMULwYdJf3jbDwyy/VeukiYP/GPG4Vu0PO+3+wPqNVdXQlWW8q/FraoFlcZ4Kq
sXqrGZ9AUYRa6nO8y+v2kCJ8PniUceo1XAKPfDZf0EJtHS/6YDMsX+fjRu1EW6B1LT3Z1rPUPQQj
tRkZvM9Jt0L1TouLHxiyiM/J9vChxY5ILYjW9JJGL4bp0BTGcbTLLGWoZRn+Ee+UqIZEnzPAhBON
sdImWeRgsAHL3eSlqGEtn7Kf514/mi5aS86cMO/xM06F53ZrB62rapBAQFldLLj7bOo5NaFohAaj
NOvjCn+ORxIbndxaQCW8z0crcw9N9Aem4s+8tsQvPahwczfMlF+jhCF8WcWixxgFiNnnDGNX5PDN
lJ/iGKZ4n0O8uFKmeqJCbXG95gmSWDaGwmHONVI5dkg7Kd3Y1r15tnOcOqFi5Ma3Vg0saauNjyHr
goXq/ZQh+UDZ9FViRhBzbl5A/f4OQ4AtjwIhtTSHyGUQjPcDusaSnLY2YIBD3cuMbanARENCpA13
/JpE+5WI/Wcqb9yNKrmdJ1xDKYbTLOI7oazuuL/El26vIs7Aw88Wh/SeiMN/1CI11ZbUNMlZ6IV3
8qKZeKhkPrhY5r5mhj3/XRSnWkI7rD0TSjyB5D4mOxVKkW9EwFjq7djHPIZh1dXT1kcen0lr5QFP
pOn0mDz4FMFFfuK7KLExTUUJkRN/R1CGH/kl2qCx6KKIerLgNde2uYC/neiZIFZnZMGhOp1yMBCQ
Jn2lhH/0G4FCKU/sv7aiAlz+VdQuoQ42xOd8Pig0kltq84sa8vHavgflGZKXKOE417tCoguG4TK6
TNqibTmyU0MTGiBA9o46IItSPKs90bZUbuxIW63Ca08+HfpocBIAxpboq/vkqkqWB5zDODbhiU4g
k1M0nASF9aTkHXwTdP8owI98eehEGWxn+VgqT2B0d0MG3zwHEoZaak+q3IzI8qWh3eON0bw/Infk
P5hW2L3d+V72Sg1SWi+8PFvjXAY3QpGYUIIOqzqTDnrzghtTrbbpZjSyPMH7V/Pam/C0+Xi3UbEw
2qstKYYr+P5HBkMvnDuPlFzQsOzn5QmcCy1ZK+PJX5G9w155F8swrKqrQQgk2KERTMiVLdWqEKVm
c90gpDxZqDpPI8mU09sm74ToJf48Ng5WiE+Qih7yt9D6sKYFN398MjQz9snyF+sc6ZcZwI4oYbBI
9e3QuWhuyHCISawCmRGwEDY2j9RwX85OZucDy/x87rsDtAjBJLFtPSwOb3jmT3QUBpdy7H1vI7Sc
WiqoGydy/pxeDu7CgMRoGl1B2C3emvPYNWUKdE/ptOUcHQ70rGF6/JXfcupvAPUr4R/131LJyaKe
pQDXcAYFhV4qu9DmXlAec/4VjV2zo0MtTmd9YevqPdrxPPPdEOOS1VMJWZ6fH8PJnM8zg1HyLfbx
nZxCHs6QfqP8SrKQJIIkDLM+azXjGyE1qW4uVxSgavg2zQpi8x4aovxbP9sG2VhS9bOy45NtH9tK
pSd6B6BVDZVuDqLRb2HkQc6xjxKOaNHvLm8NTNMVQECvNcEp3/jAsbGjoIepLjjmzVRmCuaJuxHJ
Hvr1B5z0DDXRyFeHV+C+aRA7U8uoaMFet+zP3XYyARC3Q3VnXQxa9STi+pm/ztDZfVbBOMjaLEez
syGY6kAjQwWMOJpi4mjgu3Vqti8r268aPV4SeanCryy7Ku3YcKa2a36Da7C02lBGGQJXA1vMLAik
MERj7Ly1PH0fXHF0fuPblrVoK7mGzO2KIa+NcZDddI0DGGnQdVa2sBCp0ekpuo/8I6Bhu+W9owL1
KrHxd1NkDiy2+N5hUUchbfofY8NduZM7QqAS9JlKkqzmxDuCp34IoghkOePF8NOM0JT3rXZ38E0N
NUzarwar3DYW8LMwioEAcX7erJffnXTH4NE5RLKIVthxoCDVKCfZJbyc887Q3P2DdCHoET33tqYv
osLyTPOy7KARY9Hq9eCpVhJgStTyBT1fQ33eJBz5NYI4xB6RhbJvIL2QGUnCYDuTGU89lGqR46Ls
WU/sm5+1kzS2Hk6AEh3Pcufy1LE9DY19Y4ZlEaYKT+nHw+ZRdORs5vxImHFUC5Jq294HnYstUAgz
uz2y+0mV4+cdCwRI90BBQiiZX3t/Hq2FNZFJGxVprDRGnv4kYANRK8NAp0SJM3+G0/+PFTOSvEUq
+7+a+U7Mqoe8hYLo2DQ8HkxjuNWclsaHqeSWspmSUNm4zNp7mRjOLZ/+zbLXWz9eBE7uIS3WG7Of
d64/utqSOYABXhPqhV2Jd5fMspNfmAQkgO9NBVOqldim8mtK98iVNdrSu3e9pvyKFD9H/w2CaFXS
4b7XZYlCKu9W8s84OZQzsTwgEc9YWp7lii7zTVnA3PVcZBR/QwaGfrT3Ge7snyUpNm/v0Gx6oM1K
GJB45w0AKiqy6O95AwdSyrCaaGha4RRa2ejDVhDr+Y7PcjgFIFEK5tu+Wkz0AQyFfPzgN1HEVoPB
gRYSTElnUtTu/TrUv4TTis5l9YPHgIMAgIoNoQ0D6pylsn5fMUaAaNOphKEcykBnRgLnQ3mruk/z
sc52Cj9lElIRD3meG0Fk5RYo65bM4CqrD1fq23CRW7nKmxbpDPucRfsfIoC/WrQi9hLCiX8y005V
sp0U+uOF/rgkTwD4/DnqzzpS/BIAEBtf4PQd5BwWkUgUeTe/98T2qc6dXzd61ioK+Q165KLMPpW+
/n+npyMp8fBA6erTVom0/RL9W04TBiVNSV+Kn7SwpFtAr2DglTOvegUTJ1Rkv0rONHgwS87HAj2D
CWmd76+bCY2MvSPl/YW2wXkskg/ZosSN68t5TiM9ZTE9DdgbotdQDpWo6KyqLowWcvql/4glfsu1
wehjlOyhHfgtaRAdr+tJIeuYxW7YVNMnDC2N5vEfvYXZ3M5dZlPVZeqWOEQ+HHqLbmusePXR3+Wy
In2Yp2IIJ1suGPc8twFqtAQLy8/WcZp3IAPnUl406aPcUHW9Mux+hm7sHciLD6n428exo8PgSm+I
p/H1i2P/CqZ0Z92X4DZau6bjy7Iyxc8p/zsnwOXuB/x6ZnHdD1qA4yJL/wEqAyJmsCOuRJfd5CRy
/x0PPoCWT09mTXU5RdJyEWrEkbUjMKm1Aqmkob4kHXTWO6voeRXTNd/LZS3Yp95UsTBN1kpLCjW0
cN7F6ngBc5gkqVpWCPE4n3bR3ArCaQMFhJqHngk0Jqan1/V1Gv/9QUklrY+oVgZlnGbjTzfVI7mj
Ff95uSfbMa6C8QJbsf4Bt1WaGAA89ZI+9HtbqsDOgtnMx2aoCVXjFvj8p2wYD8I3kgan+V8dynvT
zIkti3s4Ryl0g21owy4COgC5fLLA2fiyu61UIBxRZcpYJTkK+OSob/oErZaed4wqhgpQQXC66Qb2
31nvdlFGtyBiRqTR9f5mOSoqblDttWKQGw9srKRSnxx00Eb7ZWl3zxU8El5PUZJi08vYF/cqc4w/
InwnBB8Fpqr84NXwKOxtJa4nFfUQpcnY9sW41vMuU5f5H69XtLemk6mGxrWxt6Cio6qLd9BtlqAd
j0nWsa6SzOlxWpNW1fSrQYMffDsoyp93KoJISOtKOL5glv8Vfkm9RcoPq9mRi4XPysmL4vLggCKU
P4s5FzLrB+Dgt0xXJhR7VR9LD0iC9xn4DeOFo/jAThnKbqd/wS4uNJvWNZ4ziITowhuSc0Qv8kwK
bAQ/TG7Gb2MmgA2L+GezDXizcCwXyf0feRT7nGKsG5StgGkz64EeSOqEYIpM0SUKz3y5t3qYua8y
jVxwFNwdD3IHHu3o/ruAlludvQtm78/WgpJRwqu8+J/JopYelwXeiVohkcM5eX8uLWuFZufSos7+
vmdjm4GO5LznQjz39jAcesAKZYtB1Yz0ZPiRyl58RAZ2TQ2+fB5Jdy4ld3deX0yPCo4ntBr7yX/L
G7TKtZXOqKlcZpw9jeG3u2NRYl3Fep8kVyHS0d14nxk3ntmLKPdezllz4vP8NaEV37k6K0j6euF7
1AXKf2/UUBVHbrcW/6LwEs15KyulyBYg7EeL4DK3d5mFxrCjiX83lKAIAqaOGvpk0J1yRO+lOwI5
gBk/msinY9xdOoc2CaGXera8TkP0bna8/DNfamW5KNcEUU7T/42PlhjE4ONtcqSBAv3SW3zKGAra
cm5x5NoLjmgG9cXMTmrDLqwSoV9CGCDy8abYjnIVdBD6G+RrV8DOnpxz398ddFs0wSjkCZ+nNfz0
gGMddaZBfTqmOOZVOSL8mIbhVBwUN8x7jDuapXPi68GUlGGPfRl5s0GhYYqqVa3TTNpO3VYdOZqj
28DnFBvD5qiypShnSednshG71GAsTkiKe9TyBLjIfRRl8ggGSpeh+XSRiWxswZIBhfhnHT+fWyzV
yuJX959dOJaW+rBmvGDR0ne701aDhR48+FT2tMLxu4mbaj3NYwd+e0iFCz57LzNlBZZDL0FEuVga
pK7i2CpoBtWKAaZZ9akWfwu4/raM+QNgPIR9x+0f4/uR3MCssoEqzTkIJsfFH5DlGV5asMTqHGk6
kEqYHf/91myzn1S7AUAM7/80ccsk3Yx3Qh/kpnbUrHwHZjt96qKNpEgxwOX73KBWijQ1JfjLsRGL
t9hKvJgmXmjfx9NSD1PkkK68t4ZY0T1H19D0N/pe+y6bzZWKAiAIh2ewZS0Stjq0d2rGKMui7z+z
IUaTDZBTzcSUfMkc1iv7PjRTAXTb8yC3gasQV4YkKqfpw5MKHi7axryU2v5js9vnP012L2RYgKue
jXretoQystR5JUSZ31dGf8egM+MwoIoMtUOcxOy+XQV4khSE/S5Jn5e3rFmSqBysy5nQ9/OdUL0D
LtoSNRPfyW4wLjQsD9nPDMmoTKcUeDL9U61DuRDT2rabptUJ8t/r0gpt4HJeXKQS1Akzvj4kZr/d
ccUNzNIrHUGONHwjA6TUl5GXd2yHu282AbBmSsO4EfydmqymjUyFaK9S29yQBRIOsc6I5QPNsW2M
yAaeMUewykNxLZBoeKUUl6LpAfIVs/a1tJFvbSBK5dYY6xPoH0l21BJvbjf0ZwXCssE0ukl+0Ln8
aI6MlNJggf4rRNJUBmAdxWe+q+iZo/gkBEBl0eXrIvFT1F/KJjolpqWBTc6JJ9zLKKHj572EdZOh
jmzyyfuIbyUjnpiRJ+xRhBpFU3f6Up3/8tTCLzEBayFmUhS+k0d1B0/ChnKK6aCckKJsh26lX/uC
w3ZqKZRKbudotvtVfGgiXS6fWiPk7KL3BODWXMQho+WXuoci9EfOLfglALyO1p0R5acqi+ySqk1W
9Ia6V892T5EgV4YGjpc677k1azw63tz9pkNAmhXZF1D0Osmjls3x8wAA9gt6IIeyYwmNVZCudPGG
TxGIybtetdNPRE9ONxeWjaYtJfn8+wGUWHsnXU4+Ajh1Plw5VRyk+X2engFjlcWYWbL5nXiUnjJV
hb0+AIHjtyXomZx0RRvutks9earfUSZQ6P3wDY5wkudtF6v/ke3EirdBJjbsNuYeDbaA+yom0hfh
0cQIGrC2335GfNdXxuCnulUzOqIOAuv2NwSXr3ZJFTVApYbcGEsMGndOOpbThcaVwCNVxl8qTJoY
E0iK7TnNXaM6j03BMKezXiok2cSlUAkln7c/y+4u9wNTXiJXZM54Rh2aN64oLsx9b/EY9Tgapi27
QDJxuyQwaQCnfEfYmeom4+ziR2PyqLjOjfWQDJDX0q0qjJkO1kasLaes0NzI7++18sX7ocmQ2mP6
aJALMtCR3NQXFAV7xcFuSuXifESGGkeH6HXgEPojLfPot/l6qPzOvzTKOaYggYc5aZrgU6tJ8M/C
FHWSoOwhwNw5L2G12Id2i0kNcemguCiq7kVfFgw2Fp+VBlJ+h1r74IkuYsgiVq5bj0tDUiXjpGiI
xezFgqkKxSz7yZGO2Lrg/QscU3YBJtA9v/7lDsgAhBk081Z7ebxGE6PANKGW3IlGr9sk4oQkYZ/g
+j1LsZ1QQtaAo5/3HgHYUPAcRqbaw3Fb7UGVhpnRmDZRRIC8pAvEacz24+Btj7pOOYvXyYCxOlk2
TU/dFQghGGR88AZJBhDwNRN6mJ9cPzKKpfdNOMfOh+tvTzbsGZoayYFQC7s/Nyri/WDU3KAzm4V1
mw5xf3JBueYJLWNCoXFhCBSdzXMA+kAhx4nY4DSIoOBp9YfTM8FvBfFbz6zakKpGCB+lPewmwuLU
g2kdryBKOHEZC+sbdUL0BxyUuCcEaT91cRySpM7++eHrMt4SNL6DqOY+uTY96bXEcq0pc9ynVJGG
CaCx+rLcrvu4As59ypgICNxU4BmYQ3GSu25CdbZ9YibxWnbBXVdpxYkOIwrbL5hkoBinfInL2a2s
QviQ5QZ+pQEOon1oej+o/OpqXdCG+cP93ii1w0GyZHIUqcMnFsqlwddkXg8nQhgFP8nIF8cVm0pv
XJ+JPJQ6+3FC9EqZY/1UA14c5G0bulWSfVwDkhAl4AWm/ryj39Wipc2rKA+nLSmqMofbTB8jq/Sw
l6bVW6PHk6qod6hvK5jD/Z14KTN7RBU39xlxZJ/cMUBFksWS8cuCdU3QpoIM4QiIqkDOBHhM7zy/
PS6m3c1KhASKOQHC3sUsVyOKLoXAIELtPunjSP0Tkpvo1xTx8x4EMxi2myiKHrWBhZ4Eb3H+Qo+u
hatyQCwUKsBDfWaHI1CA3zRWcZ/frxp5lBE+lDd9ggYr0df8FyWbS3JmuBW34iCPKEq+z6Zv0XVD
t09qgJLi1Y3X9DnOogUWTCWWznhq8svWy7s5e4ylubrm8BJU7KMuiCIF0HAitcA8ucF+cB32VZUh
MsyWwYV5kkmpGOPn+x2m48T3MPe9A+X57hK8iXvV2DDf0y171y4+mdmLfDYJ++OYYidgDYhUJ5n/
z7u7SLfQ0BHlHR7RZeOZTBIUuuJpY4ZJl6k8ZAu/ZNLonrNz5O10QvvPmfDe8QzSU1zaF8os4gjs
5seZnPIN+tEGoC5P9bL7nUpu4/YCFtgLT2MaUL4E8o0SRBsDlOxYj0NvStOdQcrFImLQvVDjM0aC
6kFgDTsuD9bl2W9ONcO7KzTPNECGu6OzfZ22izch+jXFXATnHepSN8dmquxiHfmVgX2zNmiTokV5
/UXJrbqbE8LiDiflV0jfmgFhPzyglwcCtiDHgjuXD/OXLD8tynWsHEvJGKRd6pfbX5DpxF6ilLrR
I+pBrPFskuK66hXdvEA9bdiAjdKe/41s7TJFyZcIE26zGx0hFHUUvUd+lYCxP388+kN1HStoIKBo
a7+HCJzwsU/A2MafFWlbFscr6I5r6ePduUna2/eB88NPH4RmyO+SMYZUbFRauJTYvhQqqNw0y5GP
ZljyVm//eg9QMBxKo8bh+gXi7t3JAIHXrz920gFRVKYLP1aa8/gzYB86BdyiyfG6Inr2sDF1NeII
JWHdGs5DnkX9pPWzov3AMbqZgvpOMRDUlkwNSYTqqrO5GLGYt2uoLgZAAp15t79foc5sxx+k/92c
dsnS+jyGRIWbwlYHLphIbbAhqDjwvLI+p/osmgQl5qb+cIaK08ipYCgWZcm/2ufI5FQiCdEraAf+
kBj50ap4O60hJEBDlBl4PrxlEmTn8kMZfRYtOx3TloPQ4yHADL8o3MyTsbKeUwsknhJOYWEP3YgW
Uxa6qndhxgUHQvZQT/N1A7XB+AZgPSe6fOJPEfGFyestaULuccj1M3zMzfw25ddOkwUx8XZUJa1k
zXUMJxRmM8kM1c9VxcyOogcx91boB+C4tG18sHGlxSQjAvqwEr52ByspT6/4vo9BFpuaxD65iuD2
Kh88xqVcgFbbQomrlOeijdXzkWRbKoQhup6xL5qTtUnJbn+4cKJP45+BReJK3Etmt3K/dOVNdOn3
c7cFS2yF8S9M0IRa33DAPqRiP+E86FCgu/IcHqV1fELuFjAG9j+uyowUTgypPj4U9XX0LDQtOXza
yFFdE+fnFxs3eD3E1YMgRCZx0a6UagCr7sqMchoHWws10lZtzdGDS0irVEIh4xJqBdJ+OC+m0Nib
KjHPsus0UwEHxOt9JmMBNforbJ6zKHQCZQP+0/aGTIYiGfyBT9K7LmhZy8KZ4LEgBjsTgdYuNX38
LXPv8CyQ4D37vZNL+CZlBw2qJ1l/Q2M9JxfT8hbIcSO1worlylxjPXSMBKNHXJIL78abW7twoV5N
k+VQEjRGEKPCzlkA+rWJlNkFVWw3gwJhVoW+M22k5RcvBmRQs2NjcUItGVDYYZzy2UKjSoKOxB8+
2GaGYwuT8SuCdb34ihbMEPs+ogW6qfvL07yI7JyqXhV+dg9D8UXsFcpjPS/d2VNZcJ3AP2pz2djn
2ktaWFAoOVRaOyff1b7vejAPD/uZA/OfTl3jN/KAjB/ai+wP98zzgrSqLEynkmaoO/I3ZJkXb4dj
rtQzkPX/pJ7/edRDadNC8W986d8HLGq81YYzfs97UptOb+bdhPIm9CryzG4a9Mzn7DbP+bNHJObM
owvddTEBVV+82W8k5X7088HrTN4zTdl7DoF99qATDlzr6VOsY4hKQaEc+odw7dO8QUhgFH3gbeuB
1yNtRBFPqMXruA9r+RvkdkfW7nT8kkrlK5NiAuuOYMNSr8Y7vQEHYRiZog0bmDZy71iY6ZWVy87v
CrNE3u+gYWIHZPV8fzYZQK17bTJeZk+lzvbXJKbRHHXOkzdZSti4Td2dPPbVKyGRtAzUZvQFnq1V
2quVnHqr6EZI6zJLX5lMIiggtbMtmPh7WjBIJLjq/1CLQmmJa15vCNmVVnTm0/maZCJBIWjZF6db
wGsxsOl1XvGdNt6gLy7Gck5vtKQbJ1RreTU3ZYOHPLrfbGE8LQTu1aXo+l+OFXDSyO3saHdf4cff
EGrjSzSPLeNSHCv3tDYIIyVwxQStIr0eyaSZJecfUm2nKKNHDIv75a1kbR5+VmOr7rZDejYQ2d1U
dikg50GpqLkgKK1FiCuw46j9lv1Fb3qgT2n5LVTRPABr/An+xvsiYeGHaVR1huih3X7tuCXjnUaJ
jNVLs8V0zsCkgxEcZ0ctNp2i7oI0S88vLwEvp2/Iwr6ppdmAb7tXE1RMm7F2Eb30Kr5qwPvI+eem
k6NcDvXN8cL5ggBWitEsc/uyw+ZAKxkVB+ZK0NDlsTF2j4uKqSf7luwJMcxrofiE4xFu0MVdpnnW
Ed+XQh2nayWgEAhbvGQiH0H0mcaAxefROApZwCoaJlq93v1znecvgVb67opgMgEZaDnZmx2MdVnN
JTY0tx3VHSupLnfaH9klsG0Ta1kEGUyqQaioRiG7m2RhfXwyWeQzeeBA0q37fia4Fx5jmCicO/56
dxvOoLl5ufz/rsOJf0hAvIB+pAaSL4/idRDN7kN1SfC/7X1+Hr4uU0Zk/r3ic3Ab9DV3bH+u7ezg
6rHt33XYX5LHd8wfYiobipgVxsWoBXOpLfn4CzVDUSp5yxjCl28USTJVtRWSjImb6+XyrCWVEvWm
pzVr1ZJw+KFvXynPYTBA0hRfvpw2je64wAyBINnac2dbUNtsxSOolaQfaUHGjUq6Y7F8ViN7Jy15
GC34YE5m56CVjlZYxJRUlFHl70TT6o/mr44BUVw4dzt//MxECxaPUFhfX0QvxWrgSLz3q5ELcVtl
LBECkjaKbFxQ9G7LID/BGDFLOXngY0MbqeA42ARxtje/qmshQE8K8SjbGxg3EiFFU8MZKBUhblrV
EWiajDN09WVhD1jCDlKCr41J5K97xyxVclD8kuneCNnuDY02OdCC5aqouyRP9tAza5Z527yKjo9v
S83HEaFwJ08bLqoatdLqALm59I5w3jm30F3MWDsBKc3lKXyDNEfZ5JbDYMNT56a1v+5PgzDor3p4
KhEqzu3j1N++Q7aDCDx50cmCR+w21sqP7ktUx3OgU35NVCV2qjq24MyWcUTSI6A1M726csGd4ib0
pGKgbt4s2L30a6sWaLrtcIIRjlw/bsYhtMW6bGRhn24yMUHPdWGlEGXQxsI8/Oc9UMvivBqpc48e
TXWq/45HLrRqTfgQwyPcFBtmWRw9EaS62wzC0jNISCubqcJS//QtKnisSIv7Zs0wcy5QRW/E4tMl
P69diMpEPBL6HPgQ9LCWw+QtwRnzGqhbwRV3YhP1h18dnWAtQTBgdn4c4geRxAB7j1iMryQV3oNN
XAorrwk3MMzLWamHsJzmj/AIhPudVJeQnJsFsAuaEbTFZxrmV+ywzdKrgoKGPcibbPEfCMpnyDyt
0+NEJJRw7aLtQjNQP9Yzp3Jni0dD8JPb2cmj1vhhzc18tyxABisR/UdX8NK1EBOFD+cHHC0vcwm5
/myhZprMPBAymLA/rbOKxXKNrGPqfFZg9jUFMtYep65WWBKrDjf+5kt+ZsNQ98ug2ywNY+rXDMA2
AyBmzX3isz6rWZfh5Smmvuv8vk2a0i8zwKQwNkevULDApy2N+j/Ecq7jqztDr5U9ouGDMslZYQBt
T3UCmNE4IvyWUKxICSO5p3eoWxtIaL5Q7gA120nEZZEZmhpZb5FDsXRNKEsmVkMPCncHudHriNVd
PKK+jZvbNt0BSnnApDAffOQCAT/Epbjj6tBWpzzfucYik+8Osr0S+Bv52i4wWzypmWZsl1ykxRra
hCEMxfgf/vADvu9cMQC+9/L9ofwdi1O/klJh5uPf/nlRkPziSq/oGNJhTUNKofkEQsxdg8gob3Zq
tue+4lSd3tvfOFn/FjaWZWK+bGOoTNeaoC4hUSOjSIlLtAEqJcWfVvQLoo1vU14jl7Hv4+VTQbot
z4rJxFV0lgsSLkM7huqLM2Jb9WT/fI9eLLpTKZEW1d+roDDw1TfMFacZXX6vcu93Sqxm945xLmVj
qIRl+2bvTKJPYtY7JbNf5vObTNT+wJhsnoeXDn/hmzTTyDUlTgb6ejOIaV2X/1iT4VgfZbq6fdnN
0GzLC0nuDUn/g7z0a+7iy2Y1+SFJcE66jp2UxZqXpQUKxX83u/ZCyySg7D5scpRsHBZMGiQrxELP
oAzWU2uFJfXUAYFkcVSUYawzkoRdxEHgtB9Fs5kS9yPJ15F4S/cEXFvrfCBEOVeIx2l6+LFMSs40
hyR7dkZv0sVn1F7hBvcua4687nVt0+2RqHWsuUhwEg3ay+qH9FwFcZHXToAd49btgrHqmNhZx5o3
kruFlq09HSeq2Zs+3WF6TGlJhvww3KXPRosRDCnLmMPIrGMnzLilFwonB0b1dIAPtBGZhfHSE07N
GIS5TqhzS7JikPfl/1yhsLUQQy9a0jxdeAVhzr7i9os56D6zRqs8rq6IxDNxIe9aOWT513UMEbRR
oCt9G1ybdKn/p0n1x/I7pmGGISjLQ/LWzh2vO6B6G4wojdAhhOLU2aNBfjoyhBEBFT372j5S8COh
IolRlCqfpRhlxTOvn39s2xbjvywGoYE6uX6OsXRHHm4TpxbIktHM5VtiFoYnG1DuXgal9jS+JRRd
TvyRebRVctLUB1Xj/elBo5uWIAPzlU80TBQ7m6pdnGaYII8qsQzKbVS5Q7yTuQbq5ZHFW2DavejY
Hhzwq815Vfx+4ti4viA1h98wmatqwMnaqn38TAMPnqapHkidUTKyOZDMsL4VFPtTwDUoE5/A489A
tgN+//nKCAy3+w3VXJ6h8jEuCdnejaemQY+q8yNeWq2/f4TFO6NgwbviMHgW0PBfLZWQGekruYdR
hVLEzJaUc3nIMoOzWtMAWC5jjgSGGnHMLYw9PDfgKhGufcX0+Y8q9blPncThkS40k1wEm6mxg5Cv
rlBmlfqWnZZkDUjxM3ujfs1zNjdXAGUQLZiBO+fF+PC/M393SBa6XTWKgcgOPahdJc1JteNtVTdE
eSZmzpmS0v8kouQWd9AilVNoItJSQCTC9QwOuHE1nCnmbTNKibUM8WdmLgPGA+MjtgAzUvucFC0l
tLpS9EGZqGTyZ64yO0VgGyp/k43CZCOWbTTJ//Z1BSxd/2eelsti+b1Sab+K5MgWk74mgZNTnyR0
a0nUTeQt+cFDQ0oK2kPFo3M6dOfPTJCurNVWKl+7A3fJRZ09hgOExNX7NlDdI86RNZzjTey73PaC
Z7nK1wf4F5EZLXwkXG+f1nOLUdWdnYEzQxUFRjQ39A6CEgEbfyZHJU1Y3TLZeg1T+bS6+7cLdI3J
dzneoaN/Wlnb6VXRyydH5K9UmfnvA5PhM3tDdqk27BolHevHPXCX5qprnkReAHP+nvEKOOqa7iAZ
udX4e5jqv8iBDbYZrEFb2O/OXjP+UeGFHKwOAR4M+XeVHcpvZX9rdpp78T17Y2UYMZIF54n1AonF
M0B4EedBWsJetKTl0ZhN/45GoHQDrsYZgsl69Xbo6QywJtt0KJxyIqSUPYVdA5znWP/YSTpmHlMl
6nu9chS5aSTK4XhxbRNPDM1W/HQ4gg4a2YyWSCgQV8fCGna8gKqXlIAsjx03sacLIF8zVJMdkzO7
rZaT8izcFiJQyiZJcTPAAiQ7nAYeRGXN4tA28OVdhnBMvKkuJOAiot+xb1voWphLBXZLhcFydozT
QzukV6cDrMbNca3Bki9E4Vhk6kBoaQ3LS3tbBrsfYNaltjWVUu6c/pEzXy8oKtRi9Lu3GGGLYq/R
HYrOHjTdhV66ScFd1FeffA5GObP07EqUgLayJsQpJZU6LCzcTAaBX7k7IKooFRlAgdt82tp26gWr
cDKzcz9oMZAmpGEuvYLAREB+SpMrgQTkdIgOuKUxTw0ZIOhwbF4aMYqgu6bZ4lGaoMPS8SrXmrDO
ynU3xEDJdBCm2TbMQihp0e2oPL2sA1wDFmVp9WgHANx6n9bFMRlp3rpa4FpN3OxbEGzvr/2slmRQ
9kNkJikUcoJmrexT2LIVmZ1Qzu11shWezgPgwT30sdBWXnx6T+mK9kgDRa3l9P+Q1vLsBjP09/Z9
D+u5QHQHJ2dBEqlulpylbO0t/K/krZs4gDOqMXmB4n/hZwGXmrAe/JTPzqkjSXiYm8kJDz3XAX2W
dQ4qiQD8dv4+eaXdfZpo/wDatAjdWTDyG+hX/ZIhMX+aV9eGkcrUxeG6RhTQ/wEVHIuQEzYybwcW
m4k9Dtijh0+ZowfthhW0Nef/PSKztxAJm6/sfsPTwhcyl0EhnTQFIz29/SsVbcFTbEv9Vb+FIhtL
sGTivAKrjy+8rMA7RgFBdXpSstP8N34ryVhJP0+/nEpq41CQ2UwdS9dfoGZtwd8m+658SKYTktaz
KimiXlp16hsEd+cW53edBTKpQbKZo8amF+OOuAtP22ns1yj6EcTguntzcxsFC5zRb6SryXgB6hRa
T+nxbNbB0O0XOmcF43hvaquFWmlwdIKKU3IAQ+Z3Lj5h68ASbOcNrTIosPVFRhOWgEeNrl2iqeC4
Iz8KL1VGYnBCCLCKjOIJ0576v8QfHXXghmeG2Q6p6o0inl3EZCtUJY8OSnNPfBf9JuuBHlDMCP98
ck7Ohfp49YxvSa7Vwoo7aKmbm1VSst053ycaWIE6LJyWe/xgj/uRRKijN3xlPe+/uyejRmwjTfgZ
zkQcfVwJ9jijNqhoTUudMlaaVrRzW19VpWsPdNxaFPzm+H+VtSFIzHb1VIyv4GdIPPsG+IC3S1rX
x4PFqQGLSXhZnSYkc3Z5vBz9BqKPRybOKSpa1ZA8U1DoHfp/jE3q2PK5hUlkYHQy74+KShJoZVke
LnSZeljIzZcaV9CqeUWLQAGeNIm2U/ka65T3ONLnfmP3OpfjGAIc/und+vqKndFoHQkonwR6LWip
PghnVKkE4PMFi8tG+5J8Sc6cpXEPWYDx3WTebDdAn5iaCCjoKg1jFlReX91BCs6FC8vvl/DaDNwX
MSyjDIMj8Gvpj4eGD4m2RMytZ+qfLF0au/RtnnSga/5MCXd9PBS/ncOiqgvsq0F64TVyQqBBIO5x
nXH3o3ZAu28IjFM4r25A5KAQsIXZxNxFN+Qs4ArBI41nk3W01ERDx4/VexiZpqPcj6N3B3BXimOk
DBIVd/u+uY65rs0y9HdNlzZsFQNv84Pde6pIS/NMyWMy5HCuSl4dvl3Nkr8gmeRMntpo+WbuaAuR
WJQxrHrrPLsE93KJBFTYIcolmu3wHcpOxzOBJxrpF8Uae4GYdlcG7PIbWHVXDopvJi7zFY8U64k7
H3OspVBZMCGXzmhxk6HnmmwS7/xAYRCYHmp8JfQd2zaRQjJdqmNJCrAzCpVKhV3Af2jvFjQytzWS
gowJnjCMFwR6nFD7DRMdNvCuXrCvKk5mrixyFzmGVFCF8ceE7coIZOVbbRpmnzPv3RfvbZ/DTSJH
jbnnLSzsHBGuixx2QZWdTf5LTeSFoBpxrob6U9GMzTbJJA5DJNALeOi8qjTvZAYhbtjw4YesaaHx
Q1ELFhO7AQZ9jJsIA3+gygh4OSc3ULXEMz2mhYRs5dpFU4bhrkHD/YNKqvRFKJSd7t8RgjVTeco6
6gmk8qft4w0JK0KcU/i60nX60EJXddvP65ZYdAentZ1XBmyqIFNvlSNYHTWlSKkU5m0ilUXzk4gv
PyFq3sxoZ6TT63EJVKyN8VBPdiDGTU5d1p94UVj7NJczNPuFbLJZmo/5AFpjegGLofEaRuGBNoYx
3UTCE0Mb4OdJjem/IjgWjmZk7B/4bdd6Mdc6MQuyJBXzSaJXmeE8qacGtCpCJ3X3GyRJYvp3ip0q
PjedmVinuDERA0CQPwYLQBYF0SrZgzM+ZgRBgfFlTGXM0H+Aa4oBjfpbH1cxVmH0T/LWWrip8/VC
8Bn3Y9vPCbVcX5CIJlXZlQKk4RPJfKKWMVzgfSotAfSILNP3789PvumjwNd5KsUCcCk2oUq1LADm
y2ei6taFURTQtXN+IG6I5wiGVi0g4k0OlhIKxzPuHKvOCybSBThSFCQHgM3DO9jZPBQnW3FRINeg
f2RQHa2aW2QSmGiDpOOmD53pvK9FWS3uq9xYkRxlB1VM/Dc+V6TEPdSdsT0nQRnOc59au0JMcnle
y/Wrhglz7oslAp5Ru2dKB6mqDSqhVPLC1ROmB9O9YuyNELNWT1K5FUdpMg1191Qktnx4bOydCDXK
oksPgxBLbmV0Z90KHgL8Xkx2OuQ3APSsWy648TlQqjhrBUZ2+tub5zUBq8li47beVmmHUBiTvxey
OV4tzYPC9DSBI+80XjX/YROvhwAmO9UEyLnse3KA8HpH3ngWzhW9/+VNYWz16pY7rqLoSwmOAMPL
4w6n93+OIB4OyBGegEi+LjXThHkmH/AgYs5BFpVjPtYpGWyUebEJWfc4+1jVEMXD2WJS7/Uo9LJQ
t7zzM636uW40xqpbYG7g8POU3rgxklKjxteFKmTRytfXfKKbqFA5sVgM6lgDwmR6QQDVCFrOF3an
gjAuyb4FEohtuSRFV7Sbll6CBhmamKhPFgpyQOLsZmMTEnJWixCT6Q+zc+3MJJC26XHzzlRlaxGD
0GwR95JMG3xrcSrxz9zitRyxba+qJ/uagoDz6zw68LWmQtjkQidkVvYjBb5jA2XuWPStqXSrkjFP
pUoBtSsa7dauZl3Zf4eclf+bI6zxiLOQdWknP70SIoUia8Aeo2RoLOMlxhP3szRg723DdajO3uef
ut+aCcYOfYne/lJTY/KrOMEx9KK4MxW35CB/RpdIFfnrwmsvwVEwL0ShzP4r0JljZVt++VQjwUl9
OVhPAIXkvYTCumsx87KWoLxyqHvONKsKqSiMW2D2FtoR6AwV0ohasevZ5fFv/1e71q8c24jZLQJy
IDprvq1R4CM4OgIioppWSMJ3SVf4SW6KEpwAYvZ22hpUEM2gmsw4euCIJRctGDw+G9WgPrLT5lgp
TvILK+WVYIlvJ0+Y7NPO3S/SbPR+r4sN0g96+hkx82Thu7ym1tN1VRfklKg/sDG/gySRY4b0lfeF
Zqm4sBSs0MC+xnEXq6idTdv4V9FDwy9zvPDexGI5PzkpyIwUVv4N4FCA19jGZRaoxm/+38NVcENA
vKeeluVwr6WMHckSb8IBMX6mXIFTFNBDSB4qVhizCa8FjrSlOM28cJ/mjQM9nFfN/0c+FzZ56+Uz
tCK2IXzBWO3HUI9kSVK0VCqEegjlSIziFWMZKu9DraE1a2u0nFx3ajJMTCmBWJqlBnytH/mKnzdf
CCIZP61Sj41tM9SL4Cr2/OXQbGhjl6D9+viLobS87wgk9NXy+oDUjXa0f5mKhv0vfEx2KCrtQtdZ
UDTdyPB4xx99DUeua3Qwsd14x/9VZeoqOUY3vkX143iDj4priFAv+5KdVUYkY55CI9+6APnffmb2
Qn85LmXMOHSHUyiiij6Ss577P1arJCDFANonBOYis7vWWs5mq5DwHsPbZB+vmA5g6rUjyt/NMVIe
S506AzIRCEgKZSrdJbnSV4VPqyOfn0leNeFd8mvsMSqu+9G3giqX3HhqgIgeZPjMvNhZQnHaJWpB
4LhwkpXf7maCt5AA8/8TD0hBiGjXENHIOE8EUNxPDt9iuy/pEXnzcLdgJQjE7zwhc02x0ap4N5jQ
Tf7IGxNBG4Sc0PBsULil70G5u/IvYc2IDZ7B2ZD5OwY3fjLAzBpmsVW+rn16gGHtH/U/3aN1J4yE
ujSh+fg/UH2Ca/JwIeABwbN8a+Mqicqs2Ucg/BjDyl4YfK6CPasMMRY/vSvbfJKHZom/o4v/u5o5
/SD3F4Xby0XqEHkRhCAcI+hSYFrE5sZSPyW+gFMDGTf6fR04/KYsxmt7tFEiKfOVbIJKuM10HXe/
CShCjxLyKMrW9I9fxE4BPk9ZrgM4J7AqtST1YbN1nortvp/gHGkX5kJGRJeTydWhwvjtd9VoRBJs
snvstH2n2KGJS0vbAjcWpm8MTT8d3y54iAEDKmAjuDtbcf0JWr7LBfEEGN7+XMPsYKmeWtAAG+wW
j3QlFegFU5kvQjYmbzEBeEwMi5ngfbuHMlXg6tM+oOfrCMLO/ajdVyZsuI8RFYzVYoK1rE7vqh8v
+jOhNS45V1mwk2tYhNRbnO87g/XAoai/ZvsjGlIG6p6QTL23s6k6oKWgwDQ8jwMveELaEQSpfa9W
49AWaoh72QMsovlqys43Qra3evDBtw+KtU7zB01b79u7ukSNOLXJg4UOHOoPx3Ox26ujiEm4bqRa
i4+/XcvSR0aR8nbgRIGF3PtEYOskzZ0pZmQddkRBULPBvUzv7qvFH9Nbt/s2Q8xw4VVUmUNt23sH
Ut3d8IW6kaJcFAjGNSt9LIjKAT6xwg1ujBOqVxisgBexZ62F7RaQkyG54QuMpprHj17cVZykotGd
ilVmFPYRlTC+ffPkK0Bx6qZ3Wru+FzK+DUFgaTTca2b5pjlDPDk6Bp7ggzZ8TbthO7MSBoMVdNwb
FkoUgXbyDajtc1+aZwBy5Sd5pirKRmpYFVfLK1n4U/dMC/10qmuMSsx8Bti55weZjAf/MkWN9Tud
/XhiLGB3lt5YvQ6gAV9VFn7FLxGRIeH5IWkWf6NXHHUMcpDsARkZ0LYogsaYleVEg/Ejfcb7m4vM
5gc5TQm4RWDrA2C6M6Ufv6ccKpflZpBbY6kGo9QmitiHJy44DpfcubyXjsXl4DWQ4OIQfZLVf4Yp
eH12sBBCK1ooXqqajDjDS2uk2Dfd8EPYmFKiRcyRugrkn4xfFSSnEzORGfGBYpKZBMl2tD7Z1sr3
2yBdrQyRutxvDYpA4KTC+JvvAGzhmBTyOZtZ0GK7oSaLJ+u165SOVMLSLWIfgYgU765QzeGYuhQQ
vgxdsX5Asrtge1DSzLRgmEsAw/IiQdOT/ux5VY75RYFi1nVBOPSU9sXq6oPxhGuMQoE6ndM/2r6F
ZeZSaNBlzmnoPaya6RFPNXhz6xYhyaNEJL/PsWYXATUIpwBY3/I0NoBIHoa0SPitmSPb4yF+GpTj
Z8gvGXGUCdtPZoOQPuAgzkCBs9VXd8lU4sbQN0kgFP5owZvu7PadXL4uav5edxsP+Y5fe6vjV18T
WY5hKep0hwm1pY2sFVREjUSR6QIXobAsTuBs/AGfd3PHBWcsL8BhKFKIaD1ESzgAziIX7ScjUWk1
QU5vsB0TV8BN4lrkMrjjitFEZJ9QqaYL8fTZgsHjNzcodaAQmOvFznspE6HBe9GIdQrxDtv7vtnj
GaCHTVPNDU4po09D0oUGYw9kupZQowvxnRJGoot2cYaiweP8bQyZRrR0oVGTqGZvV5aOr4PAJAOk
NlxepOxlZVJdj+JwLK5l7E1PNVdIGJzGIropY5QaiPgZrapLAbOBN+6PjiO3Lcbv6SySpoaVoQQo
o4CyroVKPNw1pQhAQsGR5sKDDfNoYiKyoGRFma2CPR4ntLaVmOnhKyp240+YsDgLVcUS4TPmQY02
CYEJMA8hi4IGZNh48ii7LoZAxNEWyWWUu3XARzRfIAJMVzRzfeI19yuwtXVaekoVvgVqCH+JMkrt
nSX3Zd9pQa1JEiFIGshxtwX7CqwtK8laZ9XXI2CLyRIQg87HxH/BG0qserDRwfFEJr75iuQdLGEc
dGVU882AfcgVYu+HBzKzJs7PfgMYP0w8Xz2ElgAqNmh9fLFD7731N4qL/EWXfc3j01gwC5q00nt0
Wr4XNiT3aFhyyy/N6MRpZ2KW4Iw3+XVK/km8Yx1vD62RuopPTdob33i25iDdMWCj3cP5iLZzF53o
WPmr2bRMWtdVjkEoEmUKrktrUvYMEHe3uzRhytVZflkFjegwbEsl3AKNVmWO++hHWi2zUetWyb0v
oZB+or5jNZEO/S9Ga8EoXyoHOJ5YHcxlIGxMA3cZOaObfw3J5EZd5zgAXyMP1RKwoRG23yRWy7Vk
tDvzHT8d3Y1vQYJ1KV4nwwtS1abeB2fS/eY9/TpzNGgJi56RMYk+eFmaG8esksPUlOuaoRYlJL4C
xlZmbEjjbByq+KrIV/YSKoPIUpBzXVTLAPKX58YJnXyNs6jblEH0T9RouAMwip0DiKgPYVvoIRLt
eICK26QX8f79QbDXcbf0wXBTo6CR84RUqrdp3c2ys2+OPrba/sPdY0Q1UirupndAe+HYhxs3J5TP
2vwDHLTTCv3djXMUCNT9FJkaCcMNGmgpLfIIWzhGi9mg+TLtjWvfXoldtaxa30V2mrRDWglF2nj1
k3rTcbk1rxULzEXwksF4my8kLFAyTirTIlTOKbL0SD+GrhUBNVMXqyVeqibBsremHHGXZ3IOCJRa
BK7IukM+YyCk3rScDXP2Ejqb5hLx1Yk8G/95ozSe703mYbC203EGNe5ccT/nVgLWsKpeVGR8Jh+m
XSD8RHMV/8x5UYH0ZVieVjI0YasLGTAOeF0/wA6o8jpjtBOuslmwqYYHmiBeCfW5rkzBWS/Fy69b
umygZPAwz9K5680cVmaKfxNHwK5/Wp7QxCT8SCENJ0no6F/yPaZIOuVmMtB39TurLvS4GjIiirlt
70C6kBpPLnjmFFE+3tWu9P2LH91b9gqi1TIp3vrTZZp31jKaOf65A7neznQyuqXy3LqUKcYORq73
uROKE8IqhqU5J9itc9Aov+KC8xduZZZK3Yy/oagpQA4HGODTWbNCE9+AZCSUVdJU8A2m1tRiO0ol
O3yrAvwX5lPzhJ9Iq+HZMA9BLY0Pe7LH+s5DTYTJJvEDR+nVl7gUtT0qxTEwUoHAL6rYYbfmQsne
Sa8PCoP+iviaP1wDky5R8EPCNAuW64+UBWq5QqCkhL/7igIrrm4ihXEG2O2D5qwl6dfJ3QXJAfza
r6kAPZcsfW9S2L7QckcJw6fChMR232armEXsr4rO0Cq8Hp/YEUOaAsKDGe8SszhKjOhkif4b5ZI8
9khpDXqrVbZaMr5nGzI2SsdJr+e2SbRk+5LdD+p3bOWoesOQCYJwcxAKd2OA+GCSCOwix4TJVAyf
e1nSqFvkj4oEKnT6PdAE/1EQtnSt44vihBX7e8d7E7ZmlC4en6eNr8hM+RaKDhbe262ZVkHg1CSD
uFWexElQyZWyce1q8EXK+h8Bpmj8USyw9hlAulJVBfO9bT96KtQZ/HUGDP1Rx6gVrcsRoOM41XWL
Px1qVWWAnuIySfDGa5vTR8D9WtrSKLqrMIKvECn2BYpPAOjg1HLeN5buAEzd+Yk+0TM5vEKZdSk/
dXdRvogFjjDTY/n75+hkU20vEImBUkSfntwn8HXFSWZup89msRfl4sIUpr54v8SFOu+O5B8mbv3v
r8xE7ZfW9XdcPSHkHY/KIYzVnFaKLEuU8SLSyyXuqT2TPlrNAURQu4ombhOSZ3jroDGVYCPR+mRW
uSPO93mbrkVVP2Kzyww4njDEFOnfcyTsohYuOtpFlfeVrnxD/hirfgpscmZViz/MJIz8BqDA5CKZ
xV4ZoC6OlUCqkonP6yX62Ih2S237CC+KdY8pa1+iuLl1hFn0+sEgjMeAULRyZz7sBckJjoIs/qmK
RhgvCGV1FGtHrSUgytDlraQ49LP/WBsNBMMyNAmS4htR4X0/boiX6vm2i/NMPcVlCr9/7aes2sfA
hvU3WYYAPsHr5oDScljCfYj9SCCQvpHHJabmJbgyrnBjjPLKVbylAmhp3r7lY8M445Olzk/LZIkx
tTRLguQx0L1bizOT9r8JYrSgFNGJjQdLu/tV3dpmgXACeZQZrcLXPWnmbzvtPav5qWiTy2T3THj2
EiZZihdSn+QKuATQ4SEE1qYD2NMJXtKpnvNoA7l5iE2aGx9QYJcLr4Nql5nG1SR7e8owdY9949iu
RsptKPJ3XTn18SkjuEMeaQ6QJ4GogjeaDwlmVP3ozQckolOSKIFCe0DDZKQErdZ5MEbbOtmUAnmt
eprUewpcZfH3w00JTj0tT+Qw72uBrMR9jngDYUcFLYW9u7iYmmjkFdYVepAnC1zM2RQtqjuCrSrg
oVY3UFEuWsvF9Qt+mOFCSEkP5v7eZXYGCBHqqwTOyh4z5sAESl40ErxGUfoV4oWtsIU3fenPkeT2
6ESCCbh1PRYcHh44Fn5/wdH1XIf+Ag/ASRogflkDUtBRWnfozLERjS3/JLjdv83lNt0OaVSNxlTl
2Xws9d8C47joQKwI21yKPC60SRjAuHX1FVWsZZnd2MjpLMfGgDOr6BHOzn2DrZsui78EuFhUAdL0
GtsiJaNEG9e9V2X4kLNECDxQGIRKdaZ7/QDZN3XxxdjCPLfmttjC60HsxMZ04tOb3JJ6QivrNddo
uqF/ZY4DXXqKqmX4rz65d0utsgmnAYWRq7UGejlWFxwZ/CnXPbCXi7hULz6D6XfDigie6JWd1pSN
hTwBm8F8KZ1ILzQRcF1UWExAysvGdpUo7HdSa2B8YKsZpLjpIVRatP61Xe0VmZ9/tXUfrmlT8bIU
n3N6eEK3WMEOVa0xWE3/R4l0ThjkCm+ZmcH8eQxEF9vwBXHWjOqSdyiDbD+hQAAGctMLoyZVPSu+
kgUy67LmrGnBc7XfFNVk+lkqBbyB1fzF9ea8bBuW5zyCpcelYgnNSSSbS/qoPKnwVhfCxTj82UXY
WIuxiyRvm3mKG3QC4KjcB34M1C2hRrUlwgWrbmC1ScqBE1TMA4TJEjJrcXB/QFN6T32T+ccB2mOz
DulINPAWfKETvgOCeRcrUvAnxmhJq2VX2ZDe4gnsLGaTJVTmj/4xAISlJXyk9raKfKSWZCrhwU+W
Dx+Pk4aGOruItWaJ2q3PlIq2wNCWabd1igZYJSmwexAObXGxJlfVcDAIOvOTWtiAInsxfjydfR01
Htwc2dtdK+vDobs2CtNZ602U+LE8A3wmxU3zkeK2LEisP1/ceXGs6ddIBZr7blbKGZKox6O5flvW
2W37256n9+N7sBx24IVCjuQ6E1dvjTZo3x1LLaODmA3Y/gt4qwxYU/5UGhNNpJXHbZlFUI9Zfb78
ZzypjrovuHuyN3vJz8hh1mThsJts+aye/dx9sbFQyfcgMUGBE4GUhdmZ/CoaCzTwtaN440D3R2ID
FJU4r5wxiL36t9EukA6heZ9TJ/dfnN+Q+DEJylNW5NcqrP3cIQwBE/IHbHLW5l69Clf6LRnxuCid
ovQ7uvbYFCMuHcPQ4k2BBnRKNwlyjilTsnlj2UjCHCViWoe0XQXeLvuObQNeDdmZe9IGATAIz3Os
3Qfw7c7LJ+QzE7bvbBoqt/TAtWkfwO+n4LT0GQ/S/jXqzP+eyg1AZhRybMU3Kmx5cSgvbstEjF9L
WA3rfumjYric3oJqH0PpPFoSyjTR+FfKfgBj7w7mJtZFUP5Pc6kGAHUH7xi9TQNVmJ+a/BfrrKeM
RMiyG13v7rfuiHxCgPrybAgIg5Jdo9zQf897dn0bEZv6Kmo6dphlNdYiQXJUmIk9kPEDN4HpoOTt
WFnQ6iJEpE2qxZHVopJ5ci+7dyjGtc1BDr5uLk5Ig5vfIZlPTLx7ODR2NvYJ6BCvBAXOezAjIkIZ
glcUKStOxdoa1UoXWbG5le9JNexIuVMsnVv74UTWZwXtLm9722jEpIO2KXjO2DZlULvy8wE5qR/K
trpF4FIPUpIsBgRGMYf/HAxv4gkknEGaVxlaU6b3M5OhIfO1SqYAh3e7TKpSKrKbHce8UCW0Mjiz
fA2ZTc05W64N1X0KqQKW7gjo/BcVxctWSU8uXi8XFR385EqQxn6LxSXH+0KCNu0ZIBYRL0Oopagk
mqnRFqYKWi5z2nP6Gr3ns91wg1qWxscOdLYnfPuiHszO+7E0xbIFd8iR5ByTA6dS7UiymqfcE5lC
2m5dCCiysxZd1X7bfdwPIV5Hv23uiMRqnDYjFyoFTMwmeoikUC6GoKDxzoqF4TEJ0L1Fysb0Yjoq
1UZP+W256wT53jP0tqnz4tQoq0KqrLgqQwqtFdrA6rIOSd3l7xvFbm84Mh1MIHR3bENy7KTqfyjA
26GdJWGa4JKYskQDnbAdrSKp41SEKxtKNMAhFbplwCAYVQnuXu7zeqWsw/EpwyZJFWyPRbx3L8KH
7CY8r4OiQ9jTDwwkyiWpQa+kD3uRkuRv1scbaZZvLesonQn+yHfcS/VNgZSuwLJKGbQrT2mDgafV
oVEJIPpC00NTxbRpW5dEbfueID/L3tMutgFXScb0cVY7Z3gzsJL3WhloesZrGxtY7ZGCFFi3mAYj
/STCzeN3PASSaF/q6pdMCIsp3u02A6Rzea49zwKa9bVdZl+/wkjRTN0HK98Qye5bvg5RKAChqlFy
MP5b6lRbMj/meyrS3ZSvUWA8QGPa0ghH9gf0Sx4To+tWGShY023btoLV4eIJAayApCzsrtXLgP8T
ieVMK3MyaPsWHfNJhYzcto+MbmKtq97BWAkXwX5hgLLeGkKtrhZ7Gu2/hdGJL1ttjxfh6/bLxy3Z
VR9sazrfD/Wt86rl/foj0LJwqbybHb2toRnFYRVAojSadw9S04X2/h8+NXHgVRLdp9tBAMYTumcT
EwAcnczhxonf5fzEXR0WyoLr3P858Y8fuyR1rt+k2zfB5jLywTMiYiZC6cEHp//UCV3tcbXrtvGt
mK3p9q/CU54wleh4MTzkEF6iruF4wFzcIiMbq9Jzy24ImIosVTEmAcIeajwHb04yrG6FSFOn41k2
0+tfNt+fZdBSRDpVp1VdZmzBzGN39pids3vIbipyBcLC+upj759MabbiZGleyHfYRp7K0TYds4AW
1hCN+8XwnTmlcd2MDM0qyztwuzFaI8KyPX887MbI+N+ABtqR22azwRvgA9l7URJRkfFMUc4dwwaK
i+oJ340eUThEuTzj9x7zxaba09SjwbEn5atsIlGmcZs8kCgUYJofjCQuYBF63q/U6YpAUR6dg/aS
MUme7diIiNVJ9Zpkd9p3c51kUod/RvTsR4XY8MY8PvccRHWXPu4eKFgH3cwiVa3Y7b1mIhiaW9Qs
JmXVwbcT3GoTmmPUwTzDTngRVAU3vbVc0TnjT+uyWrDG+Ba/6Q27AGUYN1W8oz4ViI1FV8OWkR5L
NFzh5UMUU7xH7HHJkMtv+oB7ZhopTYlOYo7feqrtK+D6Ow7DXoJ5b9Ubur/1ajEtn6VmAsrEjOfV
6sHryDpOi29ytJfcGtRCkSBQsgtG5XB0PKrkkGVxxw+kBEZokTsl/+kxTTbaJyKMaV4N5Rxy908H
5TkqTpCPJC7nMTNFJAi2NiMVmYIXoATZ/fwIEe0sCD8oN1HsnaNQj9EQd/lxbFiUa6wwIgY+3Sul
mRUpF2E6myKGfq34ek0DYlFrK1rz97J721b2grjd8LKBK7TBb/9vZ7mlcH5tBAa2NOv+eQ9GbZba
A355EMAnKNfqrqQjUkgiaKg3MvADwOLKRfq5I0VDF5mQT0LyriGH8PW5OcpoHFNHxycZaKYbjQ+x
hC+VL3jWXVbM4I8My5cXuI5ZQ7JhIbN5JpoS945SHx4lbLjUR3ezmuMh/3Eh1iB4udzguFlUMHHQ
thsMlPmlkWvJ+VGQbmszkTURrb5emRT5fC8a1UVwoWLkY2aVyKBMCs6dMFi44tPIG5xjQD0GZnzI
ZKbepNk8Xbc0w91PMajI3ESgBBdFfH2ug7BTu2kzOrQZ02M0Kkav1oMtmHGCr6K3CTn/WrasTYbV
wOLSFnFiDfBiSzAEfZwimrIf1zlIprghbW4BjiZPEw0iuhIt8ILd1vhP9E5AJqi6SFgUczqJCEEV
WK2pD9iBf6Ev4gQPDIrXdiWN2DVtldTyhzcpeah1plSrQKmcbXFTwt4HPpdSLLqF6GVEnBY5DtU2
hAxpVIthPBywX5ySm3kMZ6Rp+O7gysd7fVL4kWAsMz338l5VuvqT4zrrrK2xd8ouO3j3AFwzHG+z
juR4PmW6LpNptKE7Qa6fJvFu5Txmao5Q4MCc/+fE3uU+yyMeYT59L/+UEzlqlVVWbYWW6wIQBhZ0
bhqyIRfIgCmE5xwZ3LhuTDxVpcANO9pyVchGvXk7ZvY8btH5YAEg165AWg/W5JlRqybPnpzEd/pE
w8uqAcvqRSd2fAJGyAAcxMvraT3pgspzfzX7KNrsfHbd2nhOjSS12CRlLhv7C7YtYarD2XJXWo1E
e0Kxgj+fR0ZpJP0MpL9IyW3qZcFaq1MRNLly7xUsk/4nz56jnIkfjoGOkX/gygXm29jrRjlBIndI
xtD9qyW6jx+vNbYylBCNw1QG3eXONwfdvpfBfJaGQE4WVs6RrnMv6Y9RJz1iyqmJJMc4J6yE0mp7
CIAvisK+5IHPXLJ9Lf3pnmsJYc+D5G+9QWEGwDZxjfrPfrSf9ydwwbw5oggPYaEf/cTugox5X1uF
FPAB/CO9U+09Vme10FZsdZq7l3Z0lt02Rkh6dm2timwAKwti/mcxY+KCAtf4VcnIemwgyS6B7lYU
sVfCWa84As3Nr9Kyc4IK5EjUz1VS4gcDlk11p5/b9ElBK8sd4xVUxK4Ga0bMlmi5yNB5mrl1VHh3
OtEC8GAtgPcEELDMDs+KF/K1fGoI9/ghTmX6yDZvbSIkysuBQLRkGpLuPNIpG8pOVZeSvMTTR4A6
V86q6DTrKoyyhx1EJMPk7ZHIzYEzoUnB+Rs80P1aNTUZP08YmNOGNktFrwKUI23pwgpc1v1Rs46m
X+RhblZXI/vNUpA1LLs1dgMIOV0koFsmr03O6cemNCbSlEeGMhOrzKOT2coB+r2FMlqcxWSf3UqM
EAx7tEcJ/kxJr8VvLLtIgCemmzkQJGCSI4LwO5DPFWF1Tj+08L6inkrYwwKm6Wx8FP1oxDPH/UVo
Wx4nawg8vuk1KS3RQP1zamXcnHtXAieh1D8vQl8B0fezBBYvXg/k4C8WGlF4Kr5NjvLJqRYlg63N
Xci9g5WhRn9fmTDPrP+nPvrQ63DFz4csScOQ9mWTEvBcY2N+zk8Ux07WdGUFLl69h3hXiPei7BvU
7IB9nW5I6mDMhIjSllOtl4NN38AeI9u+L09sDTH25McBUiZ2U3UfNtwl/SXwI6sOL6AFJNk0p/1z
XSg36kUhNU3h1mNCK3Iif8mSfUG77z2MBlpx2HvXwD1Y/261cPZIckYSZxvcEG+HSSB84hswn6Xx
fHBxrpgIT5We0MegXZ/krn/AeB19tgGUgSM3oT48o8g7X5eRJDkzBGN82q0RcELkri0rJPYhzY88
bNb/k7cpzm48EWdLAChTbiLrnvIjl5MwVtXOakiX0eVhvnSK05aN12QrPXvqQw3HfvVe7FP0DdNW
A3LA8RMTonRHIAX70Zhl7OdZGIlV3DjbZLN7Jl9POFVu03JyWXh0SAEKDtV3juzRixQxhr1VKV4l
hXSqhSw6IcIzXwrMsQ9rTX+t4fVkOozy7pOAwmjXeKIcOF3zqwJ2BmlTRX1acYMFBskr3vNgIig5
U3/+dw6WhnNeufEHXKuMZ+qfXCOc9jxlj4TeK70y48zjo/IIrjjvmbbRP/vWZ8MfQ2+Hq8p+uYQZ
8Uf4tCuEqy94PRgZVGxROmy23j4WckT9TYl4P2YH3G0Iz49g6h9/9eUFAWM2KLLTyRC91swi9Ex7
4E0streEibxvP901bQr3i/CGuSIe78U/PMrc/mwelmQqMV7Z2hZXBu3S+93OxZO8db9hlEf1xlRu
VF3ZzEwUBgIPhjDfVViO5L9jGheY02KQGsh5u9ZUzDsDl4xJS7Lt9Oovl59V4iX4GsCtNbn0NIx7
cXSlLIjB1aamYL6TYxdNAkXifduoucP7cRHblIm0koqZZqqWN/OtGD6oXCO0mJ37qtzSmAfeC191
uXHmV9GiEAvn+W/ld+15YLbfEbA67fiB7LU64iAWm/wUV16oegf6a67WGZRvgdb1fuq6PGnrmLKu
c14V3hHmtg2OUGLvC6u7ZPEkm2PgUh21rHmNkJdBkiL5Lkkfvz+WL+Zfaw8xiwLFi9Y2DI111qG3
uKkb1+iPd4vzStnXp6YwWg6CvfOZI6WDZpOumtWjihsZiU2LETq/Cp+YbMcd9VHguSKZHZUtHIFz
fuRocCUm+jEcXJdCKq6WU6wpdnY3iLdcQx8nMTrDjQTpX+Z6YtJDfxzU9yRLZgvGcQevRHOQmklb
AjASb91BhibOS4cqerZndodNZc19k5Ko74suIK7cXlJwLv1IBFwJcAmmHWfO+gTa9Xdgt8/fVPQ3
CGQSRaAC/tAQeXQpb4x1CwMqV84XTpqrq4ruUon2e5hfTtbYvOGQCvcWgsNG4iZqeuD0kjhXb/xD
9tn52nHLdWqvsiE0VCcKFD1/gTCYbZuliWpqex7xZy6Gk0O9RvCNwZ7o+/VN8rUgA1ZTKuu/Qwxq
cjoZ9h+M52h6deq9z06mXekiT+45aBOfruKQkqxjj7jojRfOYq6FkFqfA+9tm9K5gdFgiLTL7dpH
+WVXCZiQf3iCxrKzBy5kprFyM840Ks1whD3nFVdg7r6Lmlk/fJGsbmANLH6vZKM4uozeTMiXGRoQ
k1CJUCDv/ESgmO9rCkD7pA8Ajbe/iH5MVD4q/8CIFkXEI/0/J3Uc7+woH20dYxgSjZRulXGi7Yyf
EtYP21jPYsvnPZvEHU6AAgk4jQbgwt7ztnjhVnRC8c6m9ARUy9lVyqu3kHXs+WK2wb+twMw9vWeO
xiGPuKo3iqEoJSuVIqCHtnTgVkLjV4mQdhAPJFyBsmooUlocUpP3iO3pArThGbkY3GAMNNUKxsrX
Vgrb3P8bFoaQMj7Y8orOCcIivYCWFqRRiqQMx9KnODK2U5RROrGdjdAjNDqQ34PRApBNdPTWmMPk
S2ayYhhQerWV4Vjwnvn/gjL9KqF7CobXArsUWa5aYXNqV5aE1wW/UNpVrmARWUIBx+DOcZDpDJNk
N6p/fFffFIdQSLJ3uhS/vBftMj91uVQg/q/csysrb40CYuTDsh/8+lEf1gLyM/cz6Xp0OhSKcguC
NQ2zA2Ril0DuAed43WDBpTBdUHzcU5CAIiLYBaShicBR5Fhk7nMhp5qNssa0Kp4j5exQJKQxuLMQ
RBBlvCdV8if1ToCn8bMjuapY5yaQGR6RCqyl5ee4i4rAzfqnQzYQ8YXrkpZCoo3P6ZFU2/XhfpTt
EDZLQZnS/9Zn2LK4DmJYRO4Ea9PVmXVHgt9jeTsYdH+2DwGvtRvfKAFD6+SO6/vpQawcPqkM1s8c
UQE/R1su8G/1Jfhl5MgtGtsnVJwjV7GiXuxFIqBio9ilhQ0snAgfr/ZDx/XoDyL2nGtIP8seP0lM
pm7H9T7LEdRtym8m68kEx49I1+RH6zJfyJSpmiIbXKJO2icbmMfZLI1quurUZcyVQ8ORsJ9b6cqG
DW7aoYl0l58xDFobv6KjhINIhQ5s8kpIs73Ph0kqAhUj4+6vTlA4JNqrZBpFFxCGk9/3g/JCwCFD
bDGQwosRjYeupIHZ4oHdmZnpqEaoUEZ54M726na377axp39+UIBYNa2iGnPdKUtTwGnAvEYaFYTQ
Hll06/A9xP+fn9dnKyZ7+PNBVKxNxtm7B3OGvHEgvGwdZ7UcJGo4W2M4J9fTX+S3rcArubl13pUY
KiPJPMuXmG94QyLCXULaPIlTXOa2zL5bBi//XHoQIu7B6GdKL4l8f1GAkKBWmLgTCWKC1Gy0VQto
eIP9IbVkgHpryoGt0iDUpmrZ0ty2RPHhqR7cJRf+6OMVMsZ6gyHg5NSbseEv7TwmGTX5kj25cCgc
DAGEhLEtxNr6Bw/YvRxRJ81ZTjZQUV9zvNIvOiUUCWv2bKsj94wFJRn1TvuyHGVuTZGFj+Bb3ZaD
CkzOctIhgbpZiDDYbXLR0HGDH296FHcynE7tMD78mZ5tryyLn8abnWIF9EZSLsqt5K7xQJl6SQ4I
khswTCxDJjaCiunSoUEquOgS+q+ZMG3qADMG1y91kyt6vP4IC8WFIMcyTMFkVTnCo2WguM8kIMuU
HDQVV3C1G9U7NhjcFhj4gdzdjmkpl4b6s2BcW6tpEij7RLcYOL3Ji2cmltRCR9uDwdpEMsKHPGUJ
zI6RRCoCFOuzgZlviv24Xh7zPprcT5daJc1LJnw2FVje0qNZtfvGBj4ZZBNMPHAFKz93J1n4UXHD
fkx4HPYAIj12V7GFc1eduLBEcpRE7N7O/Td6dMUCf3H1q4/qizzNdJAAfyDSyrpQpioYXN2nQ8ac
L7YWa/tX1S1oc74mr1lk50H9vER4camFHZ4awCQJQWVJ7Px4BiJrqSFaSo+dE0Sd4RbRCnxwuZXM
d35D6bdv8pJP0AeFqqANyfOJyAumcYMr3LHufxBpdtGAAUGLQXo6YPYR5Rk2ZsT6Fr012hXnzXWz
eA5rXnqUs+UT0Gi9eLyJCDR3q/7DzeYbR2AM6K7KViIDuoRSgxZwVG4WcAKZTkrtrTANIZ2222fo
FCmKxWfwRvSrib/6EV+/AVs8+lCPoEUR746SYayMVn0ol8/q87kgpSBbvORYem/5SeVrPzat+e8T
h1yd+ltRxOKxsMchIHvkZVby5bMzi/2n67K2+Ns//m4Nx8Eu5ioY1YhZwBIGIoZlALPzrGZNwTui
wUT5p+l/Q6l9Br7V4+OSZEnoHl6coMAjnCGTJQR4adnFMrbSCmWOXXLoxgSY+3l5C3pdeHrpjFVT
3BPj2/KX5jHMu3Fvuzl25U2HJ+XuREEcZxkpoiYNPThsZywLoYkN6ibPkn+gn+fH+0v47Xr9GQcL
oSTFYcRmF8L7KFXR69CnsGg83+S0YCDvZbnMxl/7ZYlYAyEpjf7mJUHhxhCxZ1iqSc1ajPTXeRDb
4EDOPaAjtaY7HOv4VuVA+PGQrbItVVuO39AT+QuOS+U13Jsv4s8ZTGpN1t7WCf8m+fVkCkbnmVjI
Lip6r4pQSbf0MBVbPwLTjB5zu1I/qvS0rGRqYoX8ABk7cX7gTIfejQXe69XeGmb3RX0dIJg8zMKA
SoyYEgNd+hpwSj5rVVm+gJmjjG3JtVEFwWD/gxMANnq3tnnkK9QfrO4Ir/FODvG7nSEnraeAimQe
Q7+qoiaepQhU0ytFR+1ACcNEUNU8ADlJ5ONlTSfuZKO6LL1QxUDMrzUzQWKsQi92L+ftq/K8gePL
b6M1dxYIqheBEHRmvQn9djwhwvzU1UX9hQwtzfaMgIkSxqrAJm/tju9fhh1AAnQXFOkvvtGqVpZq
IOELlZMM9+F+DhLGNzNlEy78KbT4T1imUTcuK7+sVt2qnVK9EZdmZmtP5s0Pxw7ICf47fX2L6bzJ
gQG7aKALvAeiOmSno5yQ/Kdyz6oIA2ZbEBCOTdKMn/7kgmA+lm/vGOO9KseCaqyJyB8zIRTbD87r
7gI2KCItuPnhdJPtf45h2UtuZENeHHzHx9gY6EUf7qnZX+M15vb6zF5g9aq1ANa5T74KWXPTVrnG
jXwzcyu4WAKCV97IKKtluykbEu1RcXGTefO53azSq2RHgzP4uM+Wtp+R45Dr1ZEBYX8ugb7WonUB
VrHaKrdfF0Wv5mSY3nXgt592O3VKnDH6GQNAQiyP+KTu10Mta/247Rb2F6Kqa+tQ5judvfFk7q2e
NgNUz+04ZmrNKWQgbHPrP6+qxLivOpRiFMC8QHKTjLAWBjoBEaCKWzRzKgWD1nQ/m5GoCbcMwqD2
HzfDvuNjnLtcpYBvKpCGyKv1SHvUM7AFGW4onvEpio5Cxm0tFp+L4TARRPFLYaJl7oUrnoNEMFXK
r1kHP5hYzkbDwgRW9o13fjrrZca7C3fX8QNeMcOjhE4eBrF6o9197mbttTaQM0/VeYH1j/4cLlzu
nhOzqItMAq/FyCGswDwboQtG8dOjw6HDIUz51KTnPVQxbtoY7E9WYwPJSpyTfz4rq+p0JbEdC1IB
HAnBv/h7cWjDr4ejsoJ7+T9OeXyE3Dva949UTlx2KorFDMj46xXETgIPqqb2u6kVP64vqpo0WPZE
cDOdNB3khImaUo+9vINZdhYXU2ejAfYGq62l8I8uZYI9sQ4Pg0vHhB+Ibc4RX+pjWD7kInGWQEO1
cSmDcTKPlOzjN5XfvK2G7jZDOAzUNMQ5jIRdii/AY0iyrg+oWRg8uxrVJvhUNJSTALIlgJW0AgnC
wU0Sy7YLn/1YaP8bMo5+wXUB3fVOMrwHdMO26Vb6z5/diN9hDezlOxE966FjYWngn41qhFlPUzUl
nz6uE6xaNi4tF+DHq+Vc3d+/YxYWUQzur5BpgEEOqWqZ+RmOvqIyq2CGgiBw/s8ebMvUaG8//xcu
ekoAu7smJIKDP0XvobrCEZS5iy0boiG7MDQEMdVMg3h8AeIzqdcjrILIbAVMSHRIjCgYuef16WIi
m8JnG618NdOMl2f2F7IUeoW1Soc7BthfI4jBY+qYSQPf6YSie+SZbK/P0UVAfA2+rNA09/2GzwNB
TSW17ek5yLU1HkCl4onxNGLS/jXJNhaEB9hMlVDGJLlCl5W7Mz0Xf9cGpL1/qBkP5k5WRjl4h3KZ
VaCOygrnFVuehyTO1/Rv3/sVOIrVO7SVeZpmIQJwSBXtj/stq3rkz8CCo3Ntnpsv+9tEE7i+GeAf
zdww5oNi6b5PlMeHhyMFAzCzGw7yTCHLWA/aXwf5YUXPdJr9aiQ64ozWL8+dUQgVNuLumjJp6HXC
UxpWp6SafSrN1qgsAKSsw9GLvEAsIjA9puVx5Wq+1lE//CGYY3LzmPOonf8xu0xmBHXyGJC8PEDL
R2Jv7kbPGG7gUZ93dChNEN+PPa9isviO5P5/sUY5aQypVAdzj4WqGHoyQ8MImmsuaazqhSsZ0o94
2+JhiyzzrxH93G8GodWT1kr1SltDhrTRowkJCbMji/eGGmnZB06eNxqRkx8Hom3Dp0UhYlCM6+Fo
QCuDAUM9U0UXdCTN6n60At1Ju6Zx28Xl1U/h1b78djdmX5pnXb3h6TC9XbqvQF3OprzsV19nbCWc
ayw/enu8W/e1eHOMUn8tVejD8d7SMAH+hfRX3a6QlL9CBpy9o6FbBf/tGXcFR/g+Z03j8t8ZFBzF
gzKrqewkh1hOf8xztYGTDlaql1faruo48YF+XMCHl/jPxTzm8ZMCOqGYTFfOjpsYFxhNLc3BxaV0
93oePk6NFit1x1mgzr4qh8+bfTC1v/VRqOxAlLTWvFGRjKPFrryhesi/lW+LW8+Upct3uY0g0s5p
R8frEID0gcldkjFy49aFPFnNz7ttZHb1mZ/xNzxRzWl4f8oO8nHxEHmTcEbnAhMw2N2QtF5/oqTn
7x65VrNgqiNLWH8bBDGxpN5umzGRejI7PA3WYjTS/jkvMFiqoS0gcNMbfkJZHn0JAmPwmJz6c7ir
jndklifTS9+kV7h8EnyG4O1AodQA5FzdmtrwNvcxpHewiQbHy+fSIsyV+0CUymhz5JR9DRuyWFld
4mwrT6C9BjFGVKVG8wl2dwx9nOAsFbX13py5HUQ1y62qA2X/wa7xX8d28W3lVV26s/0KDVYSCfm2
sEJNGaLySW1p/Ykvq7j9cW1+frPj/F/C6KGasejuDqi0JHBN4ULaDWFlB5LRE2pAQayi8KQOoJqK
ME2oNujjOvMmXmwI7SjBvpUm+51edjA/npND8JO128BmjbPQG23Cy3IGo3KyuqwmGQLA17q37V+8
1IRrDvdciei6SlhrxujXMC8yfddGjVYSyNnb/91eDIhGK4tV46p2esAiC/lIXG25HKLOX97oyZHY
egUu3m5tuyLljMVKje2fu1qr5RQTis/2FoNagGGYM3lDm1Xr7jXxcoKbLBCy8kK0NV/v4LAFci+T
Zxx3PvRr9q4FtYbip/tA5CVcTcqwcoyuskqcB/Nl1OxL0CeY3+2BBl5rSLRZZW9y0LU0oBdNFISv
beIQTVAHW6wz3Vd6ss9MfoQ6aZCTYWvMoZLXqvUW9bRn95IgHzZLebqzYvcVQZyTmvXXyonrwmI9
8IEUEaCczsONfsmmoD7lLgvK3NbEjzOcQyyHMEHfsLUza904TSZvyWYS9hTh8nGQbKWL5aEkJiQH
k1UbY1ayLT+0jdxQfAmCTHDGymHxNnhnBwCmoaS76y7V3yLN+9lvZJmhZ+H2YHGybHsh25BApaxa
hYfP31HiiRf7YpbrZhukZeoUghUDcuAaCevmDYSj0L3QfV+MhiFoZic0RcPYsfF7Kc/V2r2rycNY
OH1lToM/28Sd3TSjSxXfXNISdIeZjr02uE2wtTr2WiF9BY9X8Zzy5DrtemBnnKc9nCi103eo9ubk
oaiKgjwwBEfqTH6mvaZvbcZfjKy/Pg2c320jTlJHbgvMj+ZRJpBE0yyHnYzyWYYYXnGYhhAGcCz2
Ui8ogJ5EDuHgCWtVcHyjfavyQApS+qn3e6AD6EVA6Wk+EkJ+/ahj8X+G4JGF2nARibeSN24pAn2S
N+xEecEVednsDsVzfp7ky1kfpKNqQ/1jKbJiYQBIBV2jN5X8e1+pq03vx3joHq3xUkoNmlvW8i1O
F9a14iCJbvttOZoSqO42HYiJMe1bANXFZydGYAhSud3dB+25ueEw0UFKb0ygCh/APXDRS0YG50B9
06Ka/owKOKAP2tJC13ZhknBX2dIlGjW8uNngI7gRjXgcF6wiN+cAPqDBxEkQtjpTnxJxWgdtWiv8
6Uv2/Yo7bTFIB74pb7jzv011CEZQ3JG4RN8xqWtf2fdZe4n5YwGWSLufhE1YWAaJc9QRx2g9YrVt
5aER74mSzxKe/2rjEH4O5aC8BpnzR/l27NxCQo32T+ycbKTMH9DaEKy9D2n1/uaMsm2+sAbLwmkl
74vLeDx/1gjjNE2rC0XP5eMv5FRHUF96ntVQ8n4boAr1CeyVBlEJHQBtl42jzV1AIWcYNceignsX
nLirOgKdrEveZvsHKARNhVVVROwAnLtLbwDyEQKAkvllutfKFJam+6zscf8lLviB7j4AREaZeyGi
9ofsvZeAwP4+TylDOUh1pgabAOJWhqkhpwofemDL99k0TXHq1sHP8R8lAbxZl6nvCWQtYqAezbTf
H0sPjbYkqLkFjbx4vp2ZAYVzP1ekJxaxQlpt12bZ9o1FM5NISwHRRBMtoeoCpRgD+rswQBiiCq91
w6+8KV53BUEokAlPl0MnhIFy0ed/vH+QnhCyv+pzppTBhVZxUOwfUsYehXvQmvSEK1sVoTFDXJVp
lfczfWK2JoZAMRR/IHKPFXYck2P8EVjzLnaJPoJh8dYoQTraTAz2Y3efz73+8WVdCGLWXsJaYzDK
mhQSIChPye422iaa7o85gl7B6NKXJ8t8WqJbac3XOyTU40+BH/b/fDhJfhMG/i/u1pmCVxhiRM65
R0FqORyjPK4Yu80sa7jl10tWjw8fampWnshG+e/+TUqU9QmsZ0LPFyVDkX9xiHnftdG4RhKjRNwe
fLbXal65RIGOZIHlqV8R/vQ/d7a60oBjo+VoU/3doAGvrzW3zd7C/6TKH81EEHQKxvXaUG0coayj
PtbcDgKHunv2gD9d/cWKzcj6lMp9e9Zsy5kr+OpVQlnpE/H79G/h+Ga/WL64YEiD0OYiD96zaYbl
SWtvAxvNmaoF7fRb+Jm2qAwwJa8ng44kMiDLP+pzh6MgkmdK72nzlErJX3sL1f/iCTdfyLfYbI28
61UYlOPl352735H6jeIqVhmW4sSQUFc1ZvbuhF8rH5uK6ByP/2ukeH1oh3rAfv0rnUI9HbU1LVZh
lKrmEN4STNBVRRsNHpILZK2DEOK9TKyAKEChTIrhndPnTK/knHyuKZMd9ZUeiYUmWO4BGPkqW5Jd
lMKftFfTqbn5EIt1/v9epI4MeUN9NLJ90q209dZRSKIuTpdmdMobR5wqfIM6bqLQ8M24FBBjhZST
ep6CGUfLdjE8g4yfbUIehuF8EdHmqJfEeONC9s8taeGniIs0jmC6kdIpOC9VFwE880BA52ioGB46
m8BRUnkYffL8qLmolLxrTdVWqAWJbKKx0wQNp8Grqzm6zV37kNz4BAbHQ/PEGIeky+wFhLlli4sq
fNPv/JxhxO6DCKDAijmMNdu/F8hepz9zKW1keiLlc0EQ3CeZczBlL8jXk9MRr07xnA0csdkEGeW9
w8tBmBko1C5juRS5MMIW1R3R9LIYXIeqGK0E6VpHOAoj/0KOpA0+cLjU2OqhR2fmcETDNS6VBZVg
/hjH8ApV/c5sI8bREypwlD6XHiFV4swiIzcOwYWctfQ2BZHfExR+O8DNXSvztiYk5ZdjFRg1s8jz
EhzfZH413Tcg4tx/ssTpynd7o1nijRN5E8t4dJOm4WxZz6vbGfteCShaWRMF4YwWJ1O/KG/J9jr7
W/dIv4FyTiGuHMetfoMkHciYpIrAdEeO8RiOW1ApwVC8HBU/EAbYl8cLsptXuAysLYvNlvPK+Mrp
M0veARpdgwJiZn1SSsyAkBMDNLLvqdfj6G1advVYXRxFKZXkfRPQMg7UxShyUdXy86E6e4mgvI4X
4OxQFadCl2PjISIWP0xQwHG0/sfabSW1MlPQrhZLT9nWbf4YHOcz3ttqbhiRzuSyc3NXnszgU0Ou
uY4Hvom+wZyXp9+W48fClKjRYGH56rdBBDf+aQ2yTlO6xbHrLPJ///2Wfv0YXo6i6aMto2KHQHT6
FldpeM74Id8twrWeKGSuxd1rlcTuUWSOa3bCxWjxz26+dnFM/g9QrmuV/QxpMRbggxtz3E1epDEE
893B/uhsQvAwxJTriwUJL6cMbL+kpQLUfe4HrXI5KW80uHejbJhzZck3/M34ep/0S2OZaKvQC+kJ
C/Jt8JK/31kVouDjLuwoQr5Xh89tHBobn3hFYumKG9NoI/LnrAZC6nwOEZ6CTCJI6jFhBxJRushF
5XJ0JgDBmHOlOuFjX/rLPjn+DFMHfMbMcPbE6pNfjHF85wrK8WLNj1fMBWsOL0/5s9ONLdXOy9mw
qYAQTFWun7A6sybVcjZHASdfhBwr7RYtv64ctrhPGJF1Pm41xL5EXrq8Bm5k2VVBf3W/lCgKEwLe
z6Wgry5XcLELn2onqcFP/lzG0dE4568GIq77ae9OlIC3JdooFElVpjeAV9aYidwQ0O4maYxshLHG
e4j2nRyWHNnLA+Ml7dW57hmkF8ZTsxU4jWYxKF2l5tm3p2jgQjJKgVfwUFabSPVlTIzUj8Lt6ZTO
x4xWWwj8jEyDwGRuDc68fgIOeSrSicNErgDebRKYjE9KLKugfb1qLd4pqQzTn1dsWsJ+1PN5XXp3
p3bWjYIRBLHTE9CAA2z+DWFSdIu8wgAEWtHwthGTOwy4Lscl2bYJO9BeNer5NVKMXR9sz9rRoFHZ
clxoRX4wUgj5usUqMsiLogZUisAr1uza5AP9v3Q3rNP/p0T//WKzRJx/UMzS6hWg/PDBdzBVkLKE
yfHQBNT9rd2vvh/G9UUW4nwd+kDbCKywC9nTb409cRjHuWTbB0XD9NtVOukxXHGcd5XEpz6U+S4H
aqZdQHgkE6aHpFJQJ39GHCD1EhcMpLAtzJgl4EVQKk52N5+BX98H0EzuTgQm72VPfCykEIG0rvAH
X31iNb/5k5SDOHwiMgXg/km7y1qwB5CCSpbTLUhtLUAydtin99siI1lR7wzpZ42ifG3FS7SOiY+Q
s1nsDMs4RYc70c1gA4pPziX/JhoIhYqrSS3L558mo/En//mPllZLNbHX9++gMiWXFJR9FE5iANjS
qlPhwiOqQwH0FGRPx+0ASK1Lf+CTavR2ns+QpMUGCy7nmAtxYsGp7W8Z09iclFroYkVICSEPkmkJ
WXtI+0+MugRCPxmdxdkayPrmmhkSA+JGI3McMTssPdlBs7aEjK1xXSLzH02r45eApECXmXASrJc0
OJ4qs24AIY6S7Qx6ruFexPdH0IyqZG+cr68GHDRRi70Cf8+sgYamiRL5pdCSQsMl3XbKC+IM12Se
cmd5h6qIzaCSuaPCizJ5aUyn5ySl9ffhlFTR+EVr20eyuq+/YjwwRSYqxDz8RVQ/UjB7biBM1tTC
FjLnpOwrbCeg04U6I7HBZmGygQnFik1RcSVZvu9/BYeTdsBWpBKEoJkRR6rkeTB8Pd4zLaJQEADc
7zLsICWWp0GxeMLbGWfIOsW2M8ItT/c+Ckg8qc8ooAFbkcjm4ifPP5H0iCRSdrlxNFa5v8hpm8ek
EPFU1NPvmBgVW8ZR6s9Gf62Kn8+403Hs1qEK/y/A2B/S0Gh3cadj8yWyarSijMFOUWIME2ek1ax9
mXMTSMdBpMpTJc6zSKetOYa62KKZ/ohPuPpmpGcE3paCPhE8ICR0FNamYKwUIIOAxaDokm8A7Zaz
v0TqY+cf9mrTex57QNqeMG0ctbL/WNKXYZuJ9o8vhZE0FHpZckln3V2ICVxoVjbOjZVMwYdiLYSD
gBa2srgJiE0QzlbdCzMJNVgKhJ7Y15hGchskoyLe4rm4WxjRGXq/ZOL+HGwniC89snum0Pz/mMyE
/GreNKiuJHZxQTA+xoHd74ckx3FN4OVQgQs5VRO/NfXYwFoB2YwkCVWvfLzNCeE7AUyEq37OCreJ
cNHYGuS60mz3gg7KfdCbvJbFOWONNJ4+5rnXlranx7Z+HwIzdPjRU6TU3eBc+RpCB9XGH0iUhGZp
4C0g8++Pma++uFMZz+ddlexYlO7vy8/RdUF0mZpQ52lDmrcSooun0BJ9lNZ38XlR+3DBfttmA83f
ESqCgEzeHebTZ8hXfA9ZyaLxAwaeD96p4rYBUSX6e5xJ2OoZRG6B4QBKjScYIFt5olc4PY+/1a/6
a8ri2J90G3P6yGl0GTs1QPq4ktVJaqMNyi367IKIxl52RRvDzq2bwAcjuCKSNMWl31uvDIy+s/JB
6waDJg7DkM7g0QY1nxA0Vat+Ov/2E0FMhoyBAe9IQ5cWCD8Ai5zE+WUWY+85sja61Op1CNMiVEcx
RQUY/jylJnFfBo6NbAPJ7jWvfPQ5yh3gznfTiQUdzwhFT4u14/XqkiyE4fr33/Iy+S/z2lY5lEp6
RpcECQ5hfd6KJaYkPzKAkBRatgN1FfSxhstargwIs6bP/nr9kfzwhAC37QMErZCiMmI5N+n7ZxUh
P5HKdcZhzcWKxuZ5KJBTjIrgO/R7+cHptQC1Enl+sspGCszOzyv5ZG6MBJJogXBBEImLQZz9Xc1+
iN07K0iOQJa8NELnQ8JuewWcQZ7JKX/PQGFEVlRau6ZW1HWCt3KUY56qncPHk23gPN1IIEgD/Uy9
n9CesYXJTGk3CNalCjS3Gb+YqYh7loMkQ2j030BQeHEQWCg0c31NPnE0VhxA+cP/2LoNRK7+ZdkG
94odmAxWYkdoWRQgERDuO94fu70p/9FYh4h6gmp04M8oS76+NMrZuvUjCTOMtHkqz+Vwy3ob5DCi
gqVV0nAPLyTWt6QkCRC0YS0cDom3cBNWczAp2/rqiaYgrWtYUTSlVOG1gbUlXFWQrnYEBO3U9JsS
A6A4fPXxeNbWxC4Gb0ZVDF+vnB6V6rO85OSIbyFMIcgeQos7vDVCFP7+uyQmUm+xnVTHWzkz1t42
cxdeuCRb4ZO0MMXkPuyEUpec0Dn5UT6W4sK7qAM+HqqS5XpNK2fumNYHUqi/+KxVcfRXLLp1PwXP
jcL9S5e/l9Bm5F2gq+b6uX3mIyShxDrC8xWZkVUKQFOgFlzJgzYM8yxwPHYk7nkDXX04bmaO+OD7
sDP9OmozvO94WQCxEKp74e897SsOtVz+iw7UpoNrvRF4gVzLMkYzBjxZt7vk650uT5CMUzHAQ/M0
TwcAf6DSSqoNmVPGjFfGXR9RhyF2QwmCXfaeiGjdJa4EN9Pj3XCsEspNtF6EsY/uyCmcvGGKWV/W
O2ERUwDeY4ra6b8EDw/Ftgr8oF9Uw6KQWcz9CcQvCYWCbHGIKJaZQ41uMAzAPmSTz+SS7aoklj2G
/aLOIWNW7Xa/K20UfMq9lGTUqKu/Pp46I89aUqX2FgGyxFG2GJF4gEYC3Bi3UyjU+GUmXxw9MjmH
jd/TYPkhe+HwywqAOqYwlUEhwoaUMuycIHfb3ds3c2ZEX8RqGRYbBQRDHhWg1jUimh7N6AquZNJr
8MT7TeAvpcjmSF1yy3NI/3HjObnU1N5/aorOIiQYNAJIph8jafmb88pjcvA8u+q8pcNok3sW+cdR
UEgJvy3oyvILBPNELpnSKy7LDiRHdFBEnPdNgUoMgmLSDv0Cou//l1mNShgLtCfvlu4vqIB+Prh8
Kdo3Qnui+KQXSV0YaL6qjEtdZti1cxWeOOb8Rl6dWa+YQR38L6SLNfD34hCBYWlvxpDbb4+34YjJ
FQlQE855En89KWm3kyqq4iaycDRnW5hu1y793kN4Mvnq0FeD7DY5fIhWt7sPj1t6EBjchINwjvl7
JvV7vws3Ys9QCIL4Rk1TYxzsnH3wkZBrQm/cbNOuN18HwkyYot8vjVXRKAEbMmQ45XSA2YtwEAKe
lRbW9Aq1NaH6aL92051ajinE9l08tfoime/Kub/KqlXjAuH04la5+xKTQz9ptotHY7a2Njy4mGz/
g8dTP9FjyAjvSCakFdRwdjIZyiESz5O/QGgBBSWIQ03KXedqBxHy2jiX4B/lGZtbR35ehCpGETuK
/FqL2s+CruDTubiPg27TJF1nJGi6lFAyBef2bqS+HmwgV93lLlgAftegAIugzxrodCFlrNKfm6wO
L1W8Wt16oqGWlRAaRWP1zGVUaWDVg+nKKn6rEw8pCiAA0KOdZ+3OFPrpxCykCjfYmKjaO4QZIggg
2VoAjQPkNZRYmFrmyJXSBfnW10O9iNjzl6No74/vrCeP86aMov4SttkeEDmdTRAEspVSsYttydAA
6XoQLyISpAIKpcquZk2pmARIot0hs8Lr5Ty1rfCDCR5uaoJXmBSJOgUjnR6xstRFmVfWXI2+pibF
MFV4UiHxGT2vB8lj5WF1IcEHZQ4HnL1aL/M3Fio4maqI+vsUHPZG9KmprBK2NAh4/XeTS1IST+bJ
ywdYue9YGosMtjOKy7qI0Ya//bzaq5O2paEb/Hf2H5NN++oVNjMFvrEdet7MSS0c+zODlsiQRFpj
TzcCi9lQBZWopewd+VdfDT9xJ32cAT4WyQKirlwoWvcVMg/J2r/7hewQR+kxkwm3j9UAlVpk9w0Y
7afjKnYgvUnxy6SSyAwXYWMENwTJrin4/UFx3d9eOp/MhF0yUHIjqtKiTlVApoUBE/n+30HV6G5Z
OUzxjXz+80e4Gb+UOa2+ueANBfjdzotW2XvYXtfmnN57XkjyN3g4a1UnbNSK/Zq/KLpjyn8dz9im
xQTMScQX8dhfMjtAE8Fto7/J+ywRNObBzVOpVxzK+vl7JXeeGTzK/ravsSys8JU3tyagrcf2XxvD
MRSaoqehAkY1KEUiHlWp8RT7IvuXY4lbCraagDOu32vLCQ6w/xOrNS2rd0yitZ6D1nBFknL1qAcf
17J4DrXM3mvwoMb1zeb4caiCMq8BVfkQXKTBSeIawGvHJrC9Xr51MNtCUGYMC5CDestNJ24BQtr9
j24O61uZ+XLFdZeqAIVDgKR/H9LjFboX/GS93UE7FHisItTMj74Ig5mykHyTqqRk20hNhvGGnzg3
RRkQ/wvo1aZgh7cYPqI/F7qLg2QDZRkC4xXRhPoSb5RLRf9sEgJphqOZ0gua9ibFgWwXmMJjuTm+
Mhll2GIJSoMVDEeNUIJ3WfQpGeSPDu6D1+EEhmRxA0i+nFUXPEmNDwMnRNa/XWWem3JxgAEAKDjY
LFuw9/MoRvj8GGlnI+pVTcE5XYzCuImx3rZkvAemoejuiQZbYuSw/CoHAWDBEqw/FHpJvT0TgGRS
Nv0aVqP16H5COtN+iWQQZzf1nZ47CWWLv13JwFZjsT1z2qNoG3SsKq5kzopck8gMHECA9KOCxBJX
UPHiusm+TpBA7aHwwXO7l5QbozkbGN+PO2QrZn341RPH6UarrzB+BQeGry5EMfiGwiWRcdVrO2HS
cLYEDtkcD0IK11DuCSl1er3rAJk6Y7ku/G5An2ZU94YSGyX3RsJHlv7LgjO2bvpB39qkzR7Q13N5
Pf4OvHEzf7QT/xnemBJZHTUD8L0AGQezIYvrd8peR3qfL7oazH/+y1uEo0KWDlGRwuBSp7Rie7ou
k3LHOTV7VXRlaJBjpNbfhMVsQtc4x3xswM7Zi/VbJD2qU7+iTTMwSJEHNcWqR34VSK+xymQXDf6Q
Y8fPaH6P4ipS95q3Y2PMWORY9/iiNEB6cZeYQ6hK8k0Bd96daXkN4VmbG/sogn9DyC8yQsD/cay6
QwkFf94CZAcuUPya2WjITUMMk6LWyLRZVNEuw7s9vhiFxpHmPYkHG7O6SyEl19+Bin2j3umWngUq
AbjfO1QsGgl3renGl2hJc8sNKjOWchs+TuTEYuU0i7NPWEE70KB51ZyyXCjC0+ZM0L/f/+/CO/lG
63lEBCC/HzD788boITsDmhEfJnbSiUubgnZasQzBu7fsy2XMNDR37VGezqUmhh54xfD4FpW3Yq66
ZnRTLU2jUqpauH7ADEloMidaiJrj+mycsyA2UenoIHNmgkkt6sA679wdIWlOxnlVa5jy3dRIazLf
DIItfFMo4B/qLn7uMFeVN3pnzlgw9272A2tgLmHwv3Dx4DpJ5fOMRIAICY16Xfz+SoWHY7/3I3J+
31f4sX9k/tc/dzlg+FNLBg7PCLFZgz4G9CcKUUKcpH6kjh6+GUKXccIeIaFpWjWEjR0VIT6rpsMc
dw5mTGzBpHv2v/wGuyqZC1qIZU5Ckt5Rzagc31Yg3oT5J3zPGZEhIq3FT0vtNDZ42izTDBKz4bOE
rkzoUXkcZDz9vKeaLvyZ+izxPeyn/9hf/YHBRufiaVzwKz2rZx3WjUeXjbDdPPf2vc9GQ42H++8Y
qzjiYZ1Gyt3FVXqNlA1qEInqxKV1YHUCAXNxZSVfvbvvbP9G7Lf9aAHYPgxl7vHJ5Hvai/exgY4O
Zyl7PoE8S1P6P4G1bOVI4iztbXEOPe5lTeD4Su3jeKadD4Oo4+2Q6beSC2EVoXQYtccyfiwYBhLF
Xzs+t1Cr9iOpGA/ZwORJ5rI8ezmz6jp/f4a2q24VS1tauer+s1GNw5SHnJK8G4mHlXNV/uYGmR27
EMp6eVhqX78XPA4Cw7SoloCiTxVAYzWf2bMi/JxrFKWdbGmyA73e1u27KcTOophfRkl1cUhUktQY
Klv1F5k/vyTKa6/Ipw7N6bnXiWAY5FfN11haiaXsWRvjFZbjSNN/5EBsbnqVX2axiW1iiOZYdLyh
RHDOrZg0u9va+Jsu2Qa5ux/bBFGhgE0Vx+TKhq4j0GplKNIQNOqxR6Ly/zzKz5xlGYzSDj8+fBIn
SCUtVTvrbnfkfHtRsx3LwHIv/SrgRA0pwr5UKkfwBNkC4Bwr6RbfDjlw/jmIWY/cUV1urqLD6WZE
y0V+I1Fym4idbZpQTbkEItDE7a87cNIPKdqJyEJHCnDq4QAFg7N9dn9OOwR9yaQK0bkLSzqDNSzg
PThJuw+s9mKU4lJhJiT1Z8CY92ILi7lN+4BlLUiLZLB85cNj+X+Dq9HIm4dMX0+3wmQ/4mt5s5oH
Nw0/KJrOelxAGkZA+s4jyfRiKLq5WUzN/CqvwE6H6RbaHU/+WKEmuwq7HsxMxMaRRBGjHJaF/m+q
0WfInrJ+l/fgBFYfCSjs5mwQMoBXsw/8genidcxlCejAtS6yiknKFSYqG5qa3Z3qRtm5WPxrBzqE
n9VBEY1stF9dlsO/3QWl+pKVq+dSprb9YcJdAhaMs36fj6nHqoDaQE60hHsgZI33WA90XwJ5AoQy
x8PkaapmIyDTldrbpmWMwmQ0BbhO82FwMa6bYZ9skQG35kNI9CdL/YyGZl//99HzU0FaKRn/bEUT
IFXgKlLkvOVG57S3Fg8WwxlFT0x/lQeSght5ANtby5vpbL0ycHiaclSphReJZOzsyRjOGdfTIOkJ
mMj6jjKLrAewf9bQXCVyvvOednJmJgNhvHsahk25g1s8OSJOmh33mOkzW8HcH8htEaH4BxMxvtNM
crXHj1nG7FGYbhzmXlRT+BAPfUgLBJvMt72KxWBLDAWP4aeMDBRWkRHiXnpyUbSA1TRXaWKteLP5
UVVHDFCcjSVwFkJEph/CtoBTYrIkFm744YhWwkAc5+kpLLYkEanfrO1kKeanYwSDuyA5RpkW+nRX
O8BDTtR4NaC0nBMeUg+rYodUbRZYbmFnLC2R4HcXrExMw3KSQYvcR0l7zIPEELiNCaI/KHPnX3pO
J/AWjU3tHWUmmQfkJpr2JR14Kwl4WS73QHIYw2g5wY6aPVuOs6P79wxz73QCiyS582FJxsUkpq3z
mQ/+feXWhPHiCvxkcpMyWU5ssYIB3FREJyD1CyVi+WkvzejtDrLzSnGqBKgNBErUaAHHJL6bFjbR
nS5tOfGFMMJ+xaLs5FMFKkdKbSZahcyN6JofY6kc/b2q5wtPr+iuktcESdqC6aDdMonHOoZzQz+F
pOqo0Q/nE0ibSwQ3R0f2717UMFL6ryXOMxi1YjAJo5LGERzmGCCRWNKsW0LlXVnXvcsnJQv4IqhJ
IYAYmmQ2YV0m7Qr72/HG+52DDOJ8Z1qs4/WezIzBqF1j82wVrlH5u07hevX9hw3/LNL0vR/8RASv
JukxQL5xK8lWhFTC0fc5ybcbbWWSatNQvGGWvvCFqdiqJMcN4/yRhi3C83ZvSa3CWWoQ0kcYv837
8EF7aR7d38CKmPJA/n7nixw/4KOspOcWB3ijWk4NsN7IOhSyCQprTD3VFR/L42k45NDrSOMieDxs
u57q3hZ8w2nz7gy7l8JCxeey7bVDoo3qYFy4zh37beAOK1QxJglwcdHirQLpPY930josrjjSmg/I
fdSMF+gDtXmPns0KmbYzRjbvC1Po1oLQ2rfhrikdQDwOhqzt3PavW9OloiedjfRifvvmi+7NV+7A
pWmIsDQn/LJrPL2+TtBF5LkMn475WK+kOk5+NTTFjq968hdVQ+TuwKngXGOHz9mDKk6Nabol839j
Co8Ja6r0bigJwe8u6fLDDV0fUwzxj+3DrJ422DdO3WaSg3uwWORSkB808h59CcsXihOqHckRCnpZ
y8iwSfOZ6puSwtvd3cBO8CVQQd9ikR0+GxvoocXQ4ZUBdD8sWRfVz8gFX/6Hfhl2juHAxqjAW038
fbgYRlw6Qs8p+/8nSvOg2l8T/K7wGcTCw2ohnz7/K5Hl/htqQJ6rPzkLQzoHttkY2FoxTHRKpTok
P0oOIYZZi6B/t/AQvHkuOvW9+KIYbL4xHuUlP7noqdE8TmlrwlUuQ8uqvdBh75zkGbX0rZkUuAiS
V0V5ry3/sRY/dfju3lUkhcLsJgtMRNZr/ubDFIwhUF6MaYc6febmCC3yDKXewndmOMsAFrMuTK5I
2iMKAcxf9MXhPfGZsg4iNRYLJNvWfXK4/F3LeoPix7QmHMesVcR5qsfxlILrzDe/1XQ2PqDgje65
5R4pG5EX8YN3uMqAwzLeEFe7YB57s1DJL7Zsckg1+4IQSe/+0bE4cLWmPl99q6FcgoYM31BRdgPk
PVUNnHT1u9syeQ2AspvmljDze/90ChPewoS1vSvtwwEu5VFr2jLD5D0ZR51qU8nvCgGaXf65Qh+H
dRydBlp/7G8/OrOb437NAofxkKPLG4h41XBT81Zp3L6IQHj6O8SBZZRwID+BmuemahzH378hk/hU
HWXFI3fwzJlU2Rq1wmUVpiapFL/D9uxHyvYO4ixaWJV3jLmVmZ/amOfEz5e811n8wgZsv8ntStV0
25fm06WgJCyPVmAViIb6D+Q+CGBI8VywLhL9ZZ3gamRDrQ5BaEqEJUorbJSSW90VF81z5BySlxs2
T22K2wpufwOsoyq9KMflyPf/9VRlaJ0ixoQiKRRc+OEyHE4ceUoNx8oO8wDy+BlIJ29w6BCaoLfl
/JGvrm6/kRg4dYUvSwae+lxZtyDCi5cY/gB3JsjRzUvJeBXu3iFg6nD3LQXMC4/t7hGsO+/LMpEj
l5AqM4NK9xDVt+tRlfdbPMjrFcYz8cLp88RDbh+NpOU7AEFIfdDxloEILXzdYbrgUb9PW/zDPg+q
3H9JWJgBpBQwjp+chRSyJV7Kzk3Umnxbe+5x6CtvR3bLfz116UQGY8Nd743r2YLIni8KN73FwCS2
hrl4UKUmsRejx9gmy/L3Pof6FfaBtpwTmXJa4KuP6KEXaD6JSyABrjKy8CefBBQP2igu38z4SZw2
UYKKGtrMgVlLGOhyjhKgdPCGoWFgCnSgxhL4TxEar7FGVEt4wdqhr1ZP6S1p3DEQimO1OOkn5LJ5
Pi13IOdT5DHzN4YglA76edUqmhphDafnFya9awwbyAfX+Quy0y/C4pJfg5nZxG/Oe90Iq5R5q0qR
vXpXqFsw5im1ctNimeAIGGS7YxN5DNsYNeotAcEGEAEsy+m4cPAPqr1V6EmqTnuAJKyc4x81eSex
PuYE+cnlVQiBgm0RObEMuIo04aYX+IA0Y97ubs9E/jHoIEsUIgQg+QEd0MohmMY2Bw+Zn+Onr+nS
uJj3nxwnwKB3sLbvMNPJthpQ4LEJ84J9mSTqd4tmsJydwI337q/vHh+TffXHbQXP5CJLVvezzk8F
ubrHjFVIy3QGEjp8aNg4oFXtK3DelHAein+9D5XlGj8xlhvk/JfnKQXppSuKkOEktvHpGZsX3+X3
HMOKapaqk2s8x/zFfAkZCLC46l3pHY+3pj8QDGXfiRKZ9aL9IleBwxiKyjxKAU5sK9Es3RDGYt/r
RsLLDn+ey0ELLjFJLKYhVCHd4SswL4BN7F0e7efyRvl97MJGUXGr2KFPEf7WbyDi+gqckDkOnZIS
cWLalCJz5/ESRrrKLQ/NEure9Z3w74UHBh0pp7aATKGaR3HNcGgwMiy2nSaOkn6O3DFebvpzPjxF
zbkl0Yt1eAyt1jI55XfVNp1xuNk8MC3HVHu2wm2gxs9vOqFnzphOnQD3h2j2eYJuBeYKgec3kgUb
ooFT0/ftqsZPCToQnNO0TLrK+tIM5pbeZzj+CHmB28kvTz1oIKwMJ7DJOo/45IgVAbeFeoS37w/6
10yJNxjJ9R6Y3vkSsogkc+p8YX+JtsMAVbiZVyJEz/k9BqU3gE/CkjYlmYCLRGICMdVctE9ekxCV
TpTwwKu4KJAfZitsEBgBuoM4wclA9wM6UBuEs+SvyyQMAbVEy2TINy4IPLnFc3FfUuoGRcc8eyOG
sQbawV225ipNH02BoB3dZF7rJWHEB4QHft7t4GHbPS8JFiR7HTRuWUqIeUhduOxnrQVwYG9KNtTH
t4YskqR4QJPFfMijLPlrwSOzCno4mjLp2rQsjm+q0IEzNfzpHZqHUleV8GtYcv6FiFomZT/pXn7Q
HpftD+SuPOWYYAuABTNkNmCxkYMPSVmkowSPYxHuOzUmiVsPQBy6bg24nzUwnFTdBFagezk3T3wC
DJrtJCF88WJ9JCZuyNnAUjs+AsoWFcS84tYm3xg5/v5/TD2EGrJ7IxXTowWV7BZ0HYyAEroX/Vwo
xwsEoewMzV0SijHC0B1Uq/LEPGgehuDaUlaK4NvI1bkmHF5tFV9riVonnxtmqIPz51lNuo1mHoaZ
RjzdGaDgFywocoG/0NxEbhaqAkrzYu1v5gzBgxV5zmiYMTcmAb53hHksNmmxYKNuZXYEVemE3uXI
L8kXWDCG2O0/w7wW5Quf5dAU1YrHPdphk1A0KNnopeR7pIze88T4PjDINii5ScyHlqNizf9vlIP6
AiYbdZ0aO5/smxpldTQxbxkyMVHjfXy/4Is4lPGFO6+zUgrQwBmTdZqs3MDXZxwfhEuG8zJw7mkv
hNhKEMS0BMFlbI5gBP0ACjpGGQYY/b9zNcXM2wtiGPweZKrk0UmiXVdGqCHM7H7gbr3jglpnu6ds
ltgDX8uQE3ZARAGSVr4CsOAkAR58zpnmuFDVlwRuY6C23TuVSZmttvF58E3YcCDNHn9/6bPgm9p7
NsxGW8F7We3EGIMIw8gdU62e+wXYpJ0sFT3ounjrWDXqc1BLGzrr7GdiMceh2LDb8JK06Mtgk/Nc
M6Vwx9xQin18guMBA0gEoITSOYMzRYAfPXo1KzpnwgCddcebhYfowW1NZ/+jvnMAkU/8usc4f5rQ
FMO3GEvujm6jlXfuG/H/vLlcFMdIgri1ceO1G82zDLxg8bO5lh3pe97vSbcB5wCD5AF4WsYMLjaJ
9k0CTFkpBL1L91bo1LQk3b2CsQ+XX84gEa6ARiP7rRM4UyOzM4C+ZlfDPDZOJG8k1w9JPval3kx1
QP966pcvNLJ0KwOI9dXOcaRLqT+RrPw7++/6qFW3fek+ZuE9MVsgfs/ugxyPBMcyLvGbeD0E5D3f
sUQAECXhzIX252jzETHIYXcd24O5/WYmWS5EdC0RSc4MWjSrJnr1Q4BoLQ7BhVdGe3KCCiwut+TU
V6HgFtmSPFuQzTKPnmzb7sAzbQHzC2XTV9xZEYEM0Z9Ly81T6vL6sLv2gCMlESXXG8NITgTjrnSJ
7s3nEM8GsgFvuwI7hIMtFcCsSPwa+coNufVJhaL6Ezw1kMMPzEI5rd6WbLxEVEQrUWRgBpoB6Us/
vxDXMN6kV0mv9YSdmcceLgc0wWBzaf8Vtre9hv0YQmJZI4fhGUiaa5vIP+obSCMQq4pFPdHaAQuj
rGJQb9Q6hC7odvq6V1iyN6rkivzYAgwD9K1+eFQLzSKzOo8K6flz4GOkz5wa4LGSCa8eLGH0cCRZ
WodA8sSv4RP9UKWyfKEW/oqGjTFQGJe1HVpgUzR2QQgdQMS7Kb+ABzQgFyATfBtbxZTU6LHVqJub
CJ+MjrgqaPI6qKl7OVa0IG2BkoKbFpR43FM44LR8P6iq5ZJK7B9D5nc6yfeswbofeOe75+V3sv2j
n/EukpZ5pcn3JId7NGXD/PtrrF2fbMex3SJEfFgStzg5leZZBgZ3gvIVFg0htpjaPR2tDRIx6YUJ
zQltxVGsk+CwEatFv9rkxE9qBIMrGIdCgYdwghZ36W39v6PMtqybV1cK9u03Z69o8mKCgUzLZT0e
/LB2zKhivz60mYjjW2AG9xVV/h6pBFAweBPdskNTGGAnk+8azUaN1wkC9w2ziM80GVB6szDXkveA
lM6mqV1nriXmwPkUiaGOV3aPmUvWFYwsbNo7Q8SWli6SavbhQWE+DWmMonvwuPgrNBetCKxvc6W5
uAWczWeQrn+gqVCyn+EW3EbNIfWw6+UupCMMAVcAeMR2spo4FQyCGFryQ+6qQwZ0PQtqUqwk3JVq
0Fk+UFL4fSQxKsfD46dLsd5XUlOn8dY0s/UYTvgqXSZt0gtWNdA+j67hEWV0V4ueRDa6z/0/bvSK
N6JSXZakUCgaXAVG8v3zjdmQ1YHQmW8RGDCAJsx+KFyiaKMQcKqHClxzZD0j9T15LTrHbUM7ov1m
4jjfQX1FnfeDwmMQKkSAr62RaFvgMiHuu3MEbzjMMHDklwAS6jJKiX++C1ZHLYdBztbGhyCDeMnr
0khIxWKvQvIHh6gBh1Hk3Am4r0072eBL8cUjmiAGq596ITgkjJ4fMbUjPsvpqGpGt+f+4qMdeUg1
+7Iyn3FGD76vdMu/4CtSQ6sepLIWR2kKs1UYam2S77lO4TokOhQB9bwg1BdzceiQC+N6piOg4aXn
PuP7M3sVLnDhl1IwYMESEgKuz17K3WRymSuaBotIW9IGmEVy2sALYvaabS/+KvKtmfqJ0v2Zb9mK
5YRKlwhJmEvrscJi0sW9YPUx85aw+IoL5/pGlnmmaDl9iOgqdYWxbceAVjeavkoYbBXuGmXn76Rc
V08T/aEDm450pimwj3rdTUqyeNnt9fVylG4KQO0y8ncfs4QPftS0bxTPEAagD9G40di9VfAN1Ly+
lGboDz8NfRX7ddyQeCeL5KfyAIqw8kH8QGyjbX6gjIATKBuYBLxE+RHZf6O9KIzzxyvxWLdVafYi
Upw3XtVI9xNjbDuhbnSeMJl50fESyINuhOtdzdPbzdo9XKUFelybGq+6mXBX+XuYjhA2qeqqktyO
MyO3HagyeAoJsRn0T4m0MS9ACLr9uUrLdoC3bhsv0Dl+LK2yoRMQCF0jy5mr7/xPAnJK3TCkkDg8
2uqmwqs4uB4z3u1itQbwy0WiDARWzQpxThG9wOSZecmK57XwH9BPzQED3sWIpkjwEL1k1YsJMGj0
Km++lxd7SbGMGWg2WfLmR/WXGJSbA9Y/EfuZci+7eB1VkHpzgT7aJP/RkwS7kY+vtE4p0mNA/nE4
dyE8abYpEMQf8a+eYRxuwkWjtGmy+vIAyx1dRtZyTOsUXHdV1cVI71f2tx89WG2Fqlcx+dtYpDS/
ncHqFgDc+l9+vewcN3jdeTw/wxblhNprzLbTuyR4kF1/IKzCp5PwkPa53OhxYVcxHrKntP76FdQo
f4IyN73c9H2+MTjdLHPfS562RXqCvA1p2exaJrEFSpsSYzlhYtvHUJcHnpRs3og/QZo6Bs9Gub2w
QFPI80d1k9oxyEYki40bKTGIOLBeNerfNxaw0wBZbo64bEYNxvPaY0zaQbN9ZgJP/iYI4itBwf8u
M1dKloCaRQ+glwGCRY9Z/v2zxVKZmTwS7UmLU8OhbBt4GXtXDjzyCUB2LxOeFnEn3AeNDhQVKpEt
FED7YYIpwjmV5G7xiejjWXqWo7x6seX+FSL7kwUwKhvgpidHy2IXqhdecnJlhVxMR+qPbblXQ7qt
UC+024CifP3csQiodn+qq8XRyR2EkKBSjvHWsXBAc2ORJ5d2FCLAdVRruEn2We66rJlwvKS+CAKj
XgCseqVBMTrCeekLh1Vzk8cm/lZJnzsiMP4yYEDZPnaH304xdOeCq1DFv3inE3q5VloBko+Pdb9Z
Fg5gQDbTnr/5pPyg98QsYsfE+ZZF34jgUennQ1YAV6RVZg/eiFHuAYDCCoORokdgPfUDEyhnBGjS
Wmc4irzBlsM8AowuVwKhrtQXQwivDpJCRUxGPQCKcQ+jJaa6GVoN4hsMrzv5GZ366zm5D+JTDLQn
Wx7vCA7Oeg0LbcdcczOoLShwCb8hOzcHqT35MjOfQAxN7PMAZLrOHT+BgIsmlAFi5nbCv5whTbCG
Rd3aIUkBxxbY8po9270JLSrfjPCA3c5ooRMY3wb7/DYLv2gjHBj9XRKtG0e+S/o6L0+yHi6XpAcs
EUGn53fXsWVoivqVN3+L4m96xz1Kj6ooI5Ra1JZV+itrIfMHJ2eDKZxzuJp4p1sXZpO2DNq25en4
Xk2E3du0wysY6zKqBCc6owfo/IlQupXbrwWEYfSKS3bdpHHx2ZmFpuZwx2ObS2CpkiOLKkSvzqLc
Af7oKVNAATEbf6TRmWUykN9kTGhhko+e5I6wJN2ExmmN7mXLipIJ2qrWpqPTSI7Sn5Pf4jvsWPh+
aYABrhbbGEHEASt5DK1YkhWAFLPx9LWRWEq4mbzhJZ5QUUbyQIhv6k0y44PUsfatAAn9LHD0Ar4Z
BptoiSzsvhFK3v88Fi5/pq7WR9ojbemKNoaaEYX8DKlZn6qNo+H3DWCOWtrHkZJXOVDefRIm64Sk
HOMl0ewoDMWEg2ytH52J3wbFltylAE+3QRLHuOMDEQLVLpekER/UEx3TCvt3sqzZDt3psB2I7sKn
WxkxEeoPViT70rT7CXg9K+/N65mjjlYed5uAuPJ067Mq4/SYssafFcBUM4dIbFS/BPDZGbb0Brs7
UTrhmwLG1zaZvifjtoJPBgyd/N3CA4pwKiPj41xPHWaUw690lS8GAEXfAMviiTDiV+f++Wx0MbSz
0z3oN1XdjMzLCUja3vhirYPSC8Q6PEifg3DS4oK7EbMK124JCJvMoGqeb5Ty22iqjm8AyGSKI51R
j+PMyYFaDNcxG9lSjme+mLMNqZn2glZHGO0Y8HoNRStFrBSKHJsBXuSOZ3hSk5OGyKIQt8/9x2B7
q1frQsAsTOnXUgHPTK85d62iMlgFrac6UVkseSga9OiIbE1HJOmb0SvKzNBzdJPGxe0odhqJ5X6q
8gMeV4SdbAjp9UbpIaMKEjpZiyCNOGkm4xXFLLjERAPrga1UnS0vqx/OuAbWK+3fjrbqXNU+0Pph
7aRgVpqlmbriExIjEn+AG+YJZVSekDieOL/l94vPBBLsJCID0Xu63IwFt8HHiDkYXSZs74RShgVR
P/doS8PytPGTrOyQndAJo+4QZX+b+B4tgKIIjltfocAip2PxjurGkwUxK1+XQ9iPelHR1EGoQ9HM
Gt6PCvsBb7aaW5gR4xQc9aioGD04roh+BiXdGXdNXSY8RCp82GmBHHoOlegU4bXfcG8xiX6q1Ern
EMkkvJFrKkq0c7Hy0SVxcwu29J6/f/V4TZI+SuybQCPry+mgWA6AqD8fPZYOixPchMYFgrze27sa
3Kn43gu5Ety40LJCA09wfMQKpvJUVgMh102bxzc1gqjUnlIGYJwkcOd3C1ffaMidFMDgPqxNJW9U
p5UELzGFaufofKeOUVmoVbg1B4oWdRzKM7op7s9ZugL29UtQ7NgYNiI3K0h1cePR5hwURotl3JBv
Gcl9BHAzWXnRv+buBVFEaudh2XnCbBW3MmridRuYm99vSp/Ysv/8FYbAd81OsPSL050WQ7ZJm+Oq
LoJ6NUf/VV5mgaqRCDU8qYK3eRQM4KrJNkVKtfFvq7K4pS+ItLQ241L/O2aSjNCXEwRTWubKEt8t
9X7SeVG5HsV/Q/YaVwaApwQWEQn7jZy1LZjJOaklef9LFVIGT/T2m8rWXTeAX4b58NwEJP5N1Ssv
KdpLm+Vr2+FaPX+wQXruCm4x48nf3v5wsG3o8FuZsv16DjSdMvPyhzCrIufvmnHJF1/1Jc/MLGd7
hUaHF/tcU8HA4qAnmB72VVzIHer+ZbImwZUmGF9WoE0NTfpXWGusMmpVwM97ObqJSbo13N53d0Fu
fNQkUvrpZmKwVKFI+2EX3q0zRKkEO3AW5w6ZA7ExDVMOjDJDbdeUH8JrmV0n8WajbPtF9aDeXZtn
cikRVpFY9WdqV/kEp7ycHvTAkk9LsFxGEhyG3Q6oeQWgnKPioSkEH3w7rWrpadzTXJTGUfVQj4ui
c26qhPVbYdiLd9W5CZ2STw0QG1HhcCMv2grD2NbHHPtYJtR/jeZeJbHLA6Ul6ksDmG4S9C3q9XNX
w5msTfp+G/uqNOhuteifeKOU0OJCi+VZYVjEny1zx7g/RShIuOl+/SrYyNbrOP7C8dHcd9sGcHom
INyY+TwmEJOr4v4/39ZF7CjSXTZ5NmTHl1J6LFewc4SSeBLPHBaDMCMm4hevyZi3oDyRk60tLIAQ
4H6BgeZrxnrEpG/X7hDOMjws8X3oMhlpOVdlCxduZ+UXyvqLyQvhhFnUQJYy4kcQ9Pio0nLl5j1l
AS8y35AoYrnN5TQq6/Ehfg7GLi6Z77sqkRsjOZBfjw3ZO97ZoJYntUg21wHNoqdNDKovcdMhBEmH
pHEOlKeHvyXs5C7rH36cpfG+q3gd9XN/5lRH6e/EU8Weq4HbLgI/ndwrbICO1JueMdOjicRH7Am6
nIZXEMf/LvqcN/S41tqYKKgySq+b4xIWCm5CVjwWLgz3SqbMXVhg4X14wz7kPczTllXPsdhHdE2v
yDrc1hNCtGP31by1U8A8XM6Pqe/J2eaWCPHOLspIQPZczXQ4LwlC88aWbYUVZFuBSE9SYIVOujIq
afuMR972wPmBw924vROpnkgiqpJvcfLO1RPyevycsLgzERKMkmJAdmABTVNXkPZdBgCMklHI98Jf
H0yXhIWgBr69d/Fk8kG9tOOip3G6q7X5rL7xheoWUcEYeIa5VtEg+FPIi8VAvgrYR36/dGHvLWpz
TVPBIsLcUrDpDx2TxD7m3ZNEFCtuHW/DUqVLr6bRDE3DSszNk5gDoBxxplGMh+aVW256kjZrTz+0
JTCmlUGSgE/keJ/+Rld4KUfKA4Xrt+dDxn2OizxDi+AnxJoPplDPj0UeKu43DpN/NWckMlEPETKc
na91E3V0xDikMrgnUGoJ+6+a77n3h/1zAPLb2MxEm91Cb2dxXncuFyD40CLGf/S8qGQtvPu4YGo3
PJtoQ4+b4kFGO/a9j2ZOoSE3z1aE8IGox/NWWvjcxnrTqb3HDr40exe/Yk6DR7rePsvWY+paDH1j
E97h7RdvRuwI2shaENSEIULDduJNu4ZVoiLgNtT/154EEH1qHgvxy4llycLeSx/SrE4sgxahWDj/
cF009VUgX5J9sF1wMcbAa7dU+fV76sd0Efq+ysyA/8LxkCmvdQMmPqlSKcAzjuIj1lYKW9yxOfJH
+fNSmcbNeU3RbSzNswSXPmr15Zypu8Q0Ea0HmAvR9k+7k5dxNlDArwCOiLz6RY5e5WWw4Qyq5POh
adj48gWBUkKuYJiaxyNlZc3Pgfk2kAhRaHLOpLpmUbLkD01lUTFUZzzRw2UepmPGgt3srU9X8FgR
RI0TNvOF/iYX2AvwXRQMHVzCzoC0Ifbjxj5D3eUOEXZMOeGxFAkkv/u8XmxaOwdsjcoL8vlEgl0J
KdpOSEIRg0//ljt8jkIT4l0qa8obey/xFJHOJ1n1SHtHF8ac2zLnn0iGmxYdwEJp4dPO9LdYkYUR
zG+BF0KR1l1Wvhtyr9LbAZqCQ/mhugwSD1zNmWd9DedM0FRf6lkHszrIh4RZ3TmVp7uoi4hu1+V+
CutTHzoPDb10hzAWq1amkfR62RA7JohuRiU792gXYYIkxI/mTsGriofS5yqmZ/JlVwj2scYDRntt
U2D4iBFC1BkK3FHe9afiPYbqJspa9zd9kBFRo85oTdixrPlihS9FzEEKmy5GRnveEFXwEVgf162O
u5+VTc52Cb0wiG5Qqy2ZOGaRKzQXk40PJFkWRmZR2qeprQKyq/uFGQ9p/r5oMktCPpq+mSEqFxYB
PZTK9bKFwspRHtsJ08wZglEoQQ88CE6bNygYwNo1lrKBQWVHKOEReQV/ve8LlCxzBj63OlfknKq5
D3imBgvc/r7Q8+/V/lhPVYIcL9l8Lxz5ZCXilxmPsC2aD7e76VO5GXtOW6wkwPUQD9zKeZyrfSAu
oDO+djUTAY04/+B5mdC/fZn6GTm7tybOUSu1ktsbs512eO6aZ0aSbqAYVgxVBG0ZVVmdzTzaWb+X
iDbf0wCFZNmqCb8Ni5OkF/9clsDyvrksYUwscTNKLFn5Mz0fwSoJ/dyws0IgZUn6f6dUvEj9Y4ev
ihNyaHsgPFCbXbisCFuly+vla9pUwfRXl7Dd4gGPSiGA0o+SHiV0KLEboJ0DMQC35nC3fwWhnpGB
HlDUqHyJh2HJzlUI9us4Z6BxbaxGQB1hCsbSnu2JFm3J/UK1v7epjkXf3lIECg4qmnfDilc+JmSj
Mxpsx18sTKXH6ZRUgjR9magrHGaLgpYmbBcKxn0RAcDM61NA1GjVm88+25b9uxrgb8zrVtidAgBH
xNSuHB3vaNBSRLc0g5PQxdiy1OoCBfmrL0IaCszVbbQIIb18HfYAzDXfaTgdaSR1yqWHrjuVS9bi
cEfRUXBSc8a5KGZ9hNHmj6gjMPpJFkRcTsZ6qunFTsrPyRcykLG7yc1GbLRRswlhToJgeJtjaF8U
meswDsVSsx1I+ZckJmENwVVuTLOqgWwDS0uC2+GiNuTBVOyuz4uyWdi28hPHf42++bOg4mPK8m0R
wdYCWvs1ImKgYUvlzfhWSX0tCo48FsLEwDVpbD4lma6x0TIaHBqPqZYqDizjctRrG/zTUJLOoLUb
qSa86gbz4yugELIW+90qqYb4IyRyLJNQl3UcsbHCJ3qUmc6Nz7QAbj2x5yhPFVMlCJv3bJF/JNHy
PRqzmb+PTh+xlMAozKiYKu7GdVcqvAHM3i9k8r1NDPw46OmcySv/4KOII3Tw+nWh3NaJkWB9RATY
5ed/zLtKoy4WyVrJNaNTFyeYFkEWlqyGD4kFFoOJRapFjFsERnspT839FD3ezCvgNJ0JMKfdB8hk
Vu9rp7VhHKBi7dFJwpP6mGGruXXPyyaOhEF25pmz/+k8lhCedj4nfFSwpe7G/Eu8ei4RqTsAqPhe
2Jr2EsBpl0D7zrff3lIKrkh2Am8Nr8xaSvWYn+6TLiKmHFm9U9kNb1dctrtjufiPD1bGGR4UjmVO
0REv/WMYbwOyEnB9FVeUfkWG4zC+kB9z/UHMREJxwyGo4vqvfUlNXEuI0wSS9s/uZk3tWN+WyKYi
70taDu/BpzYXZ9UIFzjeNCVZhQHXEKtv/eN87MVLOc9hI1PGACbUvZmMB9dZJCxqY7kHRjFVn3d4
eEs2GMEm3J5tbLG2LR6jh0Mj3z0KOlfiy+CuQ7R7usURyPFGnzxtTyz5TDyt+gqZHw/xFM+GiFPK
0mw7FU/zc5CsMCSH9v5Iw6YzrgYG4SiCLtyybqV0N/LZTQFbUwafEHZn3z0UNIZjm6uruYMy1ja5
BIC4g1+dPkIybblcA73We91KWWkhos6Uz26RqLoQmA3hkrlybT/jhdeLkywIFI4R/zbL9vmpPbJ3
nXnU8wN9x2KEcQc8FNE9cbnBOgXB15in/9IXysAaQgeUgpEK3MMI0OW6Kw/FswcYQ+pL8XTL86G1
uh26s1Np3Gc62Njl0XS//YGO0LD0OZHtVQU4hfMDJ9bvOiSrk+PwW0hzwtB0L7QvvY4WhXvrmXpK
+e6P8//FhVRoKETm1+uOpDFH12wXWyT7t0HR+G5jTlmTN1IaK23drgcD/Std1mQ+JkSYCBHyBdwN
TlaONe4iqWJzGx6PaTNZYjpA6cSuVuslGIX7nCbRdRAVz9VBFy20nrnN1IQ42e82IYeqgL4NuALk
YVs9Tv/FT3MoIMjrcfAc0kqA8vmuUQ0ubrW0EWS+efHHB1I5A6+AVXZ85R/KM2GjIRzuPiLV819O
Xhh0kEatlMIMe0nVyYbcSQByh1y7lw9EmMwNCuyGNW6HoUJy44l+czHIS5ju7IN+bRsoRrP44nKR
0wUuXbKBCdMptuAZVs8X0W63qE9BXFTIR/g/oyvKiIaeOUDqIvKsnpCZ2VpsRVFZHulBgLTcejCB
Xg5uyId3On5ocqzMplMJlFa0r947kNCVcIbBE3yNm7XvznDzVHXxW3z3GaiIWbLNfAz1+vTX1xA7
ofkkLauN1mAPSIwyCclh0csy33sQJ8vkllJ77MpXaBsGdWOkooOWM97vm2uHSP4lWOxkAlULXjJ1
0GjK0u6iywlFDRq/rVjyg/sBzS9OKVrAcWpX8sQ+IRUcSACB0J4bRWkgmw7vsrge6OiijGiuwbHh
aKBkZz0a+eNHkWT8SEItk8IC2VhXYLjO9/Jc9dWhgtfbtKV7/eUB9k20eGSUf4/4r6znYPVTPXxX
OtdRkbfqwkzwDSo8LoJEczZEp2Zib2Gw4yhIx30CW9c/ni3DAQ9kLu1yzxcFuKAWoRAYwlSkwWNj
GU0fVLNYk0dzUKkCozIdhgSoaosba+s5tcm53TUKjJU3qTPb6V2VMzL/aTOAi6PcEeOK27lQX63s
pCHtQcpy8HQD5/zn96gP7PsQsK2WiSif8w0GXi+ZieRXaLkF/aD7bsSgq2LFyu4fk3oUO1nRHnLD
1goSl+JGrSnrVhhmUImaOj2qsT1e/nWUUTwSYPSXT94ksH6BxpzOaA54+CcHE0E98CW1hLuyxhKN
i4W9D2UzGZSm2uGGjVjtySzNRH1Zw6FwR/MEGJUL24fV4Ge9lArAcnAJB1Hpu87vOh1mEZUABfrs
Fh2XVDwPGMtAJOU8hTsF1Yim1RB+a5h24R9QN7zpRhytxkBmVAyLCBD6tWJeNs0GhxazCeIqdTZP
ZJau4ei57vBDtnjnd/+9/As1ZudT7JxUqyc+0CvoS/Qcrw6exLvSROEx1xzbVHFbh0Q9CO26MKBh
Eev+e1IYjDQ9AaFMcGPvwTmOGd8AV9c9NpA2vJvj6d/lurMd+0CnwQ/uyuqSmw0PMZs4EnKWmbAX
Hs+++LG4Gxu2R7qqbCpO3YcZE+xUll3TNGMw8CQjsb70Le9FU0qR5275uujZ2x5M5fdQAgv+nSCk
FniMrDL8URU4RA9QsCdW16fW/HclQooD+406ZYY2nI/XIHzDZtU3xOpqkbr2z5U3txGSKkymyf/1
I5elZibAafb/LRh1mVImE2GiaBd5kjhA/a/UUiiToP1kMEgA0kjqkCSeuO6530JJQW7B7XYBvCbN
bMBTMiVMjnZNs2F84uVUdXiETsvMsbK+fSgOGDuUoVeyy4MR4Irru13WTub1a7IEhqF4wK7zIg56
fysVOHfvchGRaKzI6IGOqHf8I2TNLkHslJj08tfET2JDD+DGPZzmJWnfHPFF7ROQJjn3u8hOLuID
tT7AKOkA/BS8LC7PDf7cRIHtTQHKq9f9Hhb03s7F7Ltxx0Bdb0lnXEgvvU8b1MLZeLv5hFeiB/Z0
pIh3q1ZCJleBwGEwU0OiltrhpFCYuVNrLuXPXhQdffcs7NjP6Oh4zFmUIYQ7uRM1B3bB3GZbQ6f4
QQSmyHIIm5ZDGzqW+dgyLaxwdp5XG6ZxRaUVYO1ms5L8ys1EqsxBvcK17TA0vPZZ4MkLRamTsrVz
GiWMKT04W4QDPgeB1S8336nYgmcMjRmC8DnaqNb2OZc7th17UmOu/5yPCx7Dbbr0fg3woKen1uRw
h32CS49SYFauGNeFYB4chhZckq4FYoSb/X0IwGZ8sUA+owcnoS8VKJXa94XqEg3JbJqxyUw4vp3o
QGXOL44yoejjVlItREevLACvC8uuCX3J5cppbn7V13GnYr7fsJSoPK1SuWg9nkQ833+rUVCHDUr5
g83Hcxg61lUX4JWusMiLbNMc4pOs0BaCxWZ27j51VOGMGeuZP/DRxrTMabxmyk5M/MrJImzckAUt
pCXrgfnAaiyFOmOPGRYgMDEw+UVfDnIKVyJJWIAtR+6pAjXwdZrhrPCUWbUnI+XOTcaVCLY7b4on
2NFF+m98FJrLohhhJtSUlY9NEmb8CcYOMRsO7pJvvfV2FkyGQSplqgXdFcyTxHRUqVJGHyUGETUo
Zppem/ASiEphQWs5DHZNfL/MJf+GnOrFXMfAFWN3si3z3w0Q/MODm80CQvC7GqmU5TNIMTdQXbTW
ueUz8iT+/Yg4rEyEzNfhOuJtUnoMeqkjlWKyvLgY3fajDrqBqjJ2sFlVEsnKxWPLsU1kNBSGM5IW
hOkQNTygCORRFRd7zS7ld5NQ//6lp9eyd4qLKBUXdkVDiA7erzJ9dNPYV3pOy8d6zr0EohayJVmt
HhGw9elwGiQXy8WU7HWGOglVH9q4KoeDHvETOIjgLARlvBlPsn2IgbwAOfIYWwe/DlVqHXWRIhlo
b7H+X3pPLuw/Wk2S2wfLpWqz/xJQnaCig2/5RYvGk6o3MKofs5mH2YBGI81FP8qACBK7bl6QS0B2
sbm7YI0haB1t+EbV2hWvmWUMqG2aiXN/kKiR2bDCGpgyfDiQrp9nSqPwNGsPZbNlfzw3BkNZwBap
y0C7m8b2ydfiZd6uWoHi1kbwGxgqpOXWlDupUCwZll30kJPqMVGeMuOoyc76dL+B/r2Z+CRM8640
d/w7qdJSURc9tBRbc89ji7P3iV8DWtTNC4N06UyIA/I/oIxU4iKn3ce40sBgJfFRKwznZP/UIHOy
DUTclwLS7Zgqgx4eo/qhss9sx01aN/0qUDk3nQdtpEqiKjBabciHtR89DDvtLVEK9eJFGMGfQOFO
cLFpu/jPhDM+BSD21TTYdfUmABOkC3OmmxdCtwdYwkIvyx2ZDwxfVnvp00bV93VXrSYTdtsp8vf0
U/QvZ04h6Ud9WhWkFKT6VFoCW0rf0Bdsx98CMhFojsdqi8X5EjGjHT4oE/iUBqRnZQ3OSrsU8PWC
+IxDwhCdfNcpolk+S4/j1+FelO2Wfyp9P9j3HHlqkatSG3TTysYxdLth8svP/tzF0lxvVGw8Pm7u
CRYPMRHZ8NQzerSA8Z4sJsXIH1LmsfQl9fRY0n7YTkBBECEiEN3wqE3GBzUbGRm+jbo5yxdX1E2O
ixYp3v+jk/KSFn75ItopGrRlTFiZzjy9GjhUGdaoEih/rl1aFb/RaDCRD4zizBpscbsIOEiQDM97
T1JXkPtFi12qiWMANMirbz983UH7yNj5cdpO/q/PncwBqrAPTXU7B/u4Epkx7YtgvZ91o6VzONkx
jcRpV/nlc6hApZh4ybx8UoiOL1VqhaZb4mJtfpwbzXHnBXLKluEStfA/lU2eV/Umt32n732fwTnv
bZH6wlyAA01i1CkjO/t4MkAGdOtwE41J+/jwYAmd4EU3k5gCuh0dWH/s9/IVgjvMWVmQJVnieLTD
XlLxraoCOOdLUnFRL7ahcLkSmEV126QzrV/eCNpML44QtOUfp30krs283k0oIxdpmyAQVCAWcB6T
kO8jessVznN8fWFhEH50vR2Y9/zzpiOg8sxJ9szRVjs25HpTk+3WsPR9zRnwERJRTKP+cpCupgl8
HyHEkHqSVi8loyK+EPUXgHvHsCAYrvDhHLuUdAx3NRlubGXUa4ZRah//1j2Gtvc9W4PytdByZSq8
yDKmsyZ7SSC3whrt4XYUQgeMf7pR7GoFagyb8W9M2ZKrsuuUWQwXMuojPjPl95rrgVthubJd007o
8MNhp3QBJzoxI6yenqyRRDPstTWc2fnHAA2GdQzyQ5NXccldM4dIEGduVStF5lIIFWL2v+O0zKSk
EFabFuL9XdpASYCr+nH3+40JAbuOBFrlheJ9NX4xxQw6Uj/lE+4dcotLWhGletJOz4OAIj/F6h49
iP3uBpj7RmRMNAmfclZ8xAR0x8Fa/Rz7UOiwsKeH4ziRGOh7t1gnzAv5ytIbErxW7hUDtFNZRl2c
KbGsvzrfT7JRL7H1toqhhYGxqBdH2vfL6ASIdG3Wf8QwF2TRr05EnZm6vtpkhv/3FWBumNUhLMR8
qaKtjR4i5PVH9O9/i75lF0+ekZ33PzBDdNAim12pkBatwl7y0srG2apyLemsJdXEYmFa13LcrPNl
TAzPtj+1wBInpBX30Fu79LWkgzwx4J1bi2f7ixMDGZzgf6G5cZtMXgGGSHHCvHg3Pt8ADpIM2FtT
3sjyd2x6sV+3+N+MAH2rOEXjrC26c5Aegk2z6mEf+enn+p7Md4jkscnDJE6n3OC6G1lFa5uHvQH3
1k8ApfPKWCaDARoOlXcuQZ1g2BRF7ixHbIqdXe3YPjBRJ9ACqY06W+hJxSjgLs5mdkbdrPnsMnif
N0FJVLBcdW/vQvfqBNgSqtxTog0ZAd912K/6DNf7Uqqe413WfAXncc2DhUOi1x0spy0lrKtOuBq9
ddbvt1qkcTct3mI7fCwm2FlcwyLS4OGHORH/1zOesOE2StaO5KqirTI44fgoeMIAAps3uESuiQ4H
iivSfq9PbQ6k6Y8ATLfTQ7XJv/iOaokDoz6yYC+bj9wnXXXjDXmmDhRnyCBppseUbNZbBBL66Lvm
UeQsJjY0UdF80w3iY9p2BzOD0dxCk7x0z4CZG0oGYkjJT+10UFqozLqzXhY4hERnR13SoZN5/g8w
gCW3eL3K8mSAUX7yazPh7KnbKYDYzeaB+Ta02gBeEE3TNgZut6SUGaLCG/EvHhZPq4OzOLgpNF9c
2c5jJjtoh5M/RqdVwB1Md8iwDcaImr2UdtGWaD0z0CAlylOqJieCITEzX8Qh7xehcGI9POGRG6Fk
ooKx68FGrKWnmJ+ctA7PIGhC0J+9N6WJipRDUxfHqCeb0kjtAsbXdsocK0eROBhYIPPYFgRGHS2T
wW/8Z7mgR7sVpiPp7kjiEZfDy3GgPDfDukwi9Jiv0KGiWZWtSxax9goQAbsnaAQA0ytAL4P72lyx
BGzjhrUJcrUn2k2Fll2R1bMOxyVxe8lIuxW2JzdXICk9rR+twrhZ+rLrqWYWdcksjq/ruGfO1WjI
zb0njqKzuCZHYWny2/Z4OwrrJme7sAmsgqpCqUl9qAXKnaWiD4bp9F9c7I8mrnxWnY96W5+RZ0Bv
a4scRW0jz52815rT7sQmST8o2HqLtWecY79tily+EFLOg9sou7MUQClhL/KlD3Adx/g1d0UQ4S5I
MfyPXmL2op80l2hZglh4XRS2qz4AGHyRLZ+n7Cx483VoTU04S2UX4EntLKYhBAmAkRVrFRBGS8Aw
V7PM020ZYzgtTA0QVfolhpiPCDWTWXcgwpNWl9N4mF03850e+Z+/RIrJLO8TsGghMVrBHBRmkhYc
4ewoALF+IeXWWcLoEOR6MzVYCytkkXNA1jcfta2NwxK62OHtiCe8W051DXWboXiW+u1C+6UjxRiI
LDTko5Za0PC4f5llGW6IZCqboilanGWtDVe2myDryWGrLkE0csCtwQSgorRwmuRPVyFauxR/jmDP
rvrn3IpIdmR+IIqqOfFlP7p8Y/fg/MLZpyqCD5CqW3oSkc6jtEQeZiOkqy1eQk/gcnQHP4SXV/u6
A+T6bzlJg/vReFYc/cpyWgpkU8yexXSf2o2Og6nb8TQ9DOabGXBIXTh+gYoEdir6n3fzk6buwyUS
iXpsOjopmN6bwER5df7lDo7cyN4zZPZou1vuhUej+PKBXtrAn5Heyyq6IDK7/dFKeEDqmsAj2Evf
kS8JCWemvDTddIIpOwxRZuvc2Qz8ZfFf20asyIZzE3qTP0a41pZEU67vtSTzvmDYszQcytMRuO3w
3vmr7nhQGL/lbAFSfJWFxdeyDzKtX7V8F3fbmujPb+6e1hpIJ93wDtkhmMaZ5xm5mukyEoC5sOc6
WSupyX5xeaEA2rs3uNvPQyVMpuLWSUnE2WCqyGL2uLMlJLwWDqP9B5lVSkTkJvdqtLQc8FHzPzv4
3zV6vorEGorjQ+e0He3XNXwJ6KmoWbtAfwMwl+MwerIIHTlB/FVhxeh/Mg3lAs0FnSfPrQbvPN+u
EQJKX6C58Mi+FsAOyQXDGvFAXzUC99ogZu+8O/+21lWxqUY8kSul/WiPPpu5VC2LcmyPIc7j8OZq
YkHmaXVf0RIOkvwVZGVXhpQsWRs+AQKOiQB4BADiNApI81z+DRCud9CfgOo7gBQ37NERyVL1esII
1AoZAaooylFV+4JQGBt5sBHWvn93K5Tq4za3Lng+5SwPJVQt9tYE3lkF1QPzKvTOcNZ02Pb0pJBp
76HOPjJQnbjbqF9oSyjFLe9+pXj6uw5MzIwHFyXlD5pRCID6OcDxuPe7XwP1LqDSqQUh1PC9svDj
CwC24qlmy9YEp6zxBTUT13ecyZFGI20e3zPP0K0+0rRui6vbf6QMPnFb2XRCuLHN9tLdQ7046ccP
o2DJEX5IBMSs0R2zZ8sFCLDEB4fhVZHmgqPift697bKBPf8/psnXGceI7v+lGzhbDdzBFrBaOZHZ
bNQbw/YjnVK77rhEEWQpLHv/O+Xoaasb3rVyVYuToDdUBTuzkH0ni86weUjLJPYyAXKKdXt00Dgc
LeYSkqUTZg+rhOhwlMmYolZZa3ya1p77vOlRQwW9T53rby+SYp6cDVyS2+qCw2W+i/uNsQsPYLjU
uKA/mGsTmPyWB2piFf9dmsHeKDBNutwkOVqCkNsDbDEEQz0Bu0WsXKn8SUGJzokHIRwVF+4FDanI
yezrLmkTfV9b3gMJEEqP4ln+xIAleqK0YyYiElu+0NR82FdzM6IuzezI7op+kF5xUrGmIElxhiHR
PGuIY4HBoG/Ju92i5/v46QwRjvjlgJAsHjVjcmoRvi9OfLm7VtbeqErgug+kIwpwOeDrqlxEIMUv
WEfmP2gk6WBCWldxBtI6eYPYHOeE6/tLcyshmW7kkeUVaE7WIQdd61wB11iAeooMjZigw9GtOTBY
zHkbYYs9FIBFqKp+n3Y8VcgEx0TAzrAong28p+UderksRBunha3ALvlvqNsZ2HJ/T+/CDVTYrR2/
Ux9cRwG51P+klqXKkO8iTzrERcgyCT+qllZDfyBhMhKriLMidawocAzLceOXMSQerpKWYh8KRIwJ
6H9H/C+V5wOhbbc6ykrxHwg/sc54W2poPLfuYH+s3KXDffQYJY2mI7vSp6gzJrEhrbrcfk8TkCGl
k76DTbpytxBHfOOYZ45ZEJ//PNkfNeCEs9w4rNtEyxw5bOj6qyyv7IbQgbS7wT9sHDphIu/4GCXT
Woz1Tw07YbS3YOuSAeVyKTzuKPppPOeMzfzjvZ2HlZn5xv7rCQzIVKzRgQ8I9gbYl7Nq+25DtKLq
00MLHKLYq45H3AFm+2LoUToHhdI0rS4Eu7jFc3kHQVfTZh77RX0DZJ2qSijgtBcMe2DbuxbTt3hN
LkgoklKD9S0QMAbC730G/aaJfh/AbstxOMMe7+JwrSwSzbrMc33pXCPjEAMQZiE/jEBKxiw51wr/
mzjOMVIBPNNAmdptJ1wvEIeYeqTGW0Lxb2u7c2sUZIo+ZHhNzqOH76YbYAYJioFyUaDimRtBN7V8
u3QnankJc1glZ6pj9nKtNVEmQBn5XJyrOok8j1lXnNFlSY1iNSbz7doBXkJH44oSq0jKew9QmzYG
rY58zBgRgQ0JY0wTrzEj6P4LXlpHJu4s4NnGpMIUdup2mZ7TjFUCCMizsdMws5JpZnbi0xry2beU
T3N1LdLQCigt9cTiveXNaFzP4byaRodMzwKMMj3Nkzk7TtXhqRSnxVuBeCsxxsuPLdiGktIm+vrm
2BfhDg3Zst0sT4+SNiqVktIKY0/w7CAsJKeP/ALaE1YXEM+1cnlkiRoXRswMhhrTP0M55HoFbi5H
ZgOQB3ToKkv+OiaiEL8Uf1NhNXH+I7IOaLjNpQRZFYMGCoNsD6egBBl7tDVpNy4M1PNri0pfAipS
x7wQTSrQbnhz4fKyWqeI2/osUrbrE0Pz6TdKLyP1iNSru2TY4orvfIl98ZPhBa2pC/ZCdvTSe0cF
hjeQzduZT80c2IRso73/ujlay/EBTLXCOchboJW08xTeyQ4uoU59AQJqHRJL1NyCYOpInXCOX6bS
gewWiFSrwRzpLao6LGkhpFrDSHrD0JhLbxSfMMJpjfIMJFT8PD8CYZf6LIloEpuU7lHyztah4slL
ulwHxveU6mDUw91HlaFT0/RRKbbE2/FdsOS4vlQtzLOYbK7T7T23C2ZEGSbOeOiOpUZj9OmnX9iQ
m8oXd2K/T4Fq1qHrpwH8SeeTe84OopcJVh2TINJKEZ+kvOgsD95DgXW95Jl5JK5wFIkiVOgR+1xC
amGceX9ZLXrjAvtE2Gw5yGE+onLWAsj0Fqsg8q5J59m3MAHOGz6qLKUo/f4WB7AJ4W0rEL0HUe7D
AK/rkXm6F5pWNiSo/yWGpca4LwqxIH4s6Y7GuN3XSIJd7G14ws9ewlfFv7z8fSdT5r1ZxnIdjW+2
8v/sqw/h6unVNabMDLh1CfShB3x/9QTgnezGWjuJPgwfTcNiHLPIMAaAm2hqn/FgkIOgSLZodETC
ebNamH9WcESyD8wwrTybAi/CO2ceeDxu4vEcH77x5Hz4j7tF8eauXYkDq2koRShkpqKumqqxj4Go
1U6fG5xl3q4rLPDwia3H+vg9gXktMREk+x5vXV1J0FapCJlycQKjxqt1YlzaZ7amZ7wyZPp4pZdj
fiSqml0VSkA96xbjJxmGvqQwt+FtResGfFsuiQHdbZY6OqDIfLP1Oi3xZbURyMs5QjVLA5p8Z5cB
sPk+hjYrSCltc6BqLlBW0tzVQN7GOIyygF5QNlUJeGkCYqxf4C1agOtZB6fPDEpub8EvZFTySi3G
RLj4CL9hr6m8KPc3F1S0Fl2heoe1WQ2+ljNYpfeWEsZaC2AkOwOtqxzaKPnFBf7YhesPspPZ/LUu
rTiDz2UKlQR5HIu7Hl3KOef3BwEEI9bye1xsWnkIAvnuYB3r26obo7OtJ6HLrVKSauvApMSvICND
1DG28aGc4e377dX4ixh8S5i2s62PeOmf9RFX8/PrPN2a5bdw4wZv2H94Yj6OOAcP+/m4uf4TvBEs
o5plJHMwgv9xILUlelOUU2a2drFt4SzvmMsRDxlBdfERmoRHy1HjZM2WVDpL75XUJofkA9zuRLim
nfLjO2zFgFNI/M1X1Ejl4j+GDtAsAyv0Npkf3hhvZnY0NSh7TIFk3lBqrB4/Kd2oOBug4UoaolgH
Xxyhc9W2ZZyPy1ySwn4pLw090Q8JlMDGL5wGNGz2mGwKMZMGvx5fnS9oPXDu0F7jMCzAVWMqtGVB
iLEP1aM6frUX/b/ve0r7hHfjncf/EGFxtPH2hPamoKDu1EFbI/jRlSAt+kJj6yo1/skpwNT3QduV
B5Z470GV1OVLEB9twlAOy7m7H+x5UdHeZvb76WYTqBuT5P8WxHX1LX2oPnXdq+bBNlUwZCpCYyPJ
V5M5K41S8Aty8DKABGQJPhqk7c5TKg2W/CXTmZmvxfomzylojPo2s1Kb16WfD17mVlfyfiO7yyZl
/JVG0e/jCujUULFn/TaaufIo6NBod03pLKX16s93R+5+3N9xxgCgfT6GkAUgoOelCEUPa+SZZPrw
SbsxYDoRmkD7OpDBEaKTmBqOOEe1GbZWBtoYSfW2ltCAu99K1qMTE45T9C78c92Wl66OlaBN+ykW
p3eImjB11gXfOUaTZYYycJNUe8eOWJQzfLT0gwFKBOVjZuPGH0iWuAUkFbiT68EDl4MA6J3lktn6
zFOdgv0wJoSpf7fYsT0iiUpVX3o/Ol3N+X/vAG0aQ3rnNTwDQ6nkkYYa8xeZsCrK+15t/3iIpB5Y
rDQl3AAGZ7QLa6XsyGl932p4FnL8kjRA5JYClQ2LKG1rFeAYBGAab8uuNllS4/OwIzKw2ASEp6sh
4BBG8LMuNFMyKXXIUfX0i/w70jfbxcSCQuqvlVn2xr549GUnijdnokdXexcXDLkfoLLtqbwW/R37
lS5CH6A9SVOgvVloKSz0lWhxdDJCfcUjM9e3CcFJt1KjZLH0GRaqgkgjOABHhSYFv6Jq+siJqLQH
+67yXRNOg1yR0eSLjzPi08laIH77ds77qKc1LNqenvVguaGdVpcfEoS/JUgMGAUgCABFtIxy00EB
5iLrZGLzijlz5yQWnJzM4izvAwTGeUb6G3M5SuhFAd4PHST8pSErg+ET0DhWvyDcxaHDiZI1KzXq
rzvpAOWfAvPCb/jY0gJ/pda/LgTscZ7zCRJxnELsVuwh92t78RsPtcZCPUnd7FbJpLy7HjYuGRLg
bPnCLVLmFjbOSW7ZsCvpzjTNlD+6lD+bR0/vnIYwBLRWFzGq2IOr9/DCGZqzzHwa79cCLAbuuGjf
MOiZS3E6X+AH1V5IAFTGmsCfj31HdXI2xwwWEfuzrV10HjHTGy+ZpvDeUHAS5gW5hRIPm9g3SrTc
gotww5enysIDJJInmYo2cj/AyRoCzVg4X2YI19azib73O2eVeqFpGZSkRYegmbUCbm6vcCzg22z3
5thSAsIB7lnJrSe85EpUFGV6mFhHP1t5rnnhxKB8e2lrY5Ysgq35Jvf+xWM2sdhQ8UNvCxPiZrEb
vy7kIQYSCKUDdmUcpIHLtMi6SH3j0+JE4i4r4NCqE1z5S9iL9fCBjS3gTvmb9VypOvgA0tyPgefv
cGGZsBg8mW8Hl3NajhQkzczZP5UbdWBzxtxdJ1QNT8FS4COs2e3OhRg6fFGCe4p8Kg1hyGhDkUA/
FFN0TfVFABldRD2nuNx7ss6ta9CZFnB8xzl6UVKOTkLxX+jufQqlMpaz38alXXSkSUbkgqGvaq+O
8IXnY2MVJY8YpUeK8CJVsd3y1Bxx4PoDnHJxPubhfGINr/dUiPuXaVPAdkWfFLcfyvEXvTmnxDsg
XJ4/BsQc2LKvKPrlbIEOpL+sYBWK61kiux7Q1AUVarnc49rs7JjrVZpn6woil5VZF0HNybjWGimX
WKI5mH7aHueAqu13GO6xC4dZli27dSRKHQU7VEriDjnaw909rjO9IrFl6x7ChUKWQD/tx15dETBf
aXdV1fAAjxXx/JTWA6Lbmj3BIoPVfH/+YDs1fjtgB0/7pAifnUs6flkrz1p5MGL2WftdRXA3NGMf
2q9TcMrEoyGpFYtpR7ujwMEiu12n2RWfekAxNpiy6vehsJKxQCbbJENzl48Oo5c7UhCKLa4SPmWu
gsGS70KfKkpREW2oz8NHQhDFeOQSoDMHerQ7LGLutheq0Z0mTlEs6liCkU1lLS8klTutk0cNKCLA
Xf+tYhsbGdhn6wmFN11zw60Qblc4WzovS//Mlb8I4FHI8XLSJFKdjQeAkC1m5/Dxb6qgFae39KmB
017cZ0Fp+7ju6wdW03OWGvTlvg2Pv1OygNk8sNOh9L4Ol+/25SL51OkBta/lKvfByv3j5XSFWQTS
rnEFQFBTmSiXkGxWRe0BCRGXtRtbLEHsrI66HmLkETd6Z4/uhGcB7ILjnVmlCaRzzezl6GCJLHC7
O/N9Jjfsz9cTCH4kVjmorQldfoP3XRgpZisXc39CoxrGD91jderLkH31sW6KO9jzRbqauMGQw3qD
EBHHuRnKaww0+98dA/r1781+lpaZJdKBMUM/CCOLhi+xsnfmMad7RdXp2oqtOTN22N7Cr3zNh9cT
1SOklB2Rx/XYHdaZcztJtOddnWoDHtApiII7nLK/RsMaR7J6GCG7OYywFv226RwC/+RgQFMqTzPG
aW/UG+gQmLQnGcRQrm/C221ykgkx7dQVUl2oP9rXX39dgwdHhVW47SHzLkV5I8xBYz424EpTtdHL
gberAz3K7z+dMri3TaKZXCVONp1c+ePke2e+P/8VazbaQWDVqQLfxfAGieMTIYfY3pubzsGbXEga
6osuVG4k3A0SfAJn7gc1bPm1OiMBfPxZnLIr+baqtT8C19O3qhGVCFBVoh8ZX07f+LS1GME0gAoh
GNnp1E7ElpdrOwd04YFz4U+nl3NB5pthzI6aD9noTLViCPsJ+GHTwZS4PbB6fzYlXDsp/bk8ib7S
eJiRNzTsVNxN0Ih+UMCiZcCKo+I7ju8JlMsCzp1ln23BB9l9N8KfknaRHNtUFnovha0J4+hPGRyz
6MelqEQ7QT+XI89EhfkUIrC+yNZ7Cm3aTEJSo9Q5G70otAJwhfSqk+XaoKEwRr+7s50HNq/0wkHN
nP95TdOlbFNzxDME4mOM6cbXOuTEO8Q7lubEx1QHn36IwBIn7Xi7x4YvookaSkqYW9ZmO4VvhGqv
EVpKl8jKTfr3WEr5prAWo4RB3u52BaRyJtrm/zD9jXCFMeBQ9ZtIcq98ITTzytxjzdxbt/bOhNss
6ftfTBUCy2LIN6c0LypRt+lA3ytpYG5qeYhfb6eCed68NLkbtN3I8ymDtssLqgiHCKYoqHG06Z6l
h+6j2htdxv23Q2GsmwmvvTz3Hh/khnuSSFG5/qVarxR431bSvIrs+SxO57bUf8/t31XmW8hQwOgh
coUDSb+cqHM0DTDf4ScMTMbdKrT/Lw4bZ+B5QoRKzdPL1zZY7fGzZ+bR8jmASR8PW0EaMII4S+PN
aR4ZcSJXV/1eSniPmrLhJ1p9WHH1ErJQLwyn4kRkqMdxVkxgyzd+qwDkHrJzJiKSklXZNtwA22lq
pbf31IcdmD8jmQIeEirv3TQ9b8UFbGzEBNunNbdeghSX5lKSYZcrGEmPisSbxD5rapXyd7g+eo80
xe2ZXAHp+nTj2BM4PrFnTQXqEsbmzGqPEoYKbxvfinlqfVZ84Fo/mdBVGbqko4vst/EqTu/hzscm
53BZP9WHFLoe2wNOjMr4NbvG5ICrENqexENBGT4nTD7QamjmGleLm7758HD0K+z76iFYJrO+EpV0
RLevkYEfLiMF2uiW/0ttEAHcsRp3i90ohA4//MVorSLP6lO8LUoNF3Xg0CcBNDiiRoip+7ngvlBa
u9F4Mz8iu0nr3i7r4NG08PREN8t/Sf6mj4VwDtQCJiiLnevU9sPG2MJPPwGp1WvC6qfhsee9KFda
uI/iSKGiRjbmHltiYfQC/0gCOA7OxyoU0PfNQ2fWkHDUKbB7TZSuaZ22NB3zplmBmDnZVkt2szTV
Z2KLiYtcyoesSIEM1Uv/dHfatMcO5idSWw/DHiVwJ5kcEDZic+1I0h8RFrSRoNwo7HJt5T44rxHX
04oJGpHNZW4UWwK93zEidYwItvDVj6H6wwNNmmLyGICBx37vLYGBUAGOguj1/l8K15nfYOvFGKNo
ojla11Z7U8PtxUe+p9aPAuz1m5retIm05DXEyJTBBQgAhleefzJ/CK09Uyi/9oo9AqtVLhRGmHHY
DeuW9itX6jHUAwqLxHaSPff6sILwz4O84dppHxqBVZKYQFb+HpSD8I/Y9Dt/LPuA8R5/mRDoLbQR
9xUaVqlI1DR1FY4n+vTkLrs5MCLVHSbqUA+dDYWK4DdVymMj3k2LqRelHGUB+ZHgEvZj1zyMuex2
C8de35OOdsVjlNyr1iH2qQMqJR/HaTTN2xNK4UnSzkK10fLGWlqh/wVcKE5QzeDkSofj7Hx1CtI8
/yYb75C90Nr1cMUjvwpyzvF02ckGN9CRvhERDAyA/bQLF9na1s4+0NvLYsw6x0vj3WjdAOhfYlcj
6H9ya8FpMtJEoe4xNoc1gL+WM8B0czc4A2oXWuZfjzBqIYAjWHTheCIgNiZLG7m9BMVwBKy2n8Rd
AhKvtG8K+tQqV1gtEW7a+JJvXYNVcRwG2gOuT9lWTwmCbkiLzVHjVuluwiv5EEi9xhbnMpDlTgv0
Xfpt46jtPuwrWx2vDruNc/ES3J1qEWch3zcWsiOOcMq6Fv1A3SbeKox8LpNaqYaYXruQxYyffA1l
2rM+tcCRb989xnaRTyq2HEuab9mO631zMA2K1umaSw80nUQxShg+ta4vDFBnFSqh+FPofF6gVHFi
lkm8gd9G3WEMoouVj/5AiN9+QX8dhT7Xs/vVYfOVX+gEB0yfpF4bvi3Op6oWGAyQLQ8cmpONHxxY
bIr3lnw2TFK/ydLw9YmlDXyAxs1LY8qQk1D6vQIq3wzEPqi15hywEpv8qDEuv85QkH4296mn1a8I
dGyiCbX+7vZ/o7r4b2vhHnmxMhD/1U62uTavd+LtMNh4WFwUddxGZM8gG1aaHzdK/7Ubu/A3CxKj
QBNJivlZ45V03AUdHE2arVGaOc9nfOhjmN4YJGsYsr3QoJaC2b0Q3uXRKrdX6ZhFHE3GgenaCtpm
rPB3FIpX1tNnMIikUTgUuK1tUQGzKSZ/dTpQUnLr7tmSsm7DEL6nrV6JZSrZgOX47KgFugEiJTyj
8cSnXdjUbqlmXDXTAvT2avXJ1IF5a5IJEHvPUbFDerh5Heer+EtQKWuUqkqxMU7Gp7EqBap5OARC
nf31KM5638WgZURBfjNvgMDJTXQQVZgiKhfDKhTk7A8l/CIBy8NTEzLC6JMcxp7Gddr66jdZShXf
+qnbVHQWHPZ8tPAps8dvGbd7IkkcWv8YCEpLwZGk7S+2amhukl+R7kUw9k4vMAFOyB9wAB5pQeXp
5pCJ3VvEcBe1Ch7xWD91d+/muVLPbGctViTCifki6GfKM0jTz0sWtOcX2TbRt2EDMjh9T3c3Ky8f
I0slsOR+yTe/hJjzJXN/o5XofFAxVU5KfNCWnAUoNhV45h6KODBqyPUjERocJXEukHjvcnh0mItT
elltUrnWk5sRo++YgTCDWBJ64Iy7uotF2UDNFNB9TduGND5z6T4r1NaBmdhkG2kQC7nKYvS16VcK
xStQymV/P4xw3TJAWifEY1BLGTMAUTiBPTjU8HLT8fk0SU6axGziLMUwzxEDalWqOeCOl/fxRPjo
jn2ahldAwawIN/W9rq8X3vnDjgvAAeOJHjNn19d5HEiBKNZlrXu7sO1EgrfBhDtAdI1KD9MN+XCY
rpdTIDPp324nZfL+5z2peHP4++EAn3WQVjqHcwZ8uUvejLCZurI31eFaKnFLtICgEAJh90ZVjw/I
NZFifD+T3NnPb2SBYj6zl6H/o7J/1Vz+Z3PXCHQmtzlkaLPIMTtVGhYFMJwfeDJazNRpaVoRPhit
2C3vUIPsUhLskrwXbWVTIbo2hQa/+dNCGvExXs8LDMdTLCb8pxl7ciU+wkSH1Aob00gU6mWVwsU4
KZ6tXXQygfSdEXQSKKYaNc99WuQXeHMC0OmBNQ2WFriWuIF0NzCF2ZGlB8SCbYd1dCxHo+W3MUoF
XuTZo3ySNvvM8SXrp7agLRPr7hv4Q6Gy7Kf3nIe7pwEry9zV924mmjIKmPsfomD+Z+tBxEuRCbnl
PXhHN5l1gQjlgjii9uuEFia0RUub0+ahT431GSnLiwa930tVaB65t406ZPcfx0SlEs4Rps8x9n3O
eX6dG8mqbOCZq3e3LsuHV6vNK3brHmHf+VLDf7ycbeGwLREiJJ0jRJajRaKcFew8+/eiBa2t39PX
pRF+AxMTjB2qAznT37GKKHd38AIvL7TFEteGGvaY4B/HzyFq4wo+1DfSg7NEFSjwEHaEqi71xs7e
mh9f/qX2KJKHAESHAY7LDXiDTAC45ucEh0MTzFaA0/KN950j5ekj4WeGxKM/EYeUgdYorcjimIql
sEg0eRZbnNj/8YPhnEFGWy7f+kbW12IuGpppontCC2IE2kHsAyMaOC1i+QlNoTKBPetzhpbxIoeE
QPKSWfKznJx9pMjeytxZ2ftdRhTHUw7c8QgLuKPvHLH41cP/dLgfikK5oKGD07cu3LOLagb4E8mb
5WMwMOdaZ5yYjwS1+7A3UlumskbzjnOutlVmXBat9fP6/xadLjaGZgI/wanWlW42f4ZqgPXFOiJo
ZeRcHVt8mEy9Xs+McsVBApgpH6D5aOHtMtI7CU9A2NEFuQbO/sY9NaFZ7j8HfB6ko+exU9Q8RPAQ
7uZOSbGAe1b3FgaJ4zZQofJiQUytTPXPxpM+FvttIQeqb7HH0CnlLiLSI1Kbca7X2qhw4NCb3QqM
xb0+8YtRn1Vboawa6KmgFMSe7+Smlh2EH/9Cjgc+HG+aGojCJjsU1PY0BXj0n0l+E17b93L3l7vb
roh317OXtrDMaEPUtHWtKDU/WtVl5ELOpCcurKp4EzNOe//MQSq2Lbx7moyhPuDUerOxN2yH/N+y
0BzApzRbvnRHgbmB0sHpkh5HKcLwJH9KlF2TexULPw+OB83uLvtEbeMOODarfQPBLiOp0Apx6vnt
Ocm65muosNHhJB9u/l/5/eR3J/BKp0rWmFWDE8FnhlPhvvoyT09BjAQ/U4UaC1i7ZnIflY+2qvlz
9P+W3sf/FzdNYidxiBaSOzigYuaV8txXYV0c5e8fprAoXNVXbyMQGIoohI/DuCcJn9Ji0/Ldbygc
fILwV8aCOyAVNZ8g5RLdV7Ssqdr9Du676SGaO/EV3aPnZbKn9wbFwbKvljMJ2rN0D6ABeCwf5nwd
k9kQvqdWq/0vDxWBQ09PdiwpTyIhcXaCkyRv0D3DUHNo4sAVfd+JZdJvjtBLopAzhAGxt0VmdxoW
oQCO5aB+WmVrhhVVxBcCGLyOJCEX8mbwKHhcy5Bg9sDN/i0giLs7K6HGbBQ+/DwjtNqMtu0EhiLO
CK/qgAtEUCT6y6cSUu5P0rsXgADMekItPAFwETV2suXdPj/7+//cwIiY8SSTwrxRZlZC+KaLRgov
CmIdydavYfxaLAdy0NbR+EYiI/aZTUEJlsp7BsDqnYsU35riNDcrIrYxuMsqSdOrURVRC/naLSFA
Ec8JrY+Q4IZullshyOCRzdDusBA8rgfpMpU2pa3R/bmiDZHXxiGLBnanQ2jgN1OJAuc4WtoyUkTK
4Mj3GP0QcTKvwobB/nbZLnWfae/+9W0aJ+fYEADb8fNKO98D50bMrnXHqwv4qnM4Z757pRHsUIbP
GLU//ohsCetqEwsLBw2dgSRK2p1YNCVunQxIiHRAcXpEIDGXpZY+z2T/PqLFTNsA/AqzEKT3+cJf
bNM97c64nMWxz+G+wd+zMee91SwIGEfcUgZBiaBIkPuy9F/WIf1RmpK2NQE4pJ3dosUJRENeZoAD
cGTp646gFl9HhRRLG3DlU6M/hGySYoL45qEZwBMb4+mnVshnpqCP7HvrnDpxhF1XjNmqDkuvJfPc
FfVv8OcjP8jDm5U/qpbmYjpVetpCiSmPvCIOu5+z1kw5U7Tkihs742PD3irMSqnsBC3eOWxafh0y
vxEDVtNFenyL8Z5k6z/aYgCKaDas8zqoSImgKnTG/f3n/e5zEv6kDTGqckH70LK0RbZOubjlOs6c
dKeiXNNLf51m93S6gs7IpwT4tvLh7S+dSGZpdKWtICGZzb312sGwTKAD1E+3RA+hiV68FRcEWwh9
DNb8HhygTIHpRH3aV0rs5dYD3c+URsHwTVsx8ODZhwVVV3dhqhJlZumn4UYUEjjidTljrTRSqECE
LlvdSgviR2nyJBe8xY0mvH3tYYG5UvPJSlTQ2Iw3dPeucbc+I75IjjQEHOHzw8Gl+ObWqnzZcZCR
Csy/oEW9/rERD6lO9CZim3iLG73M+Lc4lSKEcvySPNBhQ3J0vBX4brbtEgsEJoda3i4B2O+u3pIc
4PoG/v95VWYmGDru4TqBajRagmV1f/6nDwLPRS8+S6vFGOmWZlYHqOD0sASWcd3c4ardukAlkpNn
nNLXgRuPpA7vB7BtcpP6e2le3JyGfjatEqJwRcoKloGG0rUOOaWO1EaOQtgyumdCasgrebryVFGh
ot77bteQX9nM+hDVnZMA5L8eRmwQapLqXPIDVVq0im7yF6qE9r4q7nZiDLKnqHq/vkyZyoDt5ZoU
xE89hX05ZsnqO+3UmtFbESyGlp9MP14uaA1S4LaC/GallMmL8dddn+a4FzZ+1tDyYP5gs/S7Ea9Y
Hz88YWdJL1Td84fu2itdR9dvDA/oYrV+jhBHL2mHPJ+Ere1elicxnWCFPAL+gH1dmI2VA5EGfdN6
4CHIyu1atDM/ga1w3yhAcVq+pTdQ4xhiKD4Xm4kdI1a3/ATTPXcOeqjvx2q7Ooy6VGPD3h7NUEpc
VTzSWTTZPf5zvocVjIr1E+2eZuhb5qwxU2XJJ0NN7a3iWq6z3yfE23AqezyNtaRovf8SXElu27g4
qsQDWjn07JgHhFISZF1vFhi4L7KKW9sU9LH7Mv6C+sCwWePpHTvBS11e3E19ofoj/S+F/qgYIlre
biEWtM7WvR9ZKlSNppxc44f1T+V8N3nKPyXCo9A1wjC94mzfVDJUO22C2AFvENbHmrIcmlpOXJx0
rAUwei/gx8cXZNBvFn/fp5mW+qTX25ByC5JfxO0ZYEn9rZllxwU2fcSHFkLX5FkpINntUBhImBpd
3/rFdJAVfvHTEwUW7vPr3ZHJ6RuGbMQbsdEAdFbDw+bu2X+FUJ9O18JIMjgLsqy4EX6tGAaRCU7k
JkyOJ4VU4NHtQRMeVLtz4Fa5fTwHiei2JUXCZjfJXSw+9dFj7QTby0Ab9GhwgLyw7JPllmX0FloJ
D2cKuGRf66IpkTUPQkMB5UtCYneK7y3lwck2RsGc8PVt1Y/LJG9Nvyn7cYoIe/jhiALGqZdf5nde
sJi4JV1lShrLwpZ8NYoOmJviTqhGXUwtTh7/oAduNgX/An9MjOk9e+JjWeEq7FDvtZ0LYAZHL2ii
zSqBb8PmEWylH6OIge3dSwZffauge1Gls+QEIXLtSJIUjO1X2czURfrO9knTRZXP0XbGlzfTQ5r0
nXsyBPIKT4dG4mHTyezt0h2jfeLXRiWzZ04GgfibX+zmG8h5f3cKzNJnrMdAO6MvLkqNVfow4+PN
w4VPTNc+mttchSAFez09KtyyxA+OJ1vpXqC77vQFf9gts4GHOR2XCQcTW9mhbB5KqKbIc+jIXjlM
xy0/alqmoETcnkmStuQzcpf10OIO0SmfmMn5Pe9hhJfaOXQI6AkfzDvKqhjURTSBM7nGYARumJEO
0qTBg/UDhoH0KCA8YjDLtvei9PV6SGmOfvfX+FTgEdQIFPTAQfdWt5qzerLtriwCXWoAwXtPWUQh
o4GPw1fTAHvBNZEBEGbHwU+/EmIzsb9mhjSYcT5htRdPN2KTRfqD84gJQYXSFG9vmer+bMsN525i
GHVeUCshmzjiezXNKthaagGcTmqcqZ7SmjCSbF2roLtZL3D0vO+vp7tCHj3aDIUlpP7Rp4OnzNCH
qdDrjOe1Wecun7JURfWZB/gZoRHxEhRBKnkAzLg+ZZ5GJ7HvqxAL7aN0G/6iCo9U1SL2Eb77gjCh
tMSi6RTU+tyJ9PwHXy6Al40MlWqQoudzI1xAyBJyfOKvufuuZMXXoTLTZs7LXHQlxF/VnpMb26nF
3WNqiFikPplM8rYLA4nG8W+zOcDjYVM7xNyN7r5mMfUlYahbM0uSKSkyFyxhqTrLKybgPdbaqdVk
e6r8V+dr+cc/NTfMaXRRcmlT3q1I+ff2Dts+0kILzwcrIZIkxNqcEUzspWCx4ZZAXsfcmFoDEay8
oYnHqk33sppQYqrpcr2bXFAtfUltTgp7aNyTg8kzC1f0DPHllKJxg8G+9nXFVfasXiMqMfjQmCBm
GZhvCZEZyFBxyREiOc494k/vfY5MqGEVf0QOZLzhTJguz8OMM3kCpeYpe9GbVSLZNNZE9zdrDA6b
iI3HlwlBMTBM/yUtXHz1vNIPuBSQ0nP/WWWTuYiHlcehj2W2tcMsR6fCyiRnrxUs6il6b3bxLguo
Ugj1z0cnN5rc5u5fxb5Cr9I1hBoda3d3ipEtx+do0DI+VW4MsY53YgCRisFgz640iiAsJp4gE3G7
quJNQbdgXDbOxEz0bhwVHDvIncAJzoBVXHLMZawxeGjPUI0ZTWO+8Xn9hWCZtsPFd2/kLtDO8MaH
6yHo1/qvD6RxxQX5KyWn4zDkRwX8B8B0FtDZvwra0SLCHsUzq5wNBU7Or0DHufZ5K7vd8PssFOQI
Uw8wyZhdrA81bcdxptGGw11kxG8UD6VWQsnq9AiXssqTvJge0/aeYv92KQuXoRSQP4kcpzngQWQi
XjBNNq8Rb31zGVkC7SOPVy07X8ryAIFngg9CQ04CgZ69uKLUlxITusw5WnJx1I7nxXDRfNxiXKxy
2G5rYgTCn5LbQNAGf3VHqSa32VsoXjtkzJCfN8FsuzOBREG3wgqMOu7t0B7jJmg+Fc+b+G0RXp0H
1OcryGrd+cGnia0Bs4oFy/7vVic6eCUeCHQydg5RYRSuJwD+J9wAhD0Gd9MclV6SuIRZb3pGXLbp
81jAYL9vLTce7I1YetKvyeboMV+ip/m35xXGD7l+jY3c3JRpFWTuulZmvb3oHziENL6GTyRXDqc4
IU5xDrYZRcGY954aH8b19sS5mqUfXKBg9yLFlK6MyNXvbIpRVv3fNCqWV5WJy7LJ8/hULwFeTk/6
B/VazPxOBV36ApiEfld1BXX8C7t+oegIcVgysQCZ4cE4rrxvi5j2sjdtV/uGgmiU2YoHU4+iILfZ
B8dMt7uQSG08bbe+EfhIqT/wSlSzVeSHgdF8xk1dVJOTczbHbT7tZDu8wUw2DtBxVZ98VrkGkNF4
1Anz+2mEdIqL1azTo0G3zilrI9CFdOZM1Eo3YRA29XIapG+BImOFSbkCRXo8hD/CP3AvgAoDrnNg
WKiXpE8YKDHoupQVtUd+dA5RTOkKUfAOFwTiLPvmfYu1c5KIq3GL+HIrFwZorIobD5qzvSqpe/jn
Yw1GHuYcrIPwg/DKMj/5+jY8GR4p7TaZe971uv0JBlxhnknbUEJLTHlUN0Wl+k44sZaun+Mj1D+j
vNR1ughwyGXNDfzMwJB6QEo6yvNGuHIHu4uscE+hAzL/4SpI2KH3ZnohpE0dtLNn8C/6+bg8X5kN
S48mqa9fE3Zn+HzQw0YsGvBKBqXbILlieqLItN5zaMr9q7E7p1Xyks1fMwBtpOB/FdtDFu1iu+r8
VavoIgOCtyv/mOnpC3qfCG6tBIWP5RJcocSqXfK0l2ipf+jmpKyGeEgRq/7aUChFcDFSGaRWnyqJ
8+IAgWnIwCmmFBsalbV9+Hdd4pjzNkMfMYX3Mw+Y6heXow/9VsGl+GgAeQgF6qiCTy6QS33QqgXf
SFgTkPNaOp+lv4grF3aafgeLzaUoegy236HVZKHFGneQOwXVWEkqnLm7B6ZO6AnddfReZauCP2XJ
0imjtJeNA0azwsAaMi2rzmXL9gccp2Pa99BSEef9/ikmVxsR9Ti4zk2T9U8hs+YbclzFAekCORwF
CComYhXN3EpFLiJJWU3EMrZRWnAjrIspMicBFvRIWswHT6C2jul5XW3QbytY6SGAn9Qc9Jx0HGwJ
SSC6pAxcyckcmAxVutjbYdE+wsBa4fk/i1ULxZeeCkv4v3WozsNs0AYzNvEJ8Iq4mAL+ZwjuQNs6
sO1hIdHAXj594rXEMd4F++JkyWz4oGeo4odsNHdUuCMQyLa8lHArcovMvkk/wIZ6G8ERfOZe1Mpa
nuHrm8Leg47d/oUm/SYz/bEC/kFV6UFW857GduUu+BXS/BBwCkc8j+yEwFwhK/fsqsUSrr11qMsB
6CLk0MpJvVYkH5ly9iJR9xEPxEc9Lt5T4PZ8K0IRRyqhAr6/qv3vCW1GGR4W+ryD1fd7Hb+1e77B
Um8e+z1HL+ev4JpI94zLWr153AJ0bxcV0LmJXRb5dhJGt85vVGPtucPp3OiGqIUVpDVbFDr34SXU
1nIuPykUaQQKvRB9xARA/Qp3o9Zlbh86y7GFlylufm/xpv2IYW9Y7WVPHNUpI8Tf1tOJtngw/mn3
y8XYmsGb0/2VT8trdSlNhvmj5NmnqFI54xUdREExsdos3RiW7NWz+JxXgFHux00hx6OPopyiB7dO
QGysZ+4FbN3nti1c03Ud46/rcZIKwJYloNGtBfnK0tIlFklTeTChU6GYeUb5Yn3EH0LP9Bmu/HwR
qbKGIjFk65SYddvFeaxu51PcetR7BAyPcdCw0YRpISHzmbl/8McDFEvbrgoNpIo/V6I8w2uU7ixk
23Cv3fpTQ1a8PNK+7YOa9WG5IimdMXfI7J5BglBfXZP0as2cEPbPKc3hw8anIv/le2DyRNCrq4aV
vJZZKfDh1FwxCUj2CXEBlaS0GiO6p1cHcrxREkOYrvAUhZSWvores63CRzzmObIEyfbC/Xunnr04
nHhl3EmZS7szp2bB3HaetRz0R6Fei8nMPkaE+bYyqXePIvICDp23rS5vNuaLkai93B6H36+IEqDX
kIDiyj+hnCZwtgBXbSQhcvRbXx50ZJR2DjHpGjBQtV3G8mCMWE47vA4PA4bN60GCTRLcg++F5U0I
ABNeObz1UuYI75ViMnHZc88WluSWYuT+UlbGurRGLOlw9DFFnezNOvO22teQJlaD5b3/AQJ/6yWv
m8eR/aLcfSY5Y0+SYvrykQLvQ3BJvQasdQN4mvEfYgFRL3jB//onHBnWnCwGUsU+cxo0NSdJP+ZH
mBYTbVzeHVlYmAjNHxjNBOnzB6kNPzLBcab2SJ7A3KINIP1vNmPm/7BM6CmCtVlu2ZdqsiIS6/FO
N5we+SvjIcRLQbu4lkQbOSIF+Xt+ZlCkPEytqmQ8UKrpMaE8/dSMxTsszjxEPrUnnV9wGpunBwIr
ng6TEpef5WtNJTE2vRasCnKEoCM1CvFRr2QyloJu4wz6bsBC+WD87/PbHkH8gaftot8A+/TSYcJM
CpADYfoj6jZgC6II0p5bmKT/YcIZMrIDbyjlsGetM7smsweOdFdp6fpDxujIH6wgHSGIPTM+abFK
SwsKTgeyo3fHLd+3xR4UwXPYSv0Z+2Zh4zHiFIiCoE8OYT8n6tMRXv7NPNDdbi2MiCZgWTRh/7uN
HF2zbB0zKSzvHVQcVnQM1rQBPpa9wq9vtUfa8xGSkWryce4LCGH+wMxo5nyfFKXoc7RJKfsFWwtn
juXMxfhYT39KxV/Iw8615p3tzfoPZrbqBXTw1K3if3UynxLMcbj03CUBZ0zsoaycWCqXoDfFQc1Z
JmLOwqKVrFZxR8yx2uJjSxFhHMlzplKUYnuxkpcK2GVAAMZvqmFX4h/rm3rPMJc7KST9hFUmCgLI
hSg5I+G5mbCk59P2IE3p66rBdLh0gCxWV00VCQVUO18r35b2Exe1haRW0GTAwocvkxeyswoVwzXm
oLvHJ4WG233tSxA/4fR9Z+Mp/AApfQntqULX5XaEi48psk+oYxTcQ6tsE5IUNxixY19Or0e2jmpQ
pR4UmuO6aaCzWGFn0ZzYgCJQXLG64EaDALFhXqCwjAkrh7EuxEgmJ0MiM9vvwd7Ye+RVwoPvAamS
iOeJSvOJmvYThYDmVkYqYJ1CLOMxd6ouqlhPvU5P5bfIqs/jKnotdPHUV0mjNClOe6VaocPRULGf
BBYbAD4gpQ7B05TP7nZ7dgkjhNqxU0leDKOdyMK5xWLRb3AiewIqWxE/cKWpzS5mR1LOgcVVJvuF
D/b3owyyw74OQ4Ze097WBNsgo2dsS44Cwmx0gfmo6CLYnU98MHlxyZHdsWHZO8SRn+Yj0ZkHxGvO
Q49ORLHS96TBr8vfwF/zfVteKHC3O8viAMTngzT7OOf99OHLa4wCYAFE5aly4ZgmTG7tr2uwMB2l
SigD41WA/K1UogMq6D7sYSpLBGKvRW1KQqv4Pe2NxR+RCNhMLW8VjwLrxCVvu1/xLTMZ4fkp51Au
uFrNBFOgx0Im/fpJOHG2QqmC9YPGPmszsYo3d9FRWoZMAABx4zDK+pgvwB8dRTnwvWFH/Xj3SOBv
xxnI9VFNaJ35gFyXeLznS6tvfAxpeKwJeRujz5L0YzHZY5VcqNBrcVnvwA9uHj2F7hHFts9mYdzH
Gf7TfTneffRAkILNQTEAM+NP6QCIbAEntuqlfVVpJ/Y8gjSIkgfeMFe72og03z0Vq6TPnS1PO8Ua
z7sVC4mz+90bAzsBhB6iJMRVeLlrXAGiGUgnduoa+3WrvfqU3MSUhUadQrz97nid3HZrLlZJKBuI
zBc2i4wwds8EXckXardAtE0ZBjbr2v8lS2dqjBzzxX0zy2euGuYSsA6+PT/8q/7g1vULJZpRhxeg
pJaTRH4SWMO3lzFm3suRErwjHY6IKD3HASS/1SannQ2vcuAUC3U+FQUMh8iIBesGy19vB2pDzPYv
KJkISbkq4rODWDyWTOyzmvwmD0somi9u0FcXgCizztbFtrFs2Ew2FZdvoI3pYjBfgsK2jZkyADJa
5KyzK2TsNzXSDL1oDjNnCYl9gl1KORMNwl1JDMIcI1yuFks547/tsli6J7pkkDSOkywKyj7WQzp0
sdf2qk+u3FwcD20Pz1t1ObFQsMaIeka2Md2y8hlGrnyzG/vEhhsZyKJi8gU/8OD32zOx7KMh1XLd
EeiEpKFPpdj8JCEl6yv0jchJ2HvV2fRCyj8CnDqyPmozB8uVgVYIGjE+jitLIwWvrIltfwnGnfI1
nB2TUM9zYaaUUuBLwYGvI+1nQBbyYS0X/OofNduazMLL+vwXTcVv+J3/wIemZoUOheyHVQ/FeiTs
wUeG3jm041CJYwb2v/f657wRAfGlORgk79HIM3XReSD/asq/BLrs7HN3fcIn6rhYjXEme9hgxKOq
E21+SZeninywUWlEc1U+hg/0mTBbU7rfs17qAX5XjWP+egNsUloAest7UDztloZ3jz4TYSn3ct5b
9GKKt/RheIeT7jdHuYHje5HF+6at0aXpRKr4hr2vOPwAumFtqu3a46lPYNkiRjWaZ5tQrkJRo3gL
aU2Ki+Znli7yTjxq+R6aF04p8ujHWkP3+6e0pt9MtuSrcab/tC6PAOIs1hCrXkHqwTlhF5L4QUKH
S5TKCmbknMqsC2CCx4/zSG9KVZZ0APWHkLSzENxaHFvqmGEC01MrBdZMtEmjjAjWccoxWQmRJ+vd
4nVDsFLdqEMXQaTQsXkCkTnKF/JplZwvMyJS/wiBNqbFTFab6KNT5vyFTgRcKJOUUK7iCvPvC8Nf
6Z/mWSQV7LvaeWzKLz7hZmpUXyf2bTfiPxodsvjNoNzg7BDjiEtnCYJo0c+sxZ4MTUTqLuQ6ajek
8s2r1win1NDCfxS23UnXQ4r72Qd7QoV4tOT+nz13nKc8LOAstLXog8EjDhKmS+NFcsrjg35RQl0W
xWqH3bVo/2xRXbRV164VIOXuMEB2yIdUeykJSCTcmGk+yY1Eo4jx1iAZ9afiiH/wqQClTU7ubqiR
dGuF/tKqFMjd30bmR2Vam/xyY3a423jWzKc6ZeaA5+FZ4+8ynOVFwtiyug3uMGDTpxqQtpeciLq0
Cy6N9WU00MoJdnkh77RL/RNOS69dONTRU63n38URqBUa4CVPZqBxKEtdESvBgz9uG3yGMclpxTLJ
XAOnExQQORguqRJXJxbkSP/fmKXGUGxwIKChoNMK9xMCnpWjlYlfN59ZKVCEE+rQbDhFjPRoxbYK
KHGhqj6S50cJOPOcO53C6u0reBqCrfhnP3pYoscyZ3zxa8hDh7KT2w9I4WRWyyRMu3LWkIJa/t64
IM5nLE+QLthTvakMz9/hnKBy6T+GCSbd55RldHVwxmvUnqgYGixMHtxdCpWAvhu8mJAyIoJ4xavm
M96U3lD2SwwagJn15943z5D4TMq0eFcmMIncV7YLWUamMCdJ8So57kQZ9QziNLHbjeUEkyq4wqsN
pe0HjYkyZRfU8QsrZ8Grk7PyvfiW46ub98qjtiyV6U/6tY0qoeXrKGaOZY+lE04O6p9opF/FLYIw
woeCXpuj4kwdRNyM0cGSG57bJImZFu9EeQZgB9eBV0w74dlq/FjYYje9mUCgawNqon2gwXFyAk/4
K5pzYNYY+IZcCgTazAi5M0NYwdeN24aI2oP22UsGvVCNKwFvNZpyIBPMq904POsw2FycaERXj04e
giWZWNR/5AC/7B0DMyk7pFj0CFqslqnAF5jxdBP4j2mFRmpEFUwmrxAS9GyBlPc+8BOW7EGTrUSv
X4T9pfnesa7Jp1CMV3ckoAOFCfqCLUxXw3zZQG8TO2O1xq4UhQptprZurIhdapCF7nWtvWui59nb
87mULmPTKtIMDhVLU7rFyeEiKvznmX+FThDYCNNRxbaC6Q80mEjQyMJfQ40WQTMLnWyQGnmp1iqC
Mf7e3XXiYb4HQ6C+y9xmUBPGeQpyU/L1whg2JEMlAO6MbyKj+ZA15OC4pL8CJik6GnJIc/5WAxVB
Q4oVT4D/cgYXHJUm+RK1R0TpgqB1p9n9POEkPrj9tbMmfsFuYx6mkzMAzVAINMNZCqnD+kL+YYiz
wHlHRdkCuiEGK0vDdzJ0L5HNqn3Bd7vZ5IeXmjn2d99u+UTY2bim7DZNwe2zwJZZKonyvaxg6Pwu
RIjoMzKJrsPPuGHgxCjYTgCLMC/2qGfvfYMDOhlgasJpTDVWVF6uTyuHBNoxO/d6zE2vS626keNs
xm666LPQDZTNpyLu6S29pSl97NElSIrCP6IV03yg7lRtlAkC+OIP6IuI6z+qagNZ2M14u2C/l8Yl
1Egmc050lPf+MRitQCKDerqBKmwS2VmQYsvPHWhdssn7pvZqqnoQ0qtuiR0sG/2NkQDW+VREnc8I
sZzurnvdT5uVQ7tk5HEly6x8Xumu+7H3JHCTSO8IPYtl5zJPs3eV3Fu/6FRrl7LiQwTXf5m1lET5
BuFEWCcQ+OJvAaaIIcGsGC2LnDVZy7UK8gxo6JkfMW0oGnG+TjmIIaZw9aQauQojeeY7mtOBKJAz
siz2CKFN11A2VYhQ+MDoRvXqccv759hA1u98Sfj/RaKmj/Fj8qEjMOd0U/6Z7/YrwoftaXRV2eDR
P9MbUd18amsF7SOtExTJnJSpAi82ruOuy/aCbjtIqZQB1xg8fuuepf4k7zLnxb6h5IQChQqvtasD
i0a5OtMlycSp0946hC0C0iUdHofqirRn7rlWH7a0A3OBNB9Aly1pDJFUyr90CAPHaKCZG8ba6OrV
90h6bD/SONl8/GnZ3ZOfHzHbrapHhv4ALAJi9WzHWKWxeOYQcBbpuC51p7Jmwl3WiuKSRFSEl4oJ
uQx2LExpxOxX64BwAgdtO4jvM6m7xVu/kXgPsidDdaW9luvRfXfJ9scKLyG7gauhhy/GYAt70vtM
6PAuHLwIc21Egf1FkdYPYUlWaqEOxCyQKZSX8opnXpvhaOyYB8+otNnfezXA8u1VZR8P4QRp0146
3Ii1+E7u+vWj4TFLTW+VBxq+vaRmu6NmmQmbPdAuxh9yeyNSlO651Lk1GcMEujGGrmFzjHDkYy7G
hocuss1B4QvCa3ndH/YjJ5urSjTCilMpHem+rlLoEGl6yy8MLdS0I2iRaCM+c7pqLT/N3fLIN5zH
NDAXXjsC5JvKJHH094D4yKyyI44/kA7q+2zfiyzcTFdlBv/n2xyi2DXniaOaThCTtaTVfgDR9F9E
+27hLIcw/jfSUnU/onO6FZgTE3wnqZZCt8BCokqhVl5B55sPSMdhOmViJVzxL+t9EIWcXYflTTfj
FsKwyuxUm25SUPcuHZ0G8HN2GMdVEsAQQc2gX1c5Kj9patfqc7MZ8iKGbfbSin20lPReEXwXChnN
EO/Ew1oFJfzq2jeioVrA+2KhgpNMN62v9+F6W0KZ7+CI7mticmCsW4Pu3ftpNuHCJ2BuJQPeDZqA
ETOcAHHWRaLpEAo+F7b16goP0nA9Y/5gjWuqlb5uPG98V3xJYhQXC3wN/7MttPDXlY1OxVLD2XD2
8w/tfydJkZOQZAB94oB7TMAT+3RZc4DfrfkRLKxBZLDxK4AAdP3C+/AYDx0xDsx+U7LxFuuwv1xK
RgKbAf95pg7EI3nQKvmKfFElh9RGn/iCYRsBpC7/Zksbpb4b02zaBh0xYSbD8pu4lZ4LmgpJn8D6
n2sr2xWrDw4LxEAx7EMekB8gmovnuX5O+W0+NrxyeqFoHlIILV5C+qVZaRyC3t3rKqov0OP1Gc49
LcRauiEACX+LY62HfY8vjwUiB9BOus1FuBlkd03b77Y2ay7Bril1Ms3xOBgWpCqIY9lTzut9n9QR
aVaDos2BXCfDkb7/t6VTo/vcTMWOOx89s9UsNQjG2ax5/ld0TVBvWZSc/ABJYu1eO0gjlYWBPlv5
IFdwKp7IBAmkaVrmkyxktfkNKdPeTHRk9vmkxEdprOd1/WucSGzg3uKS8AgR0Uz0c/b7CmG7MP4u
yqtcEB0EsPlo+wAbxjl2XqaMH66Fjk3EPpiLpdtUZWxQOVxv3XrIIY85G5qDhnLmsWV8aE9ugo5x
wpGsQ7EsJxVHQvA0rwl5Ui3TLJQKE1ZzTEpVXBe8yAjU+g9HM8VbnSSk5Qr/YG6w+gKbYkhRG3qD
bFMNSZsv/PGd3yx6++okfbKRw9gNjjsxXiX1jNG/ASwwnJfe7rIxyV0fZqiFGbC4ti0/mOwNSU0K
bdbdMJVzdzZ5iBrt5I6Nik6B6iEBpdxTwL+vbTlgP3JN50eqHbumFPh6SnPpo7Yr9YFMftTpOA09
olHNfdoxGWK0vlEzmLRg5ilepkt0GJM7z9uwG770CtnWK2RuGrJJbKhCCOJXh7GP1Sq8VIpK7jT7
Vg+L42f2s6gUcjjD+da9Z5W+KNA8z7gGsyqWOZuLCtXjfF/+zLxmlDUgeWFCIlVQAkv1eQisRFnJ
yNvCaFNq6M0nEYKvBZJf/6VqJE3/BkRv8NemjVzv7Ze6FBVJokjvHGmzQDIkN81oF5HgnbnQtHNO
QsJ9o3jk3eseaqr4CMD7Bb87t9ieM28PPcqPFUqklrd5iTw0cGOgDNDsWtP7PDCao6OzZgcv7cUF
BV8CyHtKgvwPvhWxS+OAXw3uNYqD+BKB3qHJ0tre9/Iqr92Ut4+zcp/gvPLLO75y9TRukZ9kPgq3
P9ZkVjQTeE8EIg50u8NEGqIeqg65JjRWLx40qybEGvMHgB2PuTt46d/MyHKflDoqXrUzBAcnYAv9
rTbKVEmNjXUSz69/M5tBlnph58pGr8vXfxJ8g/81dwm+e+08mMqd8KzslnZfPIzsxNHJKhuFjJOS
SdLjvoPVuwtBl2QDEwLtA+VnsDw//ZJwMck2yl0ZhY26DtR06A/NgVrVerOfHWf8vylHjz1pib/W
s5P59ruHcWcd5nmCQ4LBTDevKJ0utol/YYWyl0m0U9v6qAhKaATR9BLUfhCM2VywtkuMjLILXB5q
lszz6YHzd2bH6B8sjI3cI+FaqdrllYRcbMGiSOJx9G38UYq13bXvInBvGTrz5qp0MmbT6EM8eRRy
vgtItSHid/6whJwBgQkpvc8e2Ch15H769NzTuB5aEh6QxLdODjbZZUtPsa/jf14iQsdMgEY46J1L
pbuuIcoZ/EUuI81BceOESC61yPMGi1X+LbPk4yvOvpKjau4tcXavvxqj8+T1FgiKag+gVMK2thOL
QQ49lIOu0ImqbQCFlF26F+H+OtVz5HswT0nRb/LycxmAeneR5m4Qri+2WqI9h4RdXBIjQgivDazO
tgrzu68OR6tbMV1xj70boidHqag8tymBGUE1CG7NYNaax/9eFYCCaztFqj6Uk9LJq9nSiuvi1p9b
iL6Kk4kIgav2evXc6Mxh0ITzn/oCWhGIkEJc+D6Z+dr/mqVCQzIIlTlX3aP9+Bkgjjen3GcnTjos
jjVXIDQuAfJ2UBPhJFJXZM8uW+CAcWEczUKoqDCWx9kGaTmdaMGBWYAqooPs4Cb7jWkiepYpw3VI
jKkeDL2vxmqxWJ7xjW86bwzLlRFYkoekwZKDCZnph0l0eriR0NiYTjhPZ5L1BMJBJkwSK33p1AAC
0M7wWRdCfc8KTQzN9hcxbFuaTGJr1LBJEFnt2pb72RZnz9z45jE50y0irgw54Y9qlO72dknDiHye
LDVIUtI3qxJWQDh2Q6qFi3YtkTcMxWLLUHM75gvam7hsy8Cj4gWD6qcooFUYJHU/xHpXEwGK1GmO
DeSB4F5fqHYu9B/v5/fAdx1ufKUDK0xynyaAq5q76t6/4n0vCHMJ6Deq5RwC/+AsJ0ZZiMV3FBpl
KEiooAVPiJiKisXcUn+Ij+eIqcYF8/+AoWsdOUvbGePyKtbkRm4G7deNcxJIxft59odD2rC7kPYY
DYyF+vI9xlTbK6Uu6ZIWMc6SvnN5dp8kVeX14j98Hh/Qn/XCcy+j09O2dGItFbgEwpg1jWk0dwwo
Gbj1J20hEZO3odeFiPp9I3u9z55qrm52Pm1e0P/L/lvjDvRbd28fQhi9OyDkQ+VRNcFeIIWLTg/c
zxq6gL6cBP3egDR9XvXoTNrWsNkdrv7iDvZy39W/Lrp0BuhFyjSwP9mEjqnStr7VrxiILdVISla7
NHHxrQHi7RMvsUzwocI4Op9CRIF9yFSBjxI5EwLC9Eb+XTnHwhDAUDB6eiOFOhxAkFB3nRSHcm+B
jolDtCTSbo6RqEqRNj0k0bVG5+H5M1qsMJ9j4P+7MhaX3rJH/UbzMfRJRigZtJGlytPJrUm4F6jN
kqg2ef640fuZzfKf2Mp2cLnwQcl0Mt/Zk86FMGzJSEs1cy17yelHzpr2X9Mo/3gmFeObLXdoowaj
n7OOQl6w06cmh1yhQ1jN5K0Sjzjfvw3na3xQbj2yLPrr11xK8fQNYbaKk9BpU6GOPqbjGchTCReh
c4Jh38bCngr84j2wJR1j0bHS6f2ZmphaMRf0G9DbVNQSDFQuYEvoL2Y8ODUkR1p9qURdrBc8Tk+i
EHRw7vazIUnGAitaijyeyDdIMmrOsqTCc8xTFP/W9woD4eVOAo5RGQsBFSKEC1Ar/oFowl+sfTEQ
d/72OrDNMmGLzW8t9c//gKRVlkyKSf68l9uv1lIiAiJPuaLWqFG86uVJMESW/SGp2INFKL4yAs/x
W4krpw6SD7dGa8z9DijbKM6NJaIII2wIwk6pTN1pRuBJ5oeITO3h5DmnGn9CF17VfK5eieFRXT8W
QiL+33r1t5qHmX0Qcw/N2UI1MlGDNSCKvOZRE8ZaWaQAT64zG+z3uuKmucup7hj0vnTUTpoO477Z
951NrmUzBYPF+ocOkwblkb2hG6jDvQ6Ba3clK/z/wHr+JxhWI2NQStiXoXR9zRaaHnY42pMOkQZG
XzEBJM49OHWgkstGZ6EJxkAoRr42hOKG1XMAP/74IwlkRAwWcDqoDI2K9CQkVOXYXQkOxOH+yZNQ
SNebeouJ4PKCkFumCgE90gjsu9DJNDZEoK+6cq6h4u25W7G26LFw5GTbniIzlCwxZ9xVDEh0g6Lx
jjxoPyFp96u21c7Hxngqv+BSU+40P/aApcwNpPCh+wWxXquDikuU9Qhh0bGmboVV4+EWGUfKYXmj
+QKhuqBUIMJteZPLN0jP2Bhf99uKiHNErlTbx8Tvb7tSgJYmM7LEcn70H7UDfFwJ1ESW8K6nmXSm
dWs5wz9Co4FVJTmHoYelhzOjEP9pLa5MjGu7C/yn1fJuP5D4Hn1kbcLz7F0m/6aR6MOu3iMeVfl3
yWR/hTUCaNeuzPpBhSRqa5USBLoQy31szZzJbfMVgTaoivBFgJnuiFtb6qiYMzHi3mZ1fRuUXNXZ
NW8jogXa510QxZMZGxP26j2ipyTVQsRpeQ23IrcULf3XRlXQGZaPJ0IoyodDQh1pNnmADAKrVS5z
KujRSDIU55SGJeB6m83AJybiq077tJvdLLPpDiz8ap3Siy+IkKLjbYdTA3KwmIQiZXAEphxwvQk6
3z9F2pKzLd/QS5ScpWX8fyibAjxeFkLGStHhJse0bz++N8iBqO1K1+yv+IISUKKX+7uyZ+eTi6pZ
Vus0hJE8RZRXDJzA21m/evtKJ+hjOQkpuLpkVmi/WGjB2IceY6EMYiJUyKqly8vypXtBBiiDYznd
eAtZEdDYSqspvr1Ojjuy6q8D2BGQvRsZPH/SAWTIATGGeiGdfwL5C0GDI2fLwPjljDXHWjugQr0S
P7GdC7FSs/RELMXAAYD/EorlxUEfQA7OztNivKSxaE8SqKOXyGRF45ipnOUKMNQJZtibaY3RRjT1
Pmgos6uJq2xifPxJS92fGhjctClipWYvyHAlzM+6mBqKv65c5FiObqlJBXqsXdn0Bbjz4k5tMfGG
l/5J2t+GsbWiQDuuZaEbJV6uR2k5SSJ/cNix165zaX05CUvDp96QAVwZh8+iGlMslCG0koF1ho6a
BQ/3f70pgbBoLEBPIBD7PA2zhgl/nXTUY/ncSfAP98AMSmGyz/Eup/lveF59DmnjNJAiWka4UrvO
gzO6BPzjkNKmZxf3Q1Z7kUldYgUyT2x/AlOe8SlAubzSuLhYc4abWglJatroNodofch9q/edPtqT
nTCMXbn2bL8Pd0XAluTiowggi7ItZ41+RO47LFvo46UL7X0WuBJc5nVS38ZyHs4Am6QN66e9hZxr
/RKIywBFOXmdJ0bYmSr5XD+Bf9wf7RW3X4byRAVaJvvNDXE2a3g3fdEWhFxZOqLU9jPaJFBPwoFU
o898LIoxUpXAlG2maxLVefj0QWp5uUcYTUkakNtNnJgDqk5MkPDyDEvnPNCtOAFtZfKLI8Rz28xZ
L8FfioFRBYVaFY0ELAX789wS1WluRCwIOc/GNlhISXuUyit0A4RkC74Sw2Sf7H2eh2dkYlq3GgoI
c7dG16LSjRM8hMlgLZdQJfM8L9bROTa5YiW3pkdbMvnpwU8fHM6+9u1jH25amRm8JBfg4LgoIsA1
prsomLZ7i8QwiR0XyI7mNzb0Z3Qk+oJRlcXJy2WOzss0x/ottXEKEVbdxK/6az78aYmKy4m4G5a0
P2IYkjZl9D+dUn0x+4FfZw2ShoOZeeu/bTpiy8Epor2wphBsJA3rujTxPoLvNaNK753bFUcLc6p7
BoBcV3/gilo/7FPoObmyDS0KpDjLuSPE6uW85mcRyGYs0/6INhJ1IcmB/OF6+s1fkHQcPrPJE/Eo
dpsotrB/20TM6wgkXVU9Hu81TSsk9LFLnAANKan5bf/iFhLmKDXa4JZg1vnbGCx86eKBCVD9j3kg
rkuehIEVcEbB1EsPu9ApYQBHajrqGELKlHPRsQbnaNMT3lPLJzZ6ncp98yNp6MoryZSL60Thombl
aGDuO5xHQLMyTC2okHwr4etx7jbC6lR34RmGQDyBRNHKYbpKkFK8fmrUqbAZV+RtnW/yI2DrVa2W
qpDibhuwJGjU51SM+zeZauhmweXx0a6v0NLeoKlqc3/FW3gk1Kqu3YqxCfxtohvp0q2xxDwHjJOL
BXAB2Srcpu/FSNTbFUCuwNXV5Lt3xjfLH/n8hq46utXvQKYWriDZdRV0doF4tqI46IfZQnJU3QoU
in5+LqK5NHAJI5srH/4kbW31tyC3KPEs/kPbw3ChcfF+6Ixb9gqJogQQYE4niy+rphJhYuUuKM6Q
/vlU4R+x3zeDGnzDSHeqm/5HQZd+JZxQn4FeoQfJ4IqwPninqAqGPAq2pVZKI+Rc67/dTVC/sCPL
LD3nXVDA+rB9yMGKxPRxv/klxm9XpaRiR+ggQRCe+L1L5qfhPAcGmPimzs9BuFcZa+YGQs7rWcP5
AzIvn1tZiV+7og1egv1yO3U215XTtL9D8g8DbRbn05TUps8XSYEa70n7Lyl/38UyFxVvwWhIxx/B
b2jfi93bMP0ovbN5Qgpm8TLi4ISC4maNKaQT72WxdQpcsoUxF+mryhkcWCfGnyJFmzv3h1euaZwj
2UQkZi1QPdP81WPQd3rm2L/+AViQaHuISo7/KNwRLw3La3TJPHZ/0SGlqakrLcW2up/OM6K2CGx1
ICae7hyMXJNtoNu2PV1fDdrBzb9HUnb5xZ8foPm37ryoLp9TaAYXcp+SksPw+SjYYb+dIjgl0bPn
7POqxJar3FMsuhTihjy3Kld0DzB4jSrTtoUxFmpvX+QTWJlgITewtE5spvHMdE9uC60qSP2bQLnb
EGObG9mjrP7G11FB2Q1twXwPDrsWiRgcrn4koqUC1ozQIGwu47q3kDAIc9bQE5zvcAcmyhwn6elc
3sqLTvPZD5gqBlOHnL4PN8gDtUe+mPg6XmsRK+Qr4eIL9sPAWoSQqOS7UMvV/luYIKw+/vTSlclN
dnMYw0H22dKLpMItblhxLzzh0NTDdNmBENP4LpduHbVFUycDQUL2GGMqV3sotWr3Aj9lTMcmyt0o
loBKDrr188qW3kue0VdlsCAIh2qhRRRMgU1F5vP9lWN7YYZ3LOv94yCCuDnsJrLP6D89ygzGtVQZ
DYTuKNY9QFMe2d4/LDkgPRnf06FHrJ7+O6XWg1porV0Ymok+2xQ+jPH43g5co+bLi6ZxKevs1Iub
zmvR5CQBQElHbhlPlSyIw6shNSg3UnA9dUIegbYW3Y7GmMYx+y4tMCBr/KHoceTDkbQgp9VBPQIz
NxU17uT1Wh7Z6C22Pw3fzZKlGnBQ2YFNSPbfcW7UuutzSLWBKLfGimTEJitg444r7kk7g3Pl7QnG
0Piogz/DMMm3aDqfD4UFU/WE43rzzJIkQxgJkkSyRtZId6fwzVJQHn6fOLJ9TabCyQG4w7Qw2rdD
/LCWi5wKxiTvneSFsg4tvK7JOOz+5cXi9Ar+Niub+EB8vQiN2jwfGWBgIv90T2sdu7VNDqKJjbNR
YIVsvG+3HXVtGVSAfvtEbD7gHOK4KTfM6Qc8gmVQsCXVTuKY+XSXURfS0qqg4DVE9Mt/FGtPivwp
Vw4eYY0guy5G3Mak6V4O+G5vqR4homn3qQtnugWf+mb58lBpY4Dloo63l/PFx4kF9etcaI7sRZie
VTAV54S0LrySmIgK75CfYwTuBybVTu2AJqo3QdHupvv+8LpMWCZ+X+D814LxLUGuLGgcuQGOddD7
6YMP7FSQ1/uBSlr6C9R/sAQ7FF0oRNg9xoF1Bqnms4T72IsB3JR12qbO1FA09EF7yRSE18ySPdOH
ds7vQ8ti/ZG3srALGbnQoU0NNbqsbrey31m38kbDI8mdy6OXtYZULMDDlRxTj8hDKxgS58OGXqyK
CGAepcsRksxJ7zJE0e4I7Q/8+vNeigfrHdU8qxVQuCEJsWVA53UwmeFV0/rCNnPR9Cofh8iJyVeN
b8JuH6GKlhIBfp6UP0Bv5pXj7cNGo1bXI0vAR6UvzelYcDrWJtGBuVa/l0r3aBau3GD9FeCmAFUg
WOahZ3i33S1Krxmv4xbMnkIAX6ak/q0GRdjG4dKkclIkwfuGoJ5RJKA9+8SyIh+RD1bS9sabzwID
MV9GM5DEsJz+zt6I8GiK6+iCrFLirnC1ZWp9VfCj+6qEhq1HIoJQoX1fq0byP11wFe6lvCtCa1Nk
HdG4ZN9nzOh6nuJtES/vMPAJuk5HdshrDsiaVlUO5xtSSj3VnreWlT4x07sfRvHX2CRJ+eaDjLNg
eyi/h9gJQTB67x3Xeq0Vu/yjkPYVI5hhUUFnDMWTRgxNbygXarpc0AkPvBhuXAl7ohLPa8Hihk3Y
wpj5IsgbdyuwTLK9Ro3AAb7dXPvmSknZj/ERxTaBm0YTmuKwewdb61n03JxPuUNSWGDbMlxItODP
8lzHV42q9HopdO4+W0btH7GL3G+oNmPl+8cR/B8o3b9noT7VyLxxWTjwJyx4A9Ws9VzxQ+W7Gbdl
iCeatAZqOi3ruApU5Whw3zmch2qAY5oeLyMor0rwL4U+5L+f1/uBrGnNc9ajf7kVbz35r199a4ZA
ro2Puz9nwFJ8ptaQcVWGeYU5XOkas0ODFUB76xXekt4OvO5jfMm07jOtFIVtEVKZvx7LyXOU+ZlR
o+aTM19OWCL23OOjrycSI2NrIAjG2qY8YVh1cJUNbFXbSyIZz5DQ54WP133EPlMh7/Bp2Y8QXiu5
5la9+ndeNufaBizzqDMvbSYD1RYJfn6KZeguMlbYiD1frQXnVT/e5ExJbVzqY6bFX/eNSkt+0WBS
UagIQbPMU4lHz1+FvECUm1mA9Mep5939/fooALeHuize1eVS+HGQnDlBmR7I6clk3LKZSl5EttXu
QAtUqRef6ct9NtvOrxo/QUcToaZSTCeWgLrmB4tOqiJ1dfmdPdg4sq9MDqXmRLoi1n/dchknBwi5
aePcTLEMuC4R+1+69b1KliP9sNCtso9rVMfs+SQRcAitA64F53K9u6h29ikkDdfRX9+9fq0Tux3c
jf9DQiFuHFJz5G1Dxj0YpiR1L6WPfq/MII6D/9CStFY3ddBZyDkPz/YOXvyKKwFc1//UnH4SsyIy
ULYse5nQvL3h+iN0ZetU3nJLI4UHcqAgkf33TDwFHgFQUwl1V0jpQYQMJD/3TDmal9SzTw40+bkR
fptCJemCB+aii+iWz/SjUZ8B86w9LRQuvJbDafjhA09729CPlBMmnxEDioBn9Ozu3CYHgdSZofs1
BBwGBXisxcx+oEsFoJKCkKfvipISSpC5SZA2hl81ltiA3ihr3dE2zzDmEOuGBie4rqMs/MEPNaS/
HMvQbOkr4W3bdoWJQFe5Q/EhOe+omyRjljYyz59AQAzU2iI2ibZJj3AXPx5+Ck44JXJcVVjI9gzi
u09D4kf6yyiBTgXXWISZkZYNJNNsgJ+uJnfRQpemBiPr1zDZ73sawpWREQFNs4Pgczrywf+Ukrcs
/rZvAQNxlE7INU+Q2+TFjyNd1Tm8c/PIrLOBHe1FFBZ+2y+YUDZsnCMK8QlPJb08L954QCglTNUW
OmLaJ9cg1gfno6fL1RChw7ZfMDOQrIul0mFKHzoPnxvREM1aY9KImoYE9AA9Gjpnosq+tJlfZvHL
4quGj90B2vQGiTuh3tLqJwUK0FpUmMLUIEX7CIvoj8s8X8GvvkjyYyxCKYseeoKuP9vmYXvo3L/A
7SSKz8xT4FDjKUhQAaBJbMXQ4h42DY1vWoHDeYQSUhUOoElFoQ2D4pAEEORxLGIrZUUNxOCQ+v/f
v543fXC0PQAiqDnMBjQ3fjNyGveocU2FF6Fy3v55UbrYduFTy+P1vIq9kKyPFMq1OlBuzM/6VL9n
4N0Mn/7ucy4nb4qwfyVxUrieyrXfgYAlH6UVXYK5gBz1cMBS95PS4zMrUHWTR1NVMSayfVDq9VIL
rqKc3QaKRnJ8ELMq/nwrAmntMpMgpI5btTgLYOCSQvdi+xCeRVKB8Ua3RZ7wYVprwhWJdKEbYj8M
IUXTVdEQK+p4NnAG05MjdBlIBIQBq29Lt3jVe21sUF4SFdC22F0qRRg1/Q1mHN9fXRufeHZxBOxu
dWr7r4uBGCLI6BkLP95DQRjN/X7ki4NQv9E7oletDeXOQ48AQ1JKnUW6jfjCQ6LVDZgoHSI13b/a
WhscwkEd0rrBP7Cix3gAevxnx8tY56WcAY13OZeWdU+w2Gkc2xZeHwabZCJj3JElQ0rI+7aYieWV
nmpJpV5YxWTMybOdm9zIVPbT0FXPyTw5LMdc+JPoYq5e9oLkEJACm077ZnrPPPPAW0+wFakq2O+8
37SK74WrKix91G58CYyf3PNUZCjb4g3jHY3a9MNTEiuKQLSTOvvlJhD2a0Nm045RLNB7f37pY8EQ
EuMNXJTFJHUMWU3vF/DUj+Vq02C7oB3ltidsMTgUw94/Dcj4akEycIGqZGRYGJFDhKvQwNUl+HzR
7GI4qJn2lVAGP56y/YpPHzuc3qPb+B43dq8Oep0UcNOztBSu7l3mzZuPdCJR+7oyvraLbsGdjAQO
bZIUtCg19Ta9Q4HgXZ/JAN1BG7Vpp+0pB1PpcVFHqFn8m70b3nXh0s086/TmicCboo4wiLXEOw1N
yDbycKn3g7Sa+Cub1e4N8750pGR6P3+3+9JjapnkZ2pTtDEoEiHCK6TYv93Yx0Rr9It6AD+WlEqQ
lDJydBBWH+enTziQGG5MTj8A4ZZsmaKVngEEvl0grvRSkmYz77Xw8QA/UpEC3difmpQyTj1/C+5l
8UIWI8Nxxocxlgu2WIaK7GGMPlp16HsgkN5QquO3vwT6BwjVhDEvFZI4Kwwd+a/7elJHOyqaOrv3
Wgen+n/g3maDUQabrMbeX0YjeFMMy9rd1zvjN1Ar/ZtuunrXgby2AEFBxuR1B2NXOPTOfbCSxItH
lv6N8N7VkLxVkOnaXbA9v769SJ4oqAR8C5P8KCWhuUg3LK0nc4DPpBf/bCvSl3qRld9tdG/kkVUC
UVbTukCRznq21zsFckZKxVMMI3Al2krf+Y0F7wqJzpCbp14IA+RC/AMdhFSWlRHN41qeM8s7NXPn
b77yMvb10UePEcEhTKyr5Bozyn98S6cs4Ng0deyxenxmthhmH+F9BBfS3kkVXUVBn3RXF1EOEnal
sX8U6Kt1XhYg5JNJVWmUomJEiUKrMxyj70ocnkptJVDcT4+qbujYsAkmQqZkpVFtKxuUde3aQnpw
d6pbRJhItKAbrJXscuFTxgY5WBwJYJaQ0+fzjKQ+y+LSQQ2VCKcuRQZwCA+27zijd6DsknrKxlf5
JzQHCHvkOFPrmf+zwTjfNVZ4Zk2y5Qf5udN0bRdCqL4MBjNtNOOgvJv2OIYt9w048P2FqXQbLX8y
WA4R3tLeQtWi9H/JHQB6q2vxWeJWGBYi9faVTU1e98AicG9VdCALouLW1dPvRZwZ7bNsLj3lEw70
naOmVuvwkJimDpgEivf/6d92s4Nql9Kjy283FjI5mQX3UFS8DGrBxBBIvDnX83IiKnRdfxkI10er
4a+kQ7ltwNX5uK4rxPpY5EqfVIhsWPGppVvtMzAuKapUzx/DK6Y5dXGEt5NCPmmoG+BXtIA4qWzj
eOsH14IYsswV0tck4h5pujy9US5eHNp5DafZgqW60jn0Rn7aBv2LZmBUUJPPhcQPvxh2j7EBmz2q
hy8ceuW70uUTS9NuraiGHdPRjViMva9OmrqOJtwVE5odE4ZhYHp+KsG1ahZUqC8oyU3/FNooy4Zo
vSZCOniI0HKyR3bAlWTqOmvJB6QmJMZ6xO/Ln39tgjx5lwoKFoln8EUGEKwG1hPjDpyBvUp7ZCzd
GoMkBcgAqkqoTTd5/8EfnlCpNcjMhQ48unzf+Kv3rDTG9o0tuN/hLCFvVBrPPa3ajOyhlJfF8PTR
2NZT7lFFcaAoRKgnpJU8E49Fx9fl3LMy3lOu75vCIrUSFuLKPeGLGAeVTOFs7MhF/v8IhfwvoSHA
rxwwOyTkmjC5mch9IDrZqE2yT1DYASKZ9YKVJBTtPw3ySnuMsMknKGYGDPTFtV0IzTSbvsGKjsQH
xmYPL967oEHigtQytrIxHILat1TkgoCCAiDuwZ/jU/3iI/I9I1mPaE4sUzO1jQ33pWy12B+hbIHJ
e30pFe145SznKm+rYOVGANBAuv/otUdHS7mQZ2GYoVp+KddcjPKV2b3A6O7eXmiTdG8x3w1CJxpe
ZLAdkUQQuM5OyBQp+41JSeAzMZx7IYVPfIu1u2e8kjG8JP9RmW6rvNwdTUDnJlMc4AISlFy1mErv
ygK2v7G0vRV6YutJV7DIoblcd7G5cUTd7TfyLb9Hbcs0fWu/Ba5UcUnTuQOs7dmGd74C9Z+zomz/
HMfuDSrjA5bIQUsARIa8jpIodKcFZvnE83tXqD8vd/nV+kTQrCltc5YyPeeijL65ym8eHXTiPWrN
0ZAAOA7PXxZkKuGhrrd2T2A+7fJRwdENAxaSG3tYyxfBu+B1eSgbdXKiWiUC6UtAdmTZV8VDjPtM
2L2LUIP/O/o4iIkL19FEz3oR5MBdPkcQ+JHApPTiHJaTKyjyyM8CItP6NbPQmLug90OFe2W7O/ia
mqM8zH1RwkvGye4OUCafaSJkjnEiw06PbmzmIQEPSlXVR7oSyvMdd5MJ/vWM+H+SzX7YDZI3D+CG
9I6pyWEg8jMzZ+tZQTfuVrO5/t/L0oMxza24dVo3wyxDxt8JHP1UnsSbB0E500mEoQXb8hUrZIj+
QsBL5S01fyxVRo9ILBkT5y/OYD6LrH/+yi7AUV+dc6T8Su9Nh4262jPnnrkVBYXpkQuxxdhSL8S+
7TpZ0CSRsWcUTIZbZB/nqmwewfFWtxkFp363jFtnk0aitIFQIRk+ocrpyh/YBtprLFPAYhmXn2/Y
mutpRiLSql3pDlkOXV9hcovVDHUe9yzRt+iK7+aTT0ZAsYq0KYtVqFh8dFKpVpyPZUckTpvxPvs9
VeRM1kbBKvb/0aFD8DoY7UWQ2yqEPkU2QNM+78Xtng9KobEnQ3bGNCHJG2x7+sj4vPDpk/7xieWt
Y4rCkxggmPxJgyh0aCljIu8gqYjZYkSIIlokOZ5Fmf96x3+cqHiCAO2vWidnFzSmC0/pSq2WVrXv
67ybtV8gIg9ilrB2r5i2+WKVlVlIHkITBjn/Fy9fSMXTbH4Alqd9b+SbSZAqxxz5KYBRTlYJUoSN
L0EdskgVhpZ7WH24wfsSS98xRtvT78y+JgedXqbVUtwKLpeyYN04V+JR21XPQTb+VdWSjFeiUuED
NEOrOBQKIz6bbAVsOqLCrqC1qM7++GVEMFR6W0K0ie/9gvEaVPB8FqBFKAAKzms30xDZFN94INIQ
H2zklASUtAtJXEv/tJK4dbG/oFAQLC2gFnI6GiQHGJorDv6gY9Do/JZfIsTw4EFqUl/R9v0ZmlTm
l/xv/UUrsTpomEE5yLAS/LDf/D6H26Rx46zlmP2X1exwHyDpvV+0xVxq+fMFgN/SZVEWyGyCj2vv
R8RIx/lM6h3SNuowibzJefb3TnMucqG4/iqMkSN7OA7Y/XyaUMX187Kfkyp25751kltpE57K/QHy
Si49SGYVy5dI93h1EjYGdVCHXef6hN4T+eeWdM8cMdQqe2CgTCrnxEcjMVJLWhOzU/M70HOu1dTF
97wvd47okIgfhNiuZ5LP9i4U8W7coWZ5yld2BGCAIqsKq9eQZ4pZYDKDc3mrtkprtFVCAPCjR+UB
H390j2hHTOL+zP/TfcV/idxbuQMduND5nXk1i8dvzfKueNBHysUyzfe7cDb3LaHCUAUNeer4SuGz
BInLBdhQ3/etyBJDqW9X+QArYGySq1W0tR0FICS43i6EjOV2r7vnxe43JXjs3OQWN2m+MWZe3cf/
TsoU0XYaNN2F2kEzgpZ3HBaErW9a8mbLJZ7yFYb3pb+qAvezEngOaYf2FCHI5AIb3MachZNYrjVR
+xACI1Cv8DNlfK2j4cs4GmOo4KuQdS1n0aWV3ADdwdELBa32M17mSglwhdgebnbW5Cjy0k4PlR/+
UMvq1Yw3/y+gl2D6QdMa/nQbnfMjlm6aDAebiU+lraEsK7ue06/wD6Xswbbb+4bVUPzUrnMMzmw0
faa06kEfKHik7r064WfRTfSuo4jptxLSW5ORdpsNL6wpMaTFahDroQcd7ntcsCHjiNwEI/XtwrXu
H8/RPlJ5LPHuBOtdzH/PAHSgFvcAImzxI3xV2ilSoDN1GKB08HHInaIWD/umPyrkXoP5u2ht2EOQ
2UGAbsioqnUeFwgqIl4RjmZ2STSvn59SiAN1GN7U0pZ21OcSCw6gypbj9vPR0GhIYyoUF/7BBGHm
CQOc2ALdvJJzqd2yMYl1sxLOpNlgketv88DEAGUtH52I8BufOMJ0AJVFHWDfwWUdHMJmqDDujLee
GGIkLgY0QVMCKXS5+NRFMVFvQCSUk/oJFUzvrZkRZtQfDY+pdDQ5psgLCagsWLyxXWJr+x7Gdlpg
6TSBDE3vhUbTX1CLJbWT5Q/8UQpXwHEFgxNZndxNw6Y2YkTlUUGmvJg7H3xGd9Ys+vad6YsWj6et
e2ydn02odRHjKIGthj7m33ZKAMfwK34WhQ//dOgkXWD0cmnoXRvbBjsrEJ7QenR//I6cATrhgViY
MDP+QllXpVYov/cBNlD34kzxIg8MzaqbcLYMddgubySQgjLCoyAFwSTCbfjt5eVQ99Pfks/DBddj
K0hgNKIMqFZQl74LO+LWMo3g5uKC9PTYcREK+zZDcLHX22G7DJiKfpCLF3nGdI0I/5kYcopdk9fF
yZa3BaQUJ5u5NWb9Mi3Y8BO4yQMEoOHJL+QwoyM1pxWGSA32Z0226rPdXwsp78bN77/Zs0mywUWZ
wF8oGED8pSCo8VFwLiju+PpgXJGNjhOQu3MARgEWN6g1YGbmWDa98VIQigJxsIwT5UgyAQPZzBn9
hnLpct+iWsBvdqoKfqo3RGdWdd53l1C3WpbwSNx6ownXC5whNzionwdoTXgvpIB9R6k8+H14Gcv3
kPYf3IlSPp3A2MzX8OSPoqo6jI/VO71N+YESjljRsyRZem5Cxmb/f1lUilkBl0NJ2AkFSFJPoV1u
IuSWTVvd9iqH/240LzW25MXOX0/wCSVgIfDDUsTuP93kOv7ss6b0cZZERyBXLKKRo9HFuG2+6AuI
JjPLxinu6FoapOfr5EekTNz5b2txjfEmWX3z40nj/tWqJ6htwyTP/+708zdtHAIg+UL2r0c6iEea
aN3Rual6H9x5Vr72stvYyrbVZMdxIkC9FLZ1AMGcoAS0G6imnxhcFm/0n83/Da3a0sYP2R42gDNQ
ICsuGewID41D3nV7JL9SpFvG0P+wOGy6Wb+/t1+8Eqefy4OnlTzsyVBkAGUNXGF58PBniLsktVK8
TVha3nGf8I1nc5ih9zeuCRKf8EK58LuG4AwToTinvdF8tAFFwEQWdZf/cfCLmAMG+HWN6vlRQAw+
egHXJ6A8Rfo3C+sGVaUIGtoOzyO0prVlEUWY60gijmvvbOPfeFddXjM2ogUun33PxuyxT85zKM2Q
KyztdgXAHDu/JlDpzcE7p6Fpau9fInZ+JHY3g4TVj7abjTHFNPQZutI3ziUMe2TKPQb2ibFwpg6d
Vzw6ZwJgIHdVfKMdFysCZ6Vny8fXRXLOhdnjtLw7SB6Ug2uGK3LwUUuEmiTSKVG3aDU3bMlZhBQP
RJXpPjcphUzIPhSxSka+PD7lCyOZMZAOZgKIo+qpdThyHyt8yn62g2FoIXUXQIksMTOkQQOJz1TW
q9aWWGvdgjduFkiFA3VzPBWCfDRr3KhwyNbnMeD3+sZa+tcXii6EIrxoAn1pnZbdge9ndKQ7+Rr9
oGs/dHAqiHIQeJGpPOWaNuKCtBQh/3BocwlxynTyGRzw0IGwpGuIxxq68vwec2v1AWVdRw1Jf4+s
m79SFgZSsanpmx2Wotkt3b1xglqt2WWqk5UO47w259c7OoEbOPmFRCwFr57nwRW/6hAVRixqb6Ag
eOFJE/toccpND0ClqG+Liyd/7Z4cJ7XJE+SsbXx91Hc1X3M/W89P3nVQokvoda9ve23TdaYM7uL6
p0Q2E30Gb+aVL9CK8SGwu0zi0nPQUkQ0GrRihKnSD93HXuxdHtVgUmAEzcj2mwJMXmApkcWNrnTd
H1r3Qsyj3XFuOWxx+TuVmjO+4XmMB2u14va1b+cpEhS2EpzeoUIGpUg9R2Ob9IGBVCxL3z+zsQL1
SfxzTkfwDaN+y2l4hP4ZcFY1fzGfLn9wURXEzAEisfHgG5Ce0JZKtztwGLrSEIqplDrQDhGHbGkU
Mfml8GOb2UZYQ0WkY+BFYHOZ6NKMUy1ALqfFenk/1JaZ5phrUDvIB0c3f2NyFN4X7YQ2/SAw4VA2
jndTE/UqJOIO8riG50xEZc4qhTQgSgYl4YMNzyHMd+WsEWT6pDoMh/P5p0qKj6XLGrbWBh42DO5Q
LCDttWqBaIc7o7lh+LHtp2kahzyI8z2XISIqraE4eYl2+vwO3cMPLTGe21jRd9F8tXqSaO0LSvdv
4nvS1+l/PuaJDTJOBxsgR96pKpGF+8Jq4LSzgFmSrxhxBJpSonXJrItKrv78mixCl+5pfap0N1dH
cIDj/PVBTB8e+yNkeEbNr+N2cRD7gW/9wH09GGdlZPeNyxtFTeu8js//dfKSXhpzCRSDYPYtf4Ux
MpmuQeS7DBrqC0ohVJ5ZYuefrFeWKH4jVMLO9wffgtYWe0QfRur5AlVQazug0781O4HPk5iOajrO
ZWsHpuKTaMAOFRzYDMjRBy/Xiz8ZVo8yBkg+pikoL57YSA0guvvGXlP50iCSt7Huo/3MrL954OJd
g+Z1XOWNq5EzZmA9hEgikiQgxe46JQeIJfr6DQyWEbb6qWH1i5JC2rGKp3F9eh1mHx3Qb8kjsVfM
AwmsjotX2zxx4bEIUhm02UwFvNeJh05Ox2KhLqVtykQWBp9ZObr5W5qA04rSsf1Bk7LBXv86EObd
eAojWandrSGfvNIaN1ItqpzEoDIz0bJ5IhVSF3/bo7TiS1AkdPxzQH+3yK5L7bGD00MBSdiHBFun
1P8lBxCq7si4ukiHWTNfVqfSCG0Ky05MmZ7iKobB/b6ycT1wX+x31kUOxO6bO66U/KI7Y2GFnTlE
GP+EV7BKlmzUGu2RRqlUdXf0f553PZgQXp/iVynE9tgmeB0NUz8hY1ncqTxZNpoMcerexyKReS54
mAU3tN/NVeJKq/uiIYittiHhzSQy63hNHTg+jxIFVynqotm9AO7DFJps8yEekY4gzPKDBZMf05Py
JRAEO+RNY74NKYmAN+Vy0hvmE5AGEzgRuA5MyPU/gBIqPPuNcZgry4uXABkusUGOOi+F3IfF+HG1
msSywfe1RaXaWjlfm/qRqbagczkl8junuT6ZYyT0sYh2Wf2bQw/M+MDC7D/wFT4OWEqkRCy4wJqB
UwffoC7OdYSTR1h3RN8eFPJBzLr+2j9umjR+fUcS2/+BsCA2x2iwVtZ9NoSwX4uhLcMjw1yBVoGH
Yw9yPe4e58yB1sNTCnP/66TPlg4PkEwqORnwcRZZhOOxGRpndxewtPOFE/b7flAHRF0Q6EXmxohT
eotCKmG2XUm27CbP1lOMtsFywnkvQv0+x3ttTdHB6IAdK0PoMXe2z2mFXLmyWEHBDqhRp0VMdZXR
4ySNFm6ZVuyMPWz4eH7lQqhNRPl7ajiZwzDgSDJ1VoHdEUb/F08lRBdi1EX0xVPrUhW5U0ZxW/d9
OXLbDe5QH7EDE3O0aq6svNe73oFJKkOql65CrMVo3UVwKB/gRRjSx+/EhH+6wc0cHKXKHp/J3MEU
LMNK8vvmODzuBbejJpBcyuyt7r+Z4jjnuo1cBMF1mpXGQamktPAyQov+SdfzJokm7d2RVnjuKRTe
H9B6G5KgwZMYT1SpcondtxpM3xIoTZuhdKppJ2f9MnimwstuwBrR5VsxGu177lceT7I3JApA2DzU
EA0CaMAUbkyNQAdrDNdHW1Vq8pYcqJdjA/0CbyweQ48+myzbv0xP++NORYzaq3YSsYnKvZKZPMHn
i3HFUBdgvuVFqgbVAcFTKv9tqEI8CJ0/qvRhZDNrvJeuVN/JCJowNOfUZv9h6szwhMmU/SWUZhUb
kA6EpNhhcxi4P6OWGOA4DVI0cf5yqzu3pp5O6O0cDI4gJIxJl74eQkSaZRyTybHjb/50RL2MNZWT
7G/IreWh5pwj9l9veKLM36rfth9/rspfQRmX2EXcFB/iFc8VmdjtBEdf/vqt6FCDxPrfEUC+9yLt
bmw5uy7G+gMnqRupTtKlqa0aO1fSsMqTQUDhgG0d69HaEGgabsYJzeWSaaceODJInvL+N44fmuSH
4F8K8J/Y0tDCrCancee3UpEe8G0R7+nGmBQC3eSW4CuujZvaDJPmMR5YhG1P0DGQZrPd1XNQe2vN
tIMsaoabAE+H1rhogXlKNQmyCgQIV2b0HjEIEQoFzZVu0fNdVN8hXlfEj7Nz2fAaVrv/+rCp4usu
YI69exqJDu/T74lQgM8t2r5OSoDT4VohKEn2F49IvY8at0G3LvxfFR2q0wLbLaM3s/+C0JCwPbDj
HPecXSPkVwm9WKvnN7i3/grELKduouE4BRUUCbx21hS5DeOGrtJ3mUtKqmb9k8hBy9bKrT/+xi/e
4H60n4U4AX7Fumm2q9lxxzumh4DLuQCoMO89t44STOXyf9wEhmQNdtHE+y4UZYi6SZk0WyCVlA7Y
badQBApIf3vRjmy9kqtkKiDOL1fA6yCML0y9GAqN3dP4tfVUBu1FCKSMr4C1buTt1sKo9HkxD5Hw
evGIKI6oBv32YOO+IcQPNzzdn0RodxasgZXJ88eYTTf65na9E4Whi7oV/WX4x0QA6ZVDpUjHhyn2
lXulkIB9qoGFWk7wBE4l38xHDzTxB28ttMcIe4ZktMYHZ+wMueAw5k7YKYxPXRl2VUHvGRogMKw/
9jkDXKwh1e5PAZNcRMYXXpzwKAiMhGUrvF9ipCb3wFGq7ZBvmF5yd+PjNyZvkjS7YZ3x5ROxtWPa
EOi74GFXY6RKWUPa9ZOmTldXXZvBONDOS4DZo+VRnqo6OWF9Qboq6egKs6zAIV5DpJlHR8YW21TQ
G0/M467YUxjW/qOU13/OwQ1om+MB4MfQOp5BWciukSm41FZQTOalVVvRpqpB4djC+9+vJPw1UEQQ
ilYKvpyZDk1lClqxQZUAMCRlBXUqlGXKKqyfmgnvJEMvfOb+eT2L9WTz9QmPL4NeA4ILAc4XaqYy
z8dgWHh3z2JCOD9OQxZypONa23mRs/jrTLcsmsW85h3wGEG9PYb+9XBVR76348eiP+JFwOqWpsBn
Oqp7NLWq/9aKUW7Kt0bjMynKXvYDya/+HWwzVeeE4VVFbszhavbZjMCCEaQyJ+f0dujgKad3iJa+
Dnol1QTPv/htaM3k/NJH1uJdx6KFvF7mBcck7gMmAcsBAj7CyMDwrQKJ5GQmyCjTZ73GIAlfYcNe
yd4VQ8VTSWNm/tHamtVdIRvz93p8KxPk2zcT4ILdmu+Yi8Z7JfewARzr/gWN2DB0vBDMnUHpWCi9
G6OYKRuvee5Nx0Gbwdc0rNBmFNMnXqy7KOVnTEeIACu6kq/JDSOh7JmP+0KKQMJCMOWMQNmat6lv
cbR7MBWPVhttoVCTNq8j5KXhewRr85C0fHuo4ya8lfC0UKvNayhpBRCnIJA/s8SuBk6Uu5JJPxme
kFV4TwxrN8A8vYEtOZn9dL6WhU+OyFr/OUQyb5ZZsIaX1lFt/7NHiinDvREW9Xm2cAVvYsuf0S2m
dg84Akf5RJddO5j1vOnOGaTSPWisWRR4E+IPMcfEim6zw81xQ7SCSzQfMFtDuN+kiGt4/57E0epR
2F/NmHOLbtPMhBsFizGfz8wSj4QWqLH2UQ60osbL3uC8vD1YmXL9fQY/ygR0JjejWyJX8ZTDFr4e
CtuQ1kjUDxKC2ewhB5FfBomNFSPl6KaK34aE9wdLM8efjbYdNYth7DAc/DNFOeA+DfHHcjRZBKYG
kcc2m0IdR2j+Msmg8jCVgtMNdztyO/DfceuqL+L67wCgTEkt3sVEAHxBAIjIQICXcuSBAZ+b+jWX
FcI6vDitXjcEcS6lzXV4Vppwwsi21nNkrtTtTnmloeReeFgFjPHt+BEYdcgSdFc2ZExwTnZYYkdd
hopshmycS1k/t1T04Fke92Z8UdzKeubNC2HWmt1D+tbbClEcgdyECuPVB56F8WhoHI5MHqPSFkH7
o935iNuH5kA/HxKCndaMRoq+9dqYacX/l7UKfiYOBLsPO7zmUtAvHguVBxcBa2x+AoAbQmLfF9E4
Ph/2MWJRlRlVgk2ih7z69WLo76Xs7oZu4Pl0jG+mTH5Ir0SKgM49BldOsRkc0Qt4c9T13iBGbYzL
9+x9edcOljYMkvufPUTT7F+0rJabJYzeimdVMld2m7PTIaOXf2HiJ8tF/CMjjzO3ICk4x9Bztw9d
s5mu6PvXE7Eyh+Exf+mNvt5EBeaQWMJkN4Jtgw9vG1nRIi2tQkQ5IX7vnF9ARKCzDCndyPEvx6vm
ax4FSIcBUHHv4TqcmeAZoggTZAs7iWv8fogMJbCTXxI3Fm3L6nN5Up9xUYZ3g2FitVkkFZ8qwwgG
wvOe1A2x5RSYDXchwX4PSfDxQKFT9LBCHDJFgoRZWs5wtSDvjQRSNL65Xk4nhY5eVwE09j3wxFdf
HsJj9HPvAps7sKQwUej9i4PcYFCjHriTOasyRcLDF0ezQu9j9+DeFh+pnl3ufTyezcBXlLzgdOTP
3PQJYVJshJz6rqDR4JbumDozSr6jnkckZMxmsGhoEA5SicIPV6Rn6u7f0fvh6FbDbl6kPYyILg+U
IY2V44g/8Ek2mrx2qUJuttA5rACSslHCRl3+32b67caUyks9OnYUF3DAFp+5bbjINXO3PEiBiwi8
6e6iNp2dZctY5fqkwdA3nNwcw7pRG5jfOgrtrceBakofAlL19i27/STiPTr4DS4LKRyL8v/4ydCi
Rly3Xi/YPAl5ysIElCHnmefb98RBGcBfcAwt9DErAGnifvq/c3PpVrJvdQZTA0sk81/qijdATYui
7Eo5xkfVh+kmgymILawPW5LxsMsk7J753gTbntvsufNSzeUSw///4FfV0EBBDVcqijShCQSQLb4+
SecAEB+OhdbBP0MebFdAVc7e/+/dy5hDulDKL2vJcBwOV3eeHEBl/i12EaAk4kKcQf2eOD16KCLx
jWYwXMhDrl1y6TOzAwdv2IO9WPrFoHfGGMlfvwVnyqbLpw+eMl14In4eWQ5EAwqxKyq4ukLIMq0L
+s+56QmnWfUZGCfnxMwEUT9snlB2ErZeMs6RZhjyh2+mA1ziS/YPpSp3g8eLy0UKE5hJjdi8xvIs
3LLBUROaO5GhILZTtVhSaYh7Z7jQn1kM0xp97eSRb+uWZNQAiPIZFWl9q5Os020vYtt4vJX+5t7a
Re44Vi4CB3neV2HoJ9890pGI1U+fgc/a7b+ws9gA3xvhw0/bCTDqWxNqOqgnaG4iGJ+318i4Xnjm
WaPii2vXgogwXplR2GBf8Y44Mw2hMBIHie+l+G2lDxiUSyNWVOrVKVqBViUHxRKmQFe1LHOW1iCo
S+jlGOjFqYU+7qUbHBuLU02js40okUfW883ZFq5kFOq6B4BO/nfLg+0Q8SRmUUyAFuOG2VGJtSMO
gPrR2Wv9KT57QgeSQhsIQktxWu1AphGvaopXz8vZla04vLA+UnBnot39NcAEhkghgiJ9BczWLlR+
t1KhNjCwP6kUv3Q1FJqSaBzZmc1zPkiISSu6L8HerpeITdUxoksbxm3p6OlYVTnuVJxaZYxDNteV
B8vTjcIbSNjzW6UG4o4i4vIQzcIBS6xaU2dAoSLzk5AI4F+VDOAztOBU37ohSBf417LxktWCviQb
SnQpCDS7N86lj+mIEue7ciEEDB6hFyFNgPxpbEsPY4xhz0/+mnk3ki7LSzsMP/P+0GyVN6dyfQWO
rIcPOfoZwBZna+QheK8QbIobfVZS7Iyw68rSACruAPF2LUuNFu0CKjzpLvmfRat6lV7ZswQtteVy
NV3Qtp6Bl6rW8NArd+hYZPzufgPFBhfsGhHsHXacKpUgR/FlCW97Q1IznwXjoENipau8jhGS+yy/
F9ObnewFTSdR2XyeztY1r81VPzveSnzdvcoZEtl/uxVOLDxitDdWkfMqwyIxnib95gKTNySaPLT1
eu7f6ThX8NldNtVmzG95bXb5dKuKKhfoMdrGUzVXhlVuR6+tcAzbh1q/rTSBLydzfMXgdEcIQWvB
OsWO6c9vV1CTsCXAP2uTLII0xcYlJrDhitHqGrUVBUa9uodD+eLqoOhoFEEx+rwtdcdALkjI4+9B
iu6TCwEqwb37mS2BkwtwH3Nbu7yFAGKFPXg2UC67jNIsGCZ2uLykuOvA54PoLdCCfbtQAMR/uMnY
jZzO79O8k74z0w1bVCZwt6eJTe3r+t20HsuAsRpQxQ8+vT7Md7i7TioVuSrjq/N/tLgcTRzcceW1
Hr9FRIhq440F20dCD6RjZ1H9U/8oG9QGGmLQqApYws7EM56vv3XWd8RkbZf4fUKKi1pdKV3lLDf1
APqL9c11/1Og6KQo1/eZbWeDzEwDNPiWa7HCKK9sTvoUuIoRZRYvSuum+Eu/lduywzMU8Fr3LrzX
F/G2svX/th1mRcfN2YHEfMAVf3kLiMnACIpR3QgWKdbcG4WS5IrD6WTlr7YgmEknEdq+CcXoAEBr
w7jV6zYsDhKxz7ILQ8qyc8KmAmhSyC61yb4Lw1itCKNczpXmBr/K3w4FkoSSFRVFSuVknigTipcs
xyhme2UB4ea2WE3Aqp7HEeP9g3pEC9JFiFGXIEXR/8SczNG07GZjK2O3LNhMqTK/AX92mfRZsDQi
YK13hwyBWf8yGywCt8y9DpNx4Poq7eFJTo58tpP+8t+T0ll5U0g3uDk3MltR3b0SOnv05vOC3t7I
lAjonXZW3ZOcfWj6NVyV3wkU84AQBNSYVsnBHMxuhRCp1g1YpQyUpSPjHUhCSudlAcNAP+QR2it3
hEpssgvcEilV5xmk4cC6+SUmsOLCd/VFneQhBX3gD8VBTlCWKcsXMDn2xlJA2898oBG2sjScHKlQ
21Ez5Bl9Ay0zcXNultZoyWADm93KrPukpy7tblQGXseLV51xo2ZGr9NdwIUKEg6e/98LNKGYh37x
3j8janbf2KayADO8kXGjTrUGqZjxvNBBZ51dQVdXZqeXMHv2a4/tI4tuXDE+iS7+4q5go/6S09BP
nyjlCWHOxfLXMGGu3tqDIfaKTlKGoy5ZB0lMxnwwm7s6p56EwSeh0yIyKrAncIj6pcMPrHaiB/iN
UPoBw6FcXaAK0nhsBEDrZIVG7B/F1zA0dS7IvBgYnYKQDGyaL+QB9LjuEvrV70+L9k0NV2TnnPlk
ASWiRSQK+AbMWPRRDwHzvBGtezEJBB5n8ZnRXSG7RCFxyFKYLMAULGhBQpRuzjtGmYkIEwHBj7Qi
x9T0N4MytXafEon9/pjnPbln5LLOnkr06vfStMfWq9z3prifc03Kk5y6o21EqukEKHkJbtFSh1AA
5qVOp1wg0TA4YpnE2sqNOq4PrnaWnfcmQk7bGA1G+rFDLPPZiTzLX6CJkw474+sZmrTsAndCNwro
srdp2sjSJ+ej4TmiapSCLxPDsyaXjTnzEE3T/IQdvXEKRFYn8S4lp1wNo2UYBN5ZQwmotJBl8Rzl
WkULsdpC0DJ4gBM5uvQ2qOpsPrGgrXveRi75aZVyUZXGnv0GS4R+gMt5m58abtUhtte/vAPwNPwt
T+hqyp30kZInfU9U9KpV7yQpUGGCCm14yTZqEl8SgjdziZ2lOZV0ZFY3Q3N+q6i6DbJiJRKQhG8D
f762eFprmq1vQT6A+/0Tyy377AvKYtxxf3pUXpZTYa5WGzTgbbrizraEiLKqV/3E25HyrFUoWHb8
ZiztPVBUhR1plFjB5dS4qiu5gtVCmYAkZuum1LGMOL+smPvVePfVUE0za5NGcUH09DNO9Bp3vkFT
A1F88MphqS9pLEy1vdlCL+GlZPTu0XzYnwPiomDRqjEdUowOco30fr1k//hzA11a46rZ2zgOQqOM
LQnFq1To+0kQ3wPMoy1Q8BOf1qUf7PNnfqdzs08v3+gY8G8K7bqrE2zZ2ULqasfzWkjF+bNQEDcO
ymygVuhQHKbsTxiI+D/kUIXooUmpbfx9UDZq0gOBnIibUWeMblSFjxPiq9T4+s8FipUzkdhDey3F
1uDKneETnYEV+QTRZVdgjR6E7UoAG7wxFHl18YZv1oFFf78+RTQDvTk7lVaSxjEK9YE5WrsiBK2i
Azi1kQ6equlTMHohkNJBnnewZ1A/sRwpCIuuBQ7IIL2XKvjhT9CJtFgaW/ztH0mG/BXRRgcwNK1v
Zc6OMMey6O5bF5GcCmouehvod1gO8jiQktx8rQeZAA4VuZb99Bc5AJqB2e1dn9AfFY13l1hmmx3s
b0/b6WxTbpaJfdvY7TzrRVl1v0iZNz9mazSSLEeuwyiOXm0QG2bpIazKKXPiOSFKGYUi2ximyHcp
wyxtGxAinGhtQjcFwEVev10cW+YgasmrGjfcPBJqjCU0ZZRvyRvvH4bir3Byv529nD0647T76vfh
1fhJQlH2GtgHzWY2PXb3AV9onSRWyMs7VjVJkXjUdxGxWCHvTJqAqKxxxCoDeLDd5/blnxvmoOte
mpfBEbGb90vAEy58tIJ1Z1JhU4QdQm5a9PeHtFcBJwjg4xi+F87AX34AMD3Vv7cQNHNcAAsvpGTb
WqbzWDU7GmiUYEu+2+0sU0c9bNe7tPUcCTsPmKsC2QoI46EU7Qo6qEJLpjkw2++5ZLvwPn+frRIe
y6VJjw4omZ5OFaBVRIcmzOvCcmJk/sa0qzxfSTvh3xvuuJfDfBiz6pLmm7AKqtBOJMXz7/rLq5MB
UhO07qX52TDPuCR9dfJg5qyOWn8Ygd3nHnwiP1Ar/o7qwECLv5hcPWWwHMR1ONZ5qJHLaNfcMyzJ
XvnLOfRupbJ3gx0zde8UzAWEw0rCX4mdZwyP8zbLjIkWH/VQjIORul/KYA87zOV39OVMl2Fily/u
ugAa0KuzRxpvjylB2odf2motq6xbxWx1A6R/cfnedILlauTxCxeZdvzLTtTYstooUkpcr324D7WT
1tBuqRyMuLbpdfc+wAv5iA+8VFOuEea5Ldek27F853H/zDcHKb8RKCNkPl194h62d1Ifr5aOqTh+
5RVyw4hXGzodmBQ+jUqYJT0Q7w5UB9POwljYgSjAqI2vC3Y60eHCbSuTlkWBp8jX6pFNGFcLd2eH
IEEe/o6H3eMp55gJH4niz4RtqKxp26FvN9/ZKtob//F7UYHT8Zt/hiskZjgPq92z8himCRFIdsfu
/uvKk2flwlWFOCuqNGob+H+2lUoAcRv6RYbjF/R38gNbS6e7Io8DP45Azlo7hD3DgxKwVSA09jrl
0JuuA/ZdbwZ/KYbJlidtYt8v1e7w0lazc7eH2mLT0FHeZIaQZDhgZUYDP0nq1vk+kKgEnKeq1Eu5
pMF0Tjz7O22Jp7PBd2Z+9HzzwpGyvrrtLdZGpAph74JHE/vL9Jt2AXf4YMYgb1uDYPe/S1UEZIvo
I1PLkvxX6q7BBchmL8C60havKTjAnOtXqyPmiE/iCXfHNj/c8DGRUEjlEH3ofj1mvuo91UWo9EAO
IzTDEFpuXa5/OipdpYUPPHBiekzpWTDjaPNbg0unOw4Gf+g0Ac5DJ/pi/qMhDOPT4yA8zeY2APve
Km9ITilpimYTZO7xQzDzElLP13pYgjWBJRjNFrLLITwlbcMfsc0+5mlpHj9Akahjx0sU1tWb12IB
FZm2XrnH+USdQXfypfvtTP3zOPtVNrjaSytudfUwJD7LFDvf8UP2AAgpxtEJVdxmOa3L4KA2imN7
K7V7xzydbSNeWwz3QSP1H3O2jML32iFGV4lfVURt4YEIXf2/he8fIUobni93HxUSXEjL7wWcREXU
rni21ttLsU8rHp6VI/NX4Miku2cUIgF0OOVhQZFeNdET0WWSje65dZprLU8ZdyFbn2MG/jsY3EAZ
vojtWNVqV5AKZcknp8dFkvlKFrmrACiJ/6Jy+zk0oVfeWqZrTfRqrEUSLA0tGTDBWQdagWuM/6S+
cPyH4rrNuF/YaYOvwsBFQwPPI8PAn192Lf9O6rS6WeUy3B4BhZ610pj7hT5etUgGIlEd3EKkkXma
sKXgCLKrtE9C7aQ3GK1s+1OortNNTRdKZSfyww3CysJxecZheqODPSvZb+ggCt+uP9yo8g92oc5W
kAb4DC5GwajaLiAm2ZuXuzqtzkuFzD9PFC2NiVcbvLlgvHm/l1XqABBN8LspjkEVIM5zLigxntmf
rVF6Y1wD7AMXnUX9mIpbrm77nNAT4Hyv37wTP+NsG69q5L8uXLoO1PICG7FdHARAY4lC0COFHX0c
n5o9Lq3avNKreNbr8JIN3VanR8arROo0K7WovimTn1Js7bAIbn+nmdMSyjXCkD71Szq4PBYT6iWx
soqY9AOxH7A4TQ+rECMaOEGCCZIk18Yscg8iOpaGQx15zcsr+WXYFRCDBLHMczoJgYDO2cLUSnwn
mbUiHTfywt6sMLWkfF4Z62m+3XIlqrtELvsA/aGr0BQRNTMq4eYOFwCMGmnGqIC7k4EWWoQyFaLs
iH5aqdUwOM1qh7z5pKSQKkAUkKBxQgjIzzCVIJjvXT9+WGpYhnUZmpwqCQbYR0FqGxlBZF/EPM86
PWTxv8LN/jSjYVx7f/Q2uy1UVBCEvbK6tWMy/X6C4aaJDWWSFtJRz7eFKTYNrrT0MHnOrslNZITE
lgQxphjgyrHUCbe4NOmQ/osBKXZjiYRcP4KdimmG6dGFXxgfixJ1m10a5YXDQD66r/jkbLgVGx11
SLJ3NTqXbKT0/rnIpHCvrft9Wffv/FSiSGznIPD82HO/RFmwPqhLbHLb9+jtrFZCUZIBT4LRlBsL
0AFwZI0fkiBYwZUUV7bi7azR7n/UFMGXS31OnroSjzgDILjPnnUKHnkF/ALv+t2FHoe/HGRWXG36
DFhrffBiAH3ER1tm6azOfqEIElqiGtGMlc9nFT41Zpyr4giYbqLn12y4pltGbHyH3Hb6i2bhVfCb
g8/fS4CF7e3U1/XxBBx4AcxUE2PDN7wBAiczPPaRfuR4gEvrtQzRiZlBe3C9bpgozYucg/EwpxMP
IvBQKNYtnU6fgXnjeuF4Gqu/olE67INOJ/KEBG+JRRyO2M7ueW9C5ahwbqgHbrCOycbLu/r0CM6i
aNTorciZYQ1P72/5T9SmwOdVFV59X7xvPPOvWZApYU2YTJshY0aluT3Dq/AZANYfprn5cxHccA0o
igGEWKEaaxKsvD4vNIucDNcITgpHsKnYOPzxJ12MDwAAYa3xgAKlQ/EJ34O44EGfqgW/f2FLVBdi
VSnz38M8PMTXkBQrambvzKMgX2XVffic+ylFNfLTk62L1DXWMQqVarTkSH2bvSFKDc9AxOCtB0Rp
IOEC7LiWJLqlvt92zwO3IA5VJfR1Mzth8RAz+fJSa0dlQLimHeQDupTRUzgN7CU0kYbNEIlHMbrA
NwJDRbbj7SVFduLkvz/QCrb9xJwP8VcL5/68JLxbpKeS32zHoe0lPX/kqd3ssh5Eu3nEUKoL7G32
BBgpck0rkQrhIdgHh435Rkg/ai8RTu0BnZwr3mv770gszJdozj7KE8lwZWobdYHcQBknJTwhJUdA
ko/jYkD+hjmykEnYmDe2s2unaeDLyCYTBIBBepa1TZREVazXKxRPmFmWueRyqR59sD7Qz6ZcGx/g
ak5t5Qphumai+QMfEMnucDonR9CB0rAfL057E/HEItniHqz8ieAHEptjVqb+5zWhu/9yqu/disqU
N9GKP04t2iEUb4eOnAn5BOXIBBf7vrJmIwc/dkepIMA6ijihAZhuwYb/ovNE6GWt7xYPLZCyf89t
dE8ehfKgEAGygb4Xal+9CXhPiGqceAf04A4Mti70IaQk764oM7UkQHq0ZOTqthJmIWF6YykJsIgo
Q8GMx+0Icf0oYREMqyssVR41vp5cq3ks0GMOG4sfGLNRbK9zuAhZ/rziN4Mv+bhpimRLbOS8j+V+
Vi+RBKgJd/0O1ssiDIiELbKJb/7p4QnpC2O3a/xuCsFafJT+ZcPbf1/fl8LDCNPQtbBeoBSU8HrU
zbVL9nScoB3p/Uzaqyza7a+vKpdf4SCX6jdJc80EYFJ+orOmSsh+R65zbtydIkqcWgbO4MX5/i3o
bgqOi/R+mo2rUoXnSg3lb7XEfaMu60eokb6imQOq/BYpodXE5Pd0RZQLP4SyFU82j1xwz2roVyn1
1pEH8ZYXk0cU67Jbzv7aW6ZHMc2WfYMAE6UWtIPCClh/VoNy7FGwlrAj0UgyLomUv6cJD8BsKefy
Lyv782/p3ufv5q+909+inpCExC0IvWrNf6OitmnNyH77aT6mtVYHIxbr9grA+vUVAy8PrZKPXvsV
ZipjoKRQBIOOC5sJWTBts7LTEpJUfunR0YzsfKvg1uR1gxo520KIvVsAwcLa5Myg68FY+3K05B1x
3uLL4EwXFv3POqn98+tx1K0zlm8h7uTYRlCB9OHzSCr0+rAss861oh7n4kfSmRJ1+jq5w63wICK5
TyxJv13vuzCj76HNZS0YC78QJzugRu6fJoF8v0RG4Qnniose3h9cT42iwEV36n40CX5gaMQgIsBW
ewqQYpRjxQn2xAJciVED6DkqEurgZSmCP3yfjRgEE4w/s2VxST/Woo4qQ70kkOFcpv1PqZ5qaIx1
RoChfA9/KXtChrQPb3DmxxW37rVqhMagFQsJaEChVABi9OnCZTKVp7K3FLteK4yogUG82xfuS1vL
6hVfrHo/rwml01iqa13pl7A/9nNYJ6Wt4OITnrkhB3mqSi1IRDfJggvgO3pXdJuqgIuETgBGDRNM
yVG45baaEDS/HKNQ0R6A3/bW8lNq3yJcVokghQyTrlAYQZTZOMr6O8exgEeyh+qo7BPMEkt8DDyS
e9wR+eHmA/K9t5m/LwZj8Qkp4qnAgXwsud+7aFsG3hdlT+CkV7S3DOZuPZ7/SfVoANXZDsmH/O++
hnzxNkHK9gjtpUBAaq4PXCHEh6AZpCQZCH6f9bmu0j2PvMZpoSzgfI066NBM3wj3U+e2Ub0nwkhK
d+IUTHb0Yrb9nfcheIrS6e5/G6NjSTHqvDuo89mE9GEX09ShRuruHNJZvlSV8fkL6viWzyeIWx8u
qPhTESbhmnt2AwVqU04ObTbcnYKDiKTcPHGUMtVpagrBY2evJcKBgH3zBBUJsExNFGKce6yOc2b2
XSU2dWZnvrk62DsQkvwKqQdhXRS+EdNyIcR3NzdDWTL6Fi7K2H8acC2qY//TcZpKpsT5Xvh3S/X7
xZj/sjA+IuRvOp/oioFhyZ1UYLPloKmSvsZhqyTSHOl7LpGbGu7UJHQw7pQ/00vRoZ4OmSSSCaJJ
u3HtaUagU0gBjuCo/dHDWFjvOq18YF+YOpkJFmyNc0iRGfqNMy6aPbciLDiFWSbfzLsLDYB3ax65
CXQMA/N+kCyUhcbqss+oGRokiyTwP4Df6w9iXPLwQFE4VJhB+Y3nnyCUHF2NiQlT2qAOJ23hXz/1
BmanyL2wF//ISeUEczeyDa2LOdSER/guPyTpMtckeaSLrTiU4zYBjwBQ3i+b+Eztd7tlctcl3y7o
G4xS9mAHwUkas7hQpXB9vHvjIB7q2yWFITFYHIaL9mv0GNk/+KqlY3u8tqjum7P6qkOG3k3J/zgj
BMrlx0gxnExn5ABCRKT7cKvNgyXwDC1/WdqalkVUO+EsRDoZPuFwgc1A8Vj2h7Sr1YPuCOopGK0m
blBNuzWsZdUp9tXrUfdyT48nGHlE696Ev8Ng8HsNQbz9msCn/c1agMvyHr35WaAbS228NbEqShi+
hInAA4PDu++I8Sns/ndb/r/j6IRN+LRq0jecl05HDIaiOssPyDBTtVb49zNyfbvw/PFPWklGkh1v
grYHnYfszy7UzjEaOU+nRHMbdUt6uRPlfy6QpSmT6UY7dIbjBOhFaNpT7ZjaoZVK5boWVcdhyRQi
2QvL/JXA0tFRvkhgHUYlUDc6SgIT8f6YuRJ2WEChdeo7oE42PAltZbs/8fpKzSfJwnq7Rllsrs+f
6Jqi86uEU41n7WBb87dSBY6+LhHntZdjzbPwvgVtsb7ImFp6mikYSLSaim51tTWbi63i2tCeZEuz
J5z4kIXjlMVznRShXAgUDzXidCeJWm8jj4TV4tVpvRbJCOW8u/q5AkHeEzrWoZZ36V9BdDNWTtpL
sTRMUql7XSSMPlaL0Spvpjy6GzLtL1pRjq9VRa3E/qWM5VIwGJWPyYBoxqRLiMLY84ybiCETj0gb
qxLjqz9ZZTUGX4EMLiYmaNn+nIHYjdCDbYVfCgI2EStpeJOryU3++c3bV0T4lpZR1WPqu/3kQzar
bcEdxb10YI1flwLX3NNv6cw2TDL8wPDI4/ULRA46SHTCW46p1QUViJEfIuJa2aZIdj7ZHPOEYbqR
Ms3SPwR1mFY2cHrYcqIAO26IA62flQRscmiRmAEeUZ8VIU3dVSS/IgGkqQk9olUjv0DR97kTnIpi
sEJKm0wUuKDtyeOzFdhaecUZYszou3n6WTPcMaDm7mnHLHbdLW5iLW+ZW+Up7TokAgowgBIuZWiR
OQg/MTC2zqCRitlH4AIWqJct6o5rIxP3fYw46/wWB9IFpTSsqzWCa/t778JHilFZfBzdIrYsMHIK
UmsVXgpu2+ihmUCosGFTmt6JYZTiaPsfGXD4uSQvbZPcnWbl81MUkFq+ze4wIr+vhmo3vWW9w/9d
S0pZjIDQHkMDWJvO3uqJwBXvIrN+9VsaeP8dRnjwD9YTHLLTaVs0FB1kiveHPOhqemvBmjqG9rYd
myIagosw694BdYF5pLrrxd+yfTm4dFKdEbFepC8p0mlBDs6kDeuVOmg6lgqsNLUAW91mclyh2ulN
KOSb3vKMV6fVL7u/hTnMOwKDiz4Zm4KAaoCfEphDsw9mVYEbNhuOqqCDx6O5v4Z8apefz5tWpA3Q
bexSt5XXNY7iqwtMx3yAvITCpghbjZp9hRggtp3ncTDNRXDrOM3opDi8ZInwpR5hI6I0TyIy5gBu
R/41nQhpEkDULzhkaJZcS+gLkGYe4DZ1Wc5pNJDaIPhwGKKkspFQ81ioEnhvN9kyDKLxLpaenMTY
lbRivKox69B+hb2+OQB2SqHr9euFofu1S1Pbr4YHFBA44Y/4UkX88t1PszdbbCa982xoz0AifjCM
nJ46LEAj4EUL8k7m12TXW02VdCK7N6f+USnXVWYOlDtlQAaR3mLDVceRV5vtK0bb9dHbsjD5Xlbg
wEtgHsTvcQVeRi43TDfHdC3R1+0TUQ5yPRoo3n+lITbbJ4erb/zZ5VCMOE9+D3vguaCRMtlg0nl/
Yq90dpBNUVSWozEXY5BLPV0wFf9zBB4xw5EoueaATOS/KwRkv8ytDADUOvN12Bkw1Dztjne8qZxE
wLjWKF+YFdx5Ozae0TpLkVWnIJ3fj5JPSE4Y2RGF+HhMXn+kWMuRs+WVHEzlwc70kLWYna0+dJF/
YtS8yM8JNGGiOu1GnEDj2D4gco8o0nMOTTaSnbjTfwrelNH0SRljv1p9avlweIvlzWNpH6C47+EA
1LqVd6krNvO7MoQtdjgQGRJwIEf1wyk85zu032f4KTaYtoGks9fG3CGdysn8MbEM7K/yIjqGWtsM
r18w/FWU9LymTDyu2cBm3dqpUs9l3hoDLpdci9nA2XXN8EaxMFOsQZp6E17LlA/TrtnxBs8jaiML
Ra3Tz2gN8X3HORa+g9fCUzcCVmZNLsFAaYwRes0FJRz2wEYA2TrPDNRsuWkqs7kxbqLr1N75U5or
sBL4rM3B7u7D65GfArxIivp2MHG1/gvtHl1AlAMoQQSR0im0Jix1KgEfgS1FIuPffgv2MB2CutH8
2QHZ+78bkPrsfD67HsD6MuQX1++uWrynO87EnBqcJhf8dSaDhw9RYSG47yxX2e2pSCgVA4mMrbEe
lMvNFA9e6wMVMXbztAhqzJOMbbQH2lrFYuqUurt1k/u1a0tB5b4UxLGqrAIoCB465ncp1rRsbXRe
6ZNx6f4BY4phTPWSuJvDcGeEmgOoIYIWlKzspbOa4YffSwS86pKMpo71sQHE/HblCmcV3iEQiJjj
IvegohvGOyNJitgbrfMCue1ve+VIO1qWoe1Qa9Nyt3NY4GX1fD18eWhMs32bs8lFNT3KUKJz6uEQ
S1ibZy5kM+HCPOC8j1MORzOUliDOqHmkMVO0qORvSchIMeH0vnBbgd4B3SjpSGsXE38ofY2iIie6
QmD2j3F5eqs2942JtKk/9ng97TBC20p0VQBqCM8T6PiZCGJV3U9c/C6+lLRGqwFkCSCJ+04mhLOw
QPjl8zYAHafo0l1l9Y0B+2b7v46td+sdQog/DcMJ7jJeAHIMu8NgHhDotGkk+3ybh47AcVYBWhV5
tNz1vKZ4PZ1Xfmy1KleHsC5+w0eBwt+zkccXf46ox+mR2+s034ozkaG2Ah2y+OBLW1kvE4NJ8V2U
RLIE9fU/nau1jHsodkE0yqzDaxSEm4/1DV9aDWWLP3FejWij8w0GcnE5aFbUcRR/KfhgOzJu3yji
3OrX3O0OvBVYH5VWz98X2H8AzvYYsmqDJzsIA2AxYSHaiAYm+G6ajNyeHaNxpUEs+1yMlDuefMdz
81yG2ZdnZivr7KE/LHJsi9n7lvuHkx2zJQ9MDJCwbh5vwjvCGNDQoJ7jTC+ruEb958L2l+ONhFk6
UV0pE1poioaaq2Ly5QTqUVE19fj9OYF6Lu+ZeVbj80JbSm6phkphGEX41hs3O8zGwl3eE4l5AhYf
c5d4dPZlIarU8meXomSUA7vhefqg8PoZAIHruZsvE6Mfw0w2ZH73jH6zbgRsoijEZjgDPXRRy1+f
DVVPePRUKFYnUMKi99LFXBf3SXNBGlE2TnqBRh60kI5QHd+R5NO/OS8/SqNwb+AlQM4bFiAwWxPc
At6wyN4s4vzzX1E/rXCHE7FL1nXfFrZVJozas8PX1TRfBhvc5/2Ip+XoAGIQA1eUPb390ao/hrsJ
HHunIO5MrE9SHYSL1asg8jSOoB9z3k7FXn8RC4Nb1OmlQtMDGTpnAGIF1+WCQDC40eGed3RLn+8i
1QLcL1H7U8FuOkXVhlZ/xOTk7EeELF919MiBvfLI9skS421ArRRdrM/JxmovyE1qAy9+GHjRAcod
G+Fh7n4y27yCn0c4WnRozoVUdOkaX666KgcR+S8OjI0RDrbJKXrU6uSOqyIHZT1JE9J5H/6rzdua
vmm5e9NIsPh7NEREC1MAOUedQul1lmhl59aAWVAa3RjhRwpoKQlqvCmGZc0Bx4bv+5fDF7//mUWf
pC9TZFPxWhk6QnJPEoqcB8R/X8be6EYfgugcsTf33xGC16a02t3fi9fCmL9fAluWgDCxtyxEfkx4
4BCRtRrQLUXhkG7G5rYwA0bOpisnRUo9LsULUAXcRot2S2/ypkcK6IypEANPCGPcGEtMTM9qBus3
tM6wa2eRO3xJxK9YJ04kMnF3ywXYv2+9XQpvaQwi4nWw3sz1HwE8uf8JYaK/MkYEJFcD3xOZVZj7
XujRKHtSh3frg1XQ5xBlTRngBPVSS5Sqprxi6bqVSomNgjDZBZOVFKzCKVreLtu7aw71BANJuweY
FmWyqKxY5n60Q6U+i3KqiKQ/wDeqDKT8TIR5ehtrhc1TNx5oEb635zmbJ9FThz9dsuzZiQ881cg5
fHMj5jkH3Jlz0T0N6aOBoLXiqVf6i6y+byXwvgSCq8BdNFKSuOhn3YKxHBsT9mulpLUtjkf2HN5F
zK/XFTfvMbz4rQOworLFKI1vggkbkKJY3mJQ1xh9Fndyb0cgvskynmfkDXYSSBMYkYfYRi/KWTOf
Odt2oa5afPvjuvxBwo8iiFi9/5OOBGS47tkf0tzvAlCWfj3Dl6jGfnTBdIqKUESoFNQggbpNAJKX
zVevkzYdPMf0griKo4VcKicW4RJvVKHWRTGArxe6tUCN8PsXFm5sWWz0P46bYgQv+nUsIqn17FO0
1lsAvpyoMH6Wz+Vkq1I7TtqQgOinQ/awoER3c+1PaeWdG0spYS1nG869bs3LPrP7CBmpZL8D1Y4V
OmO/rxLVCIcZYG+Gpm4k4WMuQshzIbDol+f2T6SZsthP8hI8f9CnbrU98aSOoyXImigIjfIaihjE
SC8kP+8/fSGsXAzCZFv3JftVj82autLuKuus6IXgTc3F4a5tHplutoD/qqUcs6TwP1UOLnOkOVNK
MFGNDDEY9hI46n1fJukDkIt+Joa2TlO7GbC+imqWZWTPrZA7B7+ybByDjaaIt609cKj8joHfFvxW
skTjN1+Jqr6RJEGYYqIJ1OXjL+JpScg5G2AaS5pLCZel3wkDxf8anuJ7HH0cQZIqIpf6dYwzCZug
sk5bBF6A6xtX9eEecNjE5yw4cN3yJ2BpTEsn/+LsIIcYGdIlefYBkIP3FFJ8P5j8+4QJQ1CO1l4i
Y8pN7Nvbm6pBTQDUlRO2R0kv23XJilA6i0BP7BpahkSOmC9HZ/Z1ddIfDoVvMQL9Cxv5s9rTtyMM
1Yivtc4hsevHSSzTVKcdldmZQCe0LP/kk+W/jctOwuEkQ9LX59THcEwT8Otrp7bBdPtkTjuRAwiV
rdKKQrQuEbHtmnkkIiekPb1KfscYXX+fQafRZlntva/HHClzTOv2UsUt8h+oNx7KWu9Ne+4DCoC4
uD1SlyzuEQ3QVsiwRYR+Vt8wikZxXsND5hZ/VeIoXMVtkpOn+CpisGy0jm2WCWfj8zSZYcJSD/J6
dF2P4hRX5iF2vxFiu2S3mWiz8SpxccLus7QRTMXGRhfRmjBsbgq1fA/lpddAuCKEMRUAkPn3KGFF
iFQy0lS5FF2ND73DtiYuPmw9THAXLoYo7SG1HHdSAoXksN6sr59wPutJ8ncwM+vc//1CjMlPscS/
i4xhs4AdsdKu4H+efcKiy92avOsIDrjD0QriqARS5dESWFxUspfG9RuTBYFQA3znLrIoSDcYyMcK
zXow2q9bwiS3f65nBGj6VvlA//UdM+wmin35v7vL371Z+4+iBU1NIQbf46Yy5k4+1VZDfuqJOyrf
66vclXrI/u3c9WVrIN3tL5lnuoRx1y8KiXgHGSV3Zr69WypC7MJKm6tmQKjdx444DH926iAfTSKY
gHug1yqRabbS/21HhMnT+snINa3SjWIqzVK6VKRSP7MFdIX21BmekRQuChdvoML38UVbF3AM2lAd
uNP50TeDWjppJEe3p/mpeLlmYokrjj/eVyuXDjqd/Znp7Hvti7yX1+fveibaNT3DmqajkGjccs4Z
BP0SqcmvCL4PnIS+8rzTAfPMea3Lx06ZbtAuKt9m+PfgIwnqLpRdoUUtgFvoGGYUanUvy3KMfBQx
96GU83CsepUtqqIroncE2qs0qdHw1d8+yntQzNukj1LRyhSNPVVmhR/T4KkABoirfe9sWpHUk3L2
Al7t5H7cvKgtElRPLHN1/NkP4JMiRAgsILPXxyxyKY8BrYQg+6WehM4TSvSteWZa78cA3NX2R8jj
Nqti+eC1b9P9S4YhXU9UsGLotOn2yrbp3hua0DwYLRLxf7iE7GFedbthDFqpHVObUlCttIrOWuI2
SWA1JrgvsM7cg6hSM+RNOnHHy6gh3YOBZWGQeydUKRJTOaXek5J6Plu560mrXX2TwTm+aF0xCQl9
6a3ZpEkVgv4c/Gq9i1ZLpT8UWV9pQ0CrzE3UGXjtd906zc8kbqsOPjUObK6enJFtbY61+WHL5OnB
uqRoMAnqGjEGxdKhEbbD31f+1YfsEq8tG6jyGTw/Cg+6xMLyl0QAZLm+zsjYjTE4zW6GdKZPaQJq
SPH9+V+ubs+nghs4HGyOHB46cdZhlHvg4l+5aqZrxe+BPlSdXL/nf9rB74Qc59yYQPt03kQ33H15
517vdMxcRdUFOtSVKj2MkGvqU9O4XSLopb1Yx7HksXQ0NMmmgDXMGYopbmn8nAtnDJQv4v77MjXH
Y4zHrIZ1iaEuNWpKJXweZWYjBBhnAwKVC5dwdjC9+c5cqy4stqUViXc1Pfcb35aPYzxv/ypt0GIE
flET4IRGJ10L16s12W0g9CByTz+LJFidBUoeNOtw+JAkGqrIV1zW5RJIiTCprrodYwZHmNSL2meA
yscRYZR6LkX9OxZWYx7S7mX4maGG6pnA4ySxHoO31/ND63LV8dLf+UdIVs9BLgqleh98l8VHhf/2
KvYU00wKqpzmDe8SqQBVplgmwMeJLsu2IR3DJSoLIRNcj2sI0z8gva38R+PmA1IVochaRaOiEERn
kwPMdrjXLAwumFzg+Hq1cTFu2HjjnPcMCQMoVI4wE1GR8msSmnhvcL1c/442MsO6164lVwNFv7CE
fEPb3OF9TAiuYx30xFp1AE3rqOuz6AlxHHYYdGFGBx5nBEIUNbCFcq3ny6Z7RTU7WbYiukEW88w0
N14N2CLzUgTXmtPd6OnoVy6j1yagIN3Fl6ki3350xlHNGQlB+qHNi3Y/8s+nXtnCJmbHiR/IWkTq
Yn9brI7lobBcAHuGfq+WWJYW9qPvSimPbNQpA/YmgQQRvTtsYyk87n2MYE4il4aZ+dKpENuQJbNb
cm2imPuHua7li0pfsCcxDY9Ywjg0KZl3Pil116J0iROJJxIExEFqRGglpMUbqmk1n0htBT5FkSEZ
HgeiRzbpEw1eCYu7WQGhEwxpqtugoOFU+lEmxHvNzbpoJHUzSXhz72COy4mf40EcYtCm8NKYex6x
bAodb/kPNde5yfNaJXTgP2gBwLITQLbckew7GUnz0zmQjnOiW7ckk9Ob2xLSFon6YSI3pKjHdjTz
1AIOAh/nxW8eAm/aQOPJp855zsU4n5C3G1WKVreBVCsSGQgliFzq1aqFWYU0z6p+LG7zrW/MaiqE
N8UE602d8N/V1yTYq4Mv7Ehyq6Sj3Exa4i9hsUcm61cOMkCLaK5M5iHnn/jkr4Zgx24QJ4Ptn6b1
KxGZN9zf9A5+GmaVd7aIFxZQfmkZlgp5mhdVC67gFVm4mTuHYAyid/eSWkpZap6Qd5xB/+z/SEzs
nVbH9ZHe5qSKQImI6xa1vGQ12owiXnWGrK63OXcZcvl5jc+Skusg1PHuT0ikQWW5i4Ecbb5xqUPy
bscAtoJDRsINWmyJCqxa+OGGeJipIypWUabbPaNSLAp1zdP0D30MlrMYRktjVmyUVEt+6q0JOfZs
FX0+yyTi3XycGLtJohQ3ibo8TFVm+QiR7x04lQRymNWxVuoV0HhCKZgHL302jaHnkWmp3E/lVbV3
2fn3XIj9csvQJyqIcxZ7ZFMxWhl9MJUcjU7W0dJg63I7CxH6X5qkZsMNSN9fWdGl9kCi9yWsCSao
FCXcg0AZxGznx0gEF0OStVEyB798SZMTpAtmkUxEMFpuNxmPxmD9BrIPv+4+4FIiuqp2SIcHJjmr
2BzrWo/VgT5jY/dBvLbLp4Yc39vwL6sfmSM4gMMhQcjifFX2sbrI/AB0+Oa8bLJ76B6yZ0WbXDtw
rouMpHttdk+Om4Znja+rSwiHukE5nygkHVibCmwErqlbAtBq7H2clG10e0L1Elw0W9C1sLFEWvGK
2GWuDHuRPbPYjjIWSUf0FfaH4nm99edc2QZ9/h48yjIRFvI952uQ8u42AaB8e7hwcjYmCnk39f5V
fwDXXRDiR1jKD97wHn2l8zfOgiT+0rGagTlZMIwPbCvtO4wCk7ciWLNw/hayqpHiV/Ce9le3reQH
cBv63yTnR12+iwfxlADjB+OcigX3EbYZEYvZdN1OSnmEwRnxpZi49RAvdONNj3OwW+yD0kaSjwOZ
rEJ0yEkRyOFeV2NtxSijnRkUwlWFJKvjeI2KCN976bQoj/VhndVTGqwLJxoT2d+IzmIUlKkoXb3N
cV9fOopcPzVoYO+5JMMwqi7QBOhSWhRfaxvSS/H309SPd6XT925tU0NJwQxi6B75LkV/9XsO01Tt
ATBQvGVdALF3ihTaaiS1ddPMwUXF84N8rC/XASvTyA53gYIMnYwX6td3NSyE4M8kB7CzsLJeXRRa
7EU7RbTh4+jJd+4tkH5zfcAlwUvz8H3uhnmoTNw4P/0fJtuR9kc5E0vGljKTGRwdIakczOi4N030
FSvUH5beimNFVVFsRWR+JVCUw5p19TNZ6DnGr3S8SbVmZQ91WlfCdj3MlNBNPuPgyjFQFh34lJ5g
Hc5+wqgRXiJGcwO+bZlrAE4bm1trk3ZwdGAhDK4IXpJ55fRX6ua2bNYmd8LZZWALKZxS6XQXBMfN
cu6Stncds3J48fWCVEVerejAIZ5LUM+Gi178OBJzPxhAW/6op9XMA03Go9BbNUGAZVGzGS0RKFyE
lN9jizgvSuCvYQ7UYKutGcE9tGiTm+GigA1mpb2tjoyYkTE3Qg5LhkAf8rMbDCXRHsVVjgsytWNa
LP2guwxW80ZFtrEZjGZzwnpRLJ1HcmwvrRfXJynztHaqW7jNk89OFQtIp08rKvRz881eQoaFc4m8
F1PUbz863CGXI4GlLcCpjbtlSXncYg1uJtrK1B0yy+NpDw/BQNtYekh14q4+yT0bMbNVRlKr8MgW
tsmW3cnBR3b/1OzO9sENBWgbWLeCwIHw7qhkSPhT7cDWHiaJMp4DeIL/A8QD+4I1eYdOf6sstNfN
BjP+yI788VMsoQC4UYjVrERLvVgqlRqj7gqNdbpqb94Zs/dVYLuc43yvrjn0p5/PEQjdspffcTKV
SfGWGkj16YwIm1xnYbdIf4XXdgEGBWqjvMLTbWCSv/4o3vdPXxpvGNP0UaRX94a9wLHDc5iXaI5O
CQy786QfIvT8LxpQggjXYbNbH1v4t7RehoIbNNMYLn2or2Jo6EXamVgI1+rKHLY+QkUPfGiVDhHe
wvGXgiviCYotj203chjc4WH8yUgHzciKJPSOdrEp25ftBTvrgAJcjyyqsh6wCsusld6iN0/U/6uJ
LR3BHc6bsk37mqHAUJ3CGIx49hp6ciNphneftZz3AIF6oGTC/ZpDO7eGL+4rxOHA+Y7F1Xdr2F+a
8gfS+3SDGNBqW8E0A6RiXTg9q/LtAYUpcWHjkwzMMfnfeKEQD9BdABYY1qH1m/ZJBC/zjyEAuKHG
VhPcMU7/vRdcmgPROULwNu5ktymlw6DCx2UAdaDn36qRwHfD7ZZ2cupBWWUdpbhWoMOq/E5/tdWg
F09erDCM3PMeRoQXDAZ9FXFhrjokL6PiLUAboyG9umh3iH27IYup1ujwBi37qGzJ59rn8hf7McQB
HPpKx/ExOAq3uh2LsFyRpCeEcTPKqJvr0SyLTYqn+rE3dgjwkxQQEtkkL23WBPJOvBDpcxAMJtmK
Iu8uZYEV76QAbJaA0JxVa32q+6H7E5YOJJkZVtrpBT+8JJCZQj9msMEkjwgKA9Q72DoX1VrrRy4e
MgSBa4pEqEPUk+UxQZrkbjKtrRacpTZC8ZuHNh+z8w2CY2z4yPMsn3znWmhKD56yvebMf+s8FXSm
WWFAlc/p4K9wt1cvxv26+JtYHABouM//aNY8TP3i8I2FeYMo39vTMe/ZCdTC5P5G0f0a/QL6UNzv
rL85nuZP8wBnACzV/iNzVtdBfYunXkYI9TYGNxPI7FXF41BePrHC5umeQMOwri1zuLJBAihlJ821
ck+T7UDYCfNif1lXbQ4hJQJ50FElEvTk3oTNhlGaE2iSDLhMMewA9jCz7SMg2MQy2ozhyp0DpGji
tmRS0R7zKKuHSiB9V2S7vzf8Jk64tq1SYpVDVcE+NhSxvQulGx6OVlxeJE/Fpw0gWHioKMzdf3FE
6xBhqlo915g9friVhy3ZS4z5gA8CiacaY8CHcsZ1L6PBwRl152M+EMt/afXYc89nSVZAitefHseV
eyn5ikG0WM+BWipcx4+7mbdHGricAIySvOPOgpTDLR3kN05bI1GZJJX5FJVyrFa+EYtZdjEtW2eW
hud6mXmIxa7niCEroAayAZij3J4DR1uPq9IcwYYVmrbDmafAVYFDAN+HcrtGwUZ0N3cGL9hmdvj9
fL3MtPw4OCf8Yen00icRGNsXczE9Mizd2OtjMNIS3QUYgCXoidItp94YvI0Ny+zKnaRtW+26IhX4
oP8hqj3OVKPnu0JbDeFTSgvCAcehhWYNv5EKXRestTrIe+yc4kZImaHJJ/IAFmlTAey+Sah3fO29
0UQ9I1onzEWZ9V4IzMTOZ87i0d2Ca6/9y7SAqH3xSkvqI/RIhdENqQSmDrKlzEs35tXmBd7Y7Sth
M6Ibs4uOe7TP+pachkYziaH4FhRgCWoNmeMRp+CtQswzEMdERgsW3iGo9Cr+cpO2N96vJalAD5Ya
o+cvWNJNEQLwaEYLUD+VUYm2Yqe856mjWgnSEWywQgoUkJerKueXzOrtNa3ZQwwjPhLF01sI+xsj
kgrEa7Jms0cq8N5iwkQkhZLnNR+y/6XDWh35CKTaP9MTzO6egN4BwI+1AyfWOs4b9vO4cVemb7tX
0EEMdMPkJL7eBKzktwVfilCdbXCBP3Nr8YDrqyiBTRGhpYrTPyDEVE2xsz1O0fhdYFe4p3asl4hF
jR5bcRJeOMnc5Uhxe9pkS1m+VgNp7GWLYktyHaXMU7KhVOG3iyJ29q+4+KRLoyDorQ3+EX8ioYIo
OoViJKTsYNzA3kKxkX28GNuZiPRDhv78c3eX4pp22D69lc3GDz069u/WXVHRwMRZlivtFkDrwmp6
RpLaLWBDvs3I5x5KojzCXsS/yXyk8BJbiHekw7Vgf4nphpYpAQrXRsXJ2KJosrqqsin2k5lNaAyo
Emtm36PIlZ+VnElwS0kF9j6Lw3R3+5YsaiZShtwjssWeLOnY4EwVytI2yRQIMElXrPQg0iYqiDxf
QYj6Fyos5BersNLD7VBxdePxaVvOhJjUNQ2Czli3YEA+T5AUz1AG4KLQgX3a7WMGTwamfOzq7e2E
64GX2Mju74QtGivwcGzL7eZP7j+l5MdgURvCNze8jbbawL8L3DGndmfH1ngd32nwSVhBZC7aus/A
X+JUbbhQnJofbKg3uxNqReFunv0pq7/h9orJFtBv0Os1D3uvnUScyW+FoJKVmUL+75o0kDIc7nw6
mIAV1GcV+3DaFVjSUCDMMiKR3iMery+4Aqpu9tMmQSqC/eAxOqgusQznbhE6vfl/JJ76upmCRwAd
WoGgwLaChvrwisF0pcfXhVxtC64gs8nOkF9l4gmQuRIb42xcpPqrit4PR53xXJzx/RfFAoNa+R3z
OmaznUDx9juRfXKdRxwo7/2fgQmmYLFJ/BjCOjLJcW5wxwkTJMygsh3YDPFcu3gfN/lpCwvk045P
5YFrHBRY1qaYOtDLdBsAtvP1mBSUdXyACYHXqSeyqdfKtazLnIiYz7TcN5nxX+o4D2hKPSjOekc2
yRfuDYJ41TJEbMSfl15BlLfLXNkvhVBndjTMCP1X9IhT3/6kWp9asIaT/olxBRrHpQMWQuRvFOFv
49pJMInHi5f8h85CuUztoNn2iO+L4UQWVESPY/QACHYD6j2Q/RINzD2qiokn2nXt/N5OsessT7oi
kHcbhDdiJf1iZn87oFZ5OUoBLlKIJfruUAqkLjZ90v1nax3gFjlb6LGQgo1Y34ZI3XLquqkGWCFP
DRbtgOtxXY+Qym8OcvT94nAzmkvISTmD1Zz1CGsK4QjNpI1wPX5OliWlgEGcNNXxulbDU8frmSCl
sGpHgGPCQnOQRNe0FE6W9MlRFOOuqgzcHkVsGyfGzmOPyWp5iWhlgZJ7qDmj0UfRYpqQPkxbNEPm
5GVBtPxiDlLDOV4AXvSV9Qk0miuyGP8wyGpY1yDwCVY8wNDnoXUkMBs84XeDD2cTmfpTsfjVRiPa
6M4Vldrruj0zyTh+67T1HDYfMjj+rmWH0cO7HomV45ggYhzNzcFhSH6+RL+lFZCX8A3JyPIlxd4Q
ePqM2c+XqjIGYdQ8NW7TlyfHDT3/gRAmkgUe090zzH0Xxgfe1bTEyv/R4RBkzeSoHDQ9G0AUM914
wEEANNPVoA+RoPXCp95sOIqTvUO1Bptkdz1I7fN0soHs7Pu75vuE9hkbQuSzu3cjvPsD8Q5FA4NU
1cL59E8jTB7yKDbqVzGp4ciNKTuC429DfcPyHrhGf7KsFQkJVVIUbbzqHussrau37UUG8b6CD56E
UNNlN2Zff4pRHLGx5XBbmf6wlnym/E52fFhpLBGDsmjWFkBCwTOfYY3Py2c95sypeGs17N6ivPp/
jyYzxw0gHJMJF29TqapWjusvU0PIez/LKdZwj89vHJI7RZMV4hD2JOUUWc1YL0GeqAUijwwQmaIw
w80YqCHE0eyUlyMrJzisLqSH4UQVmv94dCmgCH2o2Fn63JYbv51RmSQofhLKROLRnDLLT3LbFp6U
CUkAWDL0i0Ko2QKhyq29BXh3Yxoi7gIWvA6dPskC914WV1CGF0Pot8C6C32uSl0H2iU9SyxPC6kQ
soSPv+C0orzml7Avl+rlofns5e6bGKh2VmicECh2D/IFUXoxdMlXXwjLqSqzmtkFpOsSchpuUwXh
ynM9ERLkk4yCHl6L1C1HWqunTtWEUIxEaW4h+BPSuW3XAMYBPY+D2Sn0oTwQRaJDkZy7vaDWGAoV
IzR3onmZhsqZeLYpVI2t5mpb4LDg8yU23pc122PLWvEtVdZ92P5zWqxg0XmqezaeWS4uRuaFnfem
meAFeCkAUMGeVJzptyxt5EnWJ83E8v32zp0otDHPIP5mH7FUoFHCX9XnqnqYHxQ1fWa7MYaU+/Oi
Yxs460s4q1tuOIVG1Y7nvu6q1QUhVd/DYJc/dDBytDfDI1mQUbsQjf29eFxGZ0O1nNTIbQUVJM4R
isX+n//RIOKn8FVYfsYNdyGix4tfE9TAqFFl/Ipnjryp8xN5FjYXjkSMQYsYLy1p+3iRqAC0VD7s
Iv8NG0EH0NdszjJJLGDSrBHCEjKAGUBYs83DSA4mnXplW2gGlfPX6kxJRhs+UnBF6nneCtJywm36
ySFdCp/MTD46pK3rSzOmLxsIC+cdDLPEE0Z0sDpNP+EtQvGNAZNux8ZFA9p+FU5wmGT6lVNkszjs
hf0CGKAhGxYV795mdykt7DBz/Ifzsw9PeUz0nhfr3Bpq0Ud2qCZgwRAk6PeQD2uBQetQUj4qKzJ7
4i516hIdbczzNYAn26WtheI5axLOJyhib0IvrpNKlV5NBaWcMsOqRq/PUsfCQD4maL1F9jqr5YZx
Zw1B/U+SM9ZDSOsMbObu2kMV1xc3gRxtGM+eGklCZJpX/XFZsI+2GfZWxSs6tMlvE3wTtfxbUYRH
xEMYYB9+UMh+GXqA+rQ6q48GFur6M9STz1kQAXX6XVt7EwczkUWLiW8MX3tF7Kog0z5JBz9QRcUa
Yz94/TaeHr4de+IsH2CUrWgqbW3dId150yJ03NSDkx2ew2HulYnTn0G/4CyfEBIn0hV0VO/UNkrI
+KUHV31pjyP6qP/Wv124H1P887m58LrDuXu1U4wNHMZ6+gKO/tMJFebkucZQnqL6vi7+4dKoHRyQ
k+LfyE76mYv+uI17kPas+Msfey92Qh5/kOErGSGfmSq/dIJkz1XMyf5r4yZ2EKQ97TQKUAHs+Trx
mVlWBAawIRou/Mc3X46Sw5LCZ8f47fkUYu0u5P0sZ7t4lTr2fKVf2T9TJ3oE26T72zxbjlRAXBbA
MhQ8bp32eMQWWsb0NBdkNv3U7h9qCrD3a4pgDDHDwueG9WXv5c2inQ5ckRx6QHU7OYcrwHQmbYeh
Hmw7xHPPUhmNfJBzhCbNG4XVxGcN/ft97EI+PuxsHwwWg8I+pobwf9WYBPUlVXrIxzXU/PUOb8h5
FHfOWFCmVxa7DCCqvV/XGBJEbCnFHGkjTXW50XeuDTxYYce4ZE0Xt65meFVbV8ouEW4wod4P7eLO
jTGxQDoLPlNbf5dotH5eWoWyCVoTnPrBuEeiw/i6uQ5COA0VNgci+m1oR8tP03JrSszdmcti6N6p
budQNvuACNYuYZXiRMr+olzGGh51HzJ59tHjlkLoaA7ftoohZiu99/Gj7W/NooWccOK7beM7d9bm
yIWfhPDFpcOlJe4nUBAco01r2irn5PdFWjCyktoDJD8y8s77X6NjOJuEzXb0Ycd1LyB04tgTaIs+
j9lueXXvL4W1N40V3EW5FPsgpjVDl0gsW/dATAP8MF2YmTopVxT9rdVl0WT0XWJ6UHr8kzk/YxF6
K9jvnZZB5iv7VRD7iaw9UP7dxK+Ym6GphfwihT46J7Rx/X9u9Hq1kC6raXp4jbFdS2RRQZoIbsSl
PqO2YhUoice0GE0LvEmTPgm5HiXD/JATa8W6pkahr7NURG5v32G0V9DNJaqHJsrcPrpo1TRQyHzB
Dfah/RadRYI4lRsN2h1SC/0HAAtYQoSXMS+bop3HihVcoPULN0rZlP+mSsb5L45rqjruwpkXjAbH
6N/qbhqXFMzfzsp6liHw3m08N56LnU5JkTaghGdA/55uc+oUbXG4xRkmoREYZMjqF1LWGVDF9Bmk
yS7QkdeKz6R2ZwoPWZH1LqHDnhmefdTGU9iGaS1mWXykrtC0wzxHyjBqv4NSu6bj+ENXNh7gXOeU
hIiSEMYrI7+Jf8AI7iHtrYb6o2nIZcm+uECOM55WOZJS744INKlNLldmiT04OvUiJjSPhvAkXle/
+J7INUDOJppyK89SN5443+FVxIoBDcRpqn6a55/EkJEvKEASHMBv1qYQya1znFbJrhvZwRzlgm3e
6v0/o8TESKPgb0h3Y8PMHDIita+W+7trEqnmvb/r0Urjtu/CYj5CTsu18iX7RcqJ9n98Qn22GIpG
4JmMM+YGLElMJI13LxovwjN8XZ5LZtEl7T2iSgiwJCQr/4vJbCplmjjefZKlipS8o4yI2GoaV0pN
TQ1vhM1p5CgIYPhiAqJIhvyjzjkJ0LVnAFaNUYASUOrQbg60cZpsUaer8Y5NESCbL3+Rq+FIbU+3
iGd5Bn8UOPDjSJv3vY8B3EWyiSdCljNuTXjcI0jbc+HpVIk/C2BDyFY4sE6olu+ju0jYOhnqcTXu
mpetpUUvrfitYyJyvK/yF2VprdpDJf7FmSMpPBJuAhY8Zet6IXaTIvqueZ7i++rMAwmSI58vCUjO
5W/jYN3ol16pAGkkTyf0xR7Psrwm1Y4OU7fOYpQ2xAU6TpxhXmry7+k6c1VwrZP7agGQteucM0/y
AvApCRICA6RJ6aP8I3rvBqpU7m6d90loqu1CYBFGPGr1ZXYK9Tb7qVqfyw4RwEnB7iUCKIJIZIYq
vUO8zEctsyh70Bc3kVWBpApuMalOL1Ss4SfvDBJY4pCdDhMpDfJghWZLpObqKOqXJ1/u4Htz/drx
7K5YabmWKRtcF+04kCkkpKclIU+NIk04kmwqqJC4OKsOjHkNFkz40UT0Z+4Qfcd+THS76lV4Bfrp
lqkFvjqqrgbiRjMNrbfTbHAcZgmOnEch/5TNPqyHnkF0dzFuUMNrE7pjay1smHolzaxOrR326CYT
x+AVCLchZZ60ELTk9ykPDp9e9wThooQWJfmrF4PFmDSkLNXKA+gPhxKovzNgwBroeyRjVFCFXC7V
9VomsT9NDKcnwNgpGI2pGOAs5cESgD/f6587orDHPjegP8bDGmEAmPhAFM3vtXYV9+IqlPiWd0R3
H1aFTvmopIUM+vQrKpDVPXK5mgdzHyj/LNFhb9ekEbIV1lTQERfRIW4QJAQqNggWmkhuj8sMdApc
sHn59tEzXC8lxEtZXbjsnc83jI5LlSJIWsgEB1fAq51OzLyrUmS9ffR77RpmTI0cKDErUi3H/9P9
N1a6CLXKfDu8+h5YcWHZRLcCftiq8VAwyVHefYkKn9ZiMMklcV5qlexQyE1cKPn9208Vl8JiOeDc
CGRnRojuWIaL4x3gwQ5d05Ug6rViTIeW1SGvbdjwxmk4eAJoUXX9Iqw3mGiPyhQPhrMf3/xSAKC/
Hopbv96hVj9++hdWXc/4ZzfTDvGr20+4SOG3JnoLrpNVI9+S+FEKn8Yv/PD8xfNQFp03ySRgMF0T
3svHJ5x+sRPCAUeoWGSumQ7t2bQ4kohtZ1aiEDDGxqzx75yxUJdB+/r15S8Lk1/K3rrE30M9I3a5
xTdcJ11DN8DHE0pixR5FwUpjrZIhCDkI0tSzD7BxYc0Eofqnu7rO9l7mL869GKiGD4WIMV6Pa0kT
DKMxd2iATBmdCG23FDGV2T8sYVGI/2jRAYCTdF+7DUuIGywWtgaukzm5xE+0lPwGPn9Skc3yw6WX
EXcqB5YB2qLonb1gVG6cB1PscCtQxTHU3vuoID0+hFx0XV+ndhJ+ebsONHR3fbcZ+eZHAQwPYrp7
wu74ltJqlZ2pAfLwyJZ7zP4ex7R8zV7QH16tccy9VYMYSueg4clsbiBzvyLG0K+IQBsLxZ30DA/s
EjL/Sw3umqrHziRT2Sk/OY5uSPQ3K7CtugAAZaVXldajLISSvLNKBU6lPqiozqrcHoRkX/B+aYHp
0G2FxR6mTnWC+ukt9UD2qOvj24bCPtKMsdiaYurI8i6MPUOK44OuqYhuh5IHQcrYQOGDg5IjY6Be
AMIGRkGq2aHscI/Y1FOFxbCkemnTG1Jq2rYuPERAJTA2jv/Lj9G1JDvw4IiHnvqlM/iha+BlGNYV
ZLQANGMDTEOISmEJCXdOPnvMarxSEgI6mv7zUg28MeYHxmklcLgGjx36ou9RMAD65jic781SnetC
DPXf7VojSQZGq91bPbWiiXzqtPtkvgsyPc5/0YIUpA30EFeFbxOqbGnErIq1XKwh6/CHIdhivafm
IRXvv788YbzgPSXpjPAakriSrRDgivuTpLIEUGxEKdn9JjXu48pgYWu9ttEVPGINaRRE8m6qqUUK
nbPPIUMcNYZTR4DY+RuLxt7RewSTmtSMMoVepkRbeK6QBb2WuGhA6M1D8+ZKFRJ/P1hKFXThfW0d
szLHWTuG5gIN3+e161udHJ1ZenZI/5WncEkYTdeot36I0o9owdIhLQKlMmD5/qaHtNTikL0cPJB1
OTM62VzSGZWy/7Gj1TNd10TQeuWtVhr1bNRI8ac5yPvXjI+qWUoiz6lmdNLwb1D9U1IJ3gGlwY9q
vyRCZYQXmqAkZAQY7L8G4RK/wt5PjeIc4hlwNpRN7pJ+23sPTbkPPLIBWKujExOHz4QtMuJdLPg0
Heu+8CH7vkiNcFaZ+K7LSYoCXg5sYt1pHPJ19WKGZB30WHC6nXgXMxtodG4yNcH5I8Iezr8+WXlA
uCxk92xECrvhLmYDOOZRqGLRSV6AS+V5kynlebca7ZWkt+VPb1sGu9MwwqRHz94MarmzxnirHK9h
MeQsXSVTkT3YYRKUtr1sehMuYCIPU4Hc0WR7L+kbAbWL5kosMG8Iw/c8qjG9nd47wcDxRzzucXdq
aBmzQN+7aXTPx21W1bYup9K0ieC5hp08CLq4chsv+br6ktOeEhKMwoGEmRBPYmIUHOJz3QIElBGt
bJBilCBU+bGBh50QEb3aA4cGp3wUU8q510JncA4+WEk+I5VBDwvUgGNkfVJwGX9O/cNxMDmtZnux
t3Xyk2fbpgszMGhIIRBUbGvwo6Vu75zClekgy9G6/KJN+LPW4XnQDJXgQdt7XHHWEZ+BFj6mbLds
kz0FXu/KO1NibeXFMXn6H8I/+6Xjfz8yn8Wy7Jx7d2nzPOeIbPJKAULmEPWBtkGC5H5woBGRAjON
3USaVUlynfB/oHEeVC6QIK9ZxWsa0lDDMw5PB6sE99x8dREhpnmoq0cmx2dK2b0yBifa7GrL0eaT
librCAY8xJUK7vksDX3Ghpjuz3iSAOKHiPocs9epiA6JGzNwOg6EtwW1wiksoDOUjubGGzBamBYu
U6L/zsV13snQfMFzn58q97G1nL64RHUDGVZzR1Xpwk18mQB9IvOHGWROoXcG0hn+s6KNfXl8h6cm
jDVVVnkZCbycaFS0MnjzKnI9mSXJH/SYCofe8qsepFCOIMMeIK0g62x9ZK7Y3N0gN88Qug5UAdPS
MYRZTk9RWfN64XcttwRByNH+0jnQS1/yTjtOQ74E/Lp28EEaBO0V+Rr4ctilcr9ml4cTwcMApnNA
ph9JZqxR4U3Ku8hFJWHvOfetxvuCPTPsn5ZuSlk5giCgDLVJxegMoln9XqqSo2tY413LpfLkRiGc
/QkdZgK/fkJK7eHlE51NvxL9cP7FbjFdjzW3/4rWYmY8Q8NpqhjT+1J2OctwfgKYy5ERvX7etfDa
0tX/5qGjxF/uTSHepSoIqonv619vySuipQqJnQLlUq6YlRSZHN+UCcuPp1TY5Ne4TzCS6Fp3zeo9
aWXioib3GmMhTr5LGvlILJ/1n3xh3niJPGRlnSHYDsK7wllIOk/yCqKzTqRWtQB1amyQhKI2eLae
AvonImAKwB9QQIzBfBy7DH43li1dKOQLAn1X8FHeej+7RjJb1WNnCrFTK/7quUINmWl/Uycw4i7P
Y2q5jUZXKdB/PEcJ+wUqOIqY2dT/MWba/2ekoWhFqwpQ+YWNj0jXzFSulVY7alDKBEsfF4HJjMoP
uNCUowE8/JTnTIpjGf2IwZdllpUxnPK11ToaYCKkPaWBmNtrPBoQbj5qYgNXhrCeOdO1Kx2ZPSe0
ZSjvCyXHuiG7vTHqExj+0OIhFGoFpzZnQLXL/+ighWt95MLsNwN53AJg2BB6SrR4ySzCCTlJyn38
I9Ug4tUE+vMKH97e0mTPNpGz0Tmr9tPCAIlURtjt1bPlq05fbkhqcEASYEFR25lc/3N6B7xi2RK1
1UgQR4wTmLRsfn8NM+0Rck0xXBO/10tde5FLF4hPeZ7IPJWHuZU5w0S5maKeV508jCDx9x1QlKo9
Xq3YahNHquoZbhqi4ADA9g87DNWU+Xu6L0XW0cRWDlrTK69BACV6NngHTldosZcxHsSRqBwJFoCr
CtFl7QEuuWf/+bAJpJDah2yB8sSkNERqqRIX/RD0vLBUcZM0PSgNR0V++DMYGx/1TZXLBQScPbXs
Rvc4lPm4J78RmkKrxjoM5PA9pKKYd2c6PZwaca6BdYrFRyX7BTtjDCA82LkxTIR1VIavI3nA7X/L
QMVUn/Nx6qVekyD12mFKAU9JIT2Dtv6P7GCTHdHRCS+Wv4qV2gFxqa/tP07jBiyWOvFFQueUzUMU
nkdbPfjamMQ6rp1e8f2Z0cm4Zozzcns5l4F9Tmuxy8LugswFXldGjq48nSdo8vld4cOt//4MTtgS
Moey/FtA+zV12yi0zg+coZVvcsRsrQQvBSIKM8pmd7+7gIiibdBdBOL+Y56jvf/ShVnqJX0m1PW1
Pw2Sy5Bq5IeBEGFwvfvMbfwf6Vp4jyneugLIOFF1B4iq6J0IEzra/qkr0hSFuFWKdOwvUcr/ZIoq
IBYv0fnWWI2rxJ0QDQNvyvXwbXCFWxxy9iGzmEbg8Lj2SzKwGi7OHX60Mr/2GoQ110k6zBoyNh4L
7OXd6442wzlH4Mf2d6YKkrT30BfjAzwYBPsS6M7o9sNdZ04WIm1GRUwkTxgRJ05UNF3aXHKwX+Jt
3HBUCv9j4rztWFIjH8JIaoloE/UVwDRc8XLu2n6vI4Eena/SGEQEajEZ4R14x2tzSSFgi6e9Y0bo
pjvtu+NjJlRAwzUesom+BDbgaiAdtcRWiaellSuRDdunlnKw0oIBdNrVAgvSaUsTsySoGXuUkxnj
qhfLkvhXth3EMyD3I7o8kaeSw98hpxs3faXRSfyZUWrItP4VY46qkfx6tUEk+NXAYS+nPyvwZIZt
6/Tbb6nWO1I4nl7mqzcOPyexTjInDfrqH9pNSwvWsnbDoOOua8t7Xh7P5PehN1RBK35AFN49OPSA
Thx5S9NwAZjk9SfnV9SWGXOIGuPs2qgIRqyuIiwJkfxImLWSdOOYvLEyOeusqoPhJmx1oif/Dkyc
kIOeruK1Ca/gsq40z2ztVnYGAdbZALrPu1wdmHlnQg0FZ1WiqswQZclecVKZJBLsXnHS7iQjW2UT
rXXQZmGkEoKMMaJaqabzpJW2jDgYAKZEAfXgMLpEyVuWjDUjrrq87dRvX0k+IvlgES8NYwOh6UAP
zM8/VgPdArx6Cz4dmtSJGftymRRbhYspBLsX9va30hPf1DLRo0/W2SRU6w3Ded3fDKLIhjaZ9I0Z
Fss6dTEEKPyEXE0NRmiIj61SbEfZKAPuevKzP5LrAqcd/4OlDQMz66UmVPt0Gj+Lil+vIQ0VzvbH
60S3P+euYN1lCsa6A2eT37Ab+aXRzFjM1OSIdZuADihjBRWvO1lLyv4tuIlFGHUWLCH8ype5K395
w/S0dTskFjAf8PgqP9smcIryzNP0L2wkKs6MRigXfFJ8BuWLXyTmi0akhcjkBfEZlUrCBsR53rpB
fiN52+Acv3LisuYYZZEIkXjJnM72LgB6Jlfl8Di8WKcSNWYQE382QHsrC+xhvGR1UOX6SXSCes6p
YLycQwhHm7JsbdbRNxY3F0yRTGEqCBarTWHjVFD7KIYLIE6KaKMa1iQRNTV6RQjtEixV68mFc6A0
rFd892Y0KB5TXInlsVTLBekjXl75Af7P1nhl0UuvkCgNgfZpD/3L5OOhvh/KCDuExgrWctNNOAFa
N2fAujy6smiBgVXPwH4IOAuWsfn6zixeB02aTWWy41/cTmLNZcQzqQtGCU1YE//0eG4Ym3ReWlVX
coDCJaHNuSdRCU7j6ngXD2J42lE4bAEI7dGIOFaYv+Oda8MsY8uPI1sMnQ7O51JE7BJiuF1eGPKv
LAJW9U2YvvpMSMiC5ooadwpXJwbuPSvjIPJ/iJEFnIdadgYXu2CFzONgNQGriJlgazWhr/6rxvQv
fPJNLdgksPK+5ybsU8Asknp4exbjNfsDLbLfH3AEfUbNGACymC977uYrbjFN+aU94UlZzHqhQDjE
aMU/Xba6pPfrd/viFQAW8/VmfyeizsX+7ef2b2/tJiEz+mcFXDxl7ZnpdI+w8Sc0fpGGXUCzMYfl
rEeXNOAPqBR/V8RRd1gaIHl/JcyFrxBX9sSrk+3P9YjUPIs2ebSYHSZhuWjnhCffIps9VqUn6lO2
J+qbow02A7dC3hTYIogm1KhjPxfZCAFB5xeQva6VOEvis/R5vyrGuEvCJsL4R6J/XRT0NNFqAnlx
6A1Vgmy9N+hC2iWBEU4T8bg3yzEVRcgyE7Rq7AoX848hhKnDiIbtE4rNXw3p3H8X2DNMb1q+P2c5
saSSJj7Lx4jFHCZKKBZatBbZezwhYEep03upN0Bw6X6fAKvidowOT+Okxzz7ldtRK1atiNZ8zS+A
LJCtNrVKh9xE54NVu8Ut8p9rhRLvUGuLxXFt+WoFj5C6uw8Z41Eb5f54JQwuI5a7UxKArT2qXMMu
G7Axyyo0/rtO0jNzZFHKoe+Lfd36yYJh46QuUUVP6U/F7/a58UFz2/bH0Qgfpc9w44MOdRtlWulI
w0ws3UUt2K65lXLUaHebqyMTMgJx5gSa9SyCVZQSv4scIk3mirPwjovumE8IFbxwj/uXmqUJZOdD
fcDcMx+QHEkqqSuKeQZ46IIK1Gxg6KUdqjiiRax9kEV55CIi+/lWk9aL/QJymAqyissWTDvyxnFa
DHAZ5XNfEmskF01rqB8nGVeZWY0t6fChQKmEFcU9w0iMR8vWxJGEseMN1Ae2EXy+jGmMk8X6XzGC
lkf97q00hTQ5gEFxqGrbwqZnj4JTdWhvUaqBI1zUELEf2eXhdxZNENpX/7vzHFg0w+tlavPEtptv
soj3UUYzgAHh0t/tPCWmKBwVLzl4JVc1/biKR6uAsELfx1X7WcbpubcUdsu0K7mftuQVzYCYFQ/4
biruiAS+85HHDavP68StEDdx3rjOwpDrDRAIZWDY4T1rgCdwWNOgPSz2eFC0tkjzS707it7bHhah
cqmdH8wr/uT8sqJ99HXe0jz+pshDu/ntoNbmu8VRnW7wXGuUGLzzPOAcj6MV6Hk+s2+MV1Ky0LgJ
Mj8NFbGluj64C2O7xPVUIGpuAXHnIlscg9ev8BQiidJJ9tvJvm9MtZPmumxcBOGOHPmlPMgN0NRk
zKW+TdY/XEyGTaROpkFJM5QGa8Hdu/9YqEqFi7DJIcDEW+5jnUlfQ9i6pQlJ+x3j2PQlBLQAGOvl
015Mn7E1JmO1fG+FwWmGrWcmaY79WzuhQN1r6izPDbvfh56aJoBXrbdy1ikPJcJZpqHzoljPPOWQ
DS901HyGqxt8YaAdmtVvjTqZxYAN0pn8RHRXxkKFTHU7kteU/rbwfmeY0uqaHGIy390+xfF1j5lJ
O3omB0mKxqDrm977yC0jiXQPtj1GUMXpyPYg/3xTJHPO3qy6sd7dqKPreHQKwjFeYsU9zp4G2NFk
QiZisEjExwbze0cPvLC4SUWmTaEMO974F0pgdUpz9u1bzXQ2MtM4RYktlDk4mBSe4hkmqdTBvl3g
nJGxx7t/1EKSuPTPfvRa/ZBnKhXESNAgLLkZ4Ppxzxokt0blrOAWBJ1PwP6iol9DHlFVdunS9d2+
Hv5XtQuydx4zQ7Z5Tjl0yDyew5TKQzxXbdu1f2jiTiMtUGnme4OcvrvYRDItSZj4RXJX0Mhqzo8l
3vBc4Oqc4FME2oQyNf1/3vB/f9bumgl0vIa+c3VOXLpNnJO7XijKiHf+AlYXapLtjPdD7QaImkBO
grobACCofwdBgUw0LsjF8JoxO4fkmt02gHXd3vaFM7ZNyNqBzSva8OLv59QK448VMKE6xxLPN9wq
C/5TMlcwgrPyF/1CcNIiCmgzW3AmreSnUTxkODL9T7cpLX0oUIIBzdqqci2haoau20V+Vusg/SLJ
aIlDhHXb4aYEApG8x6v7f6PWzL/UJItNZzxMrCQiWxgfqO7A7AlSin5jAuUZW0XU5GZV5l6Gl84L
mb3D6KT/hjVJ/OdohEAQhIe8/qqPj2CqlynE0/Ri9y4gd/wyPB57G//v44zQEihrNALDOh2tFF+4
xGSxKyKmKRDTx+N40CBw6jgFWMVqhOD60mE4G7WelcfHQwqNyK58K6WX+NGBTyH258bvYBDHZjac
cnj0lf8YP9SxqzzPpGGa+z5DbeO2NcutMZUyD5oqgUC0N6A543b8V/sUc0W466Q9EH6u0HJP4EAd
zOCEEDKgakwB4/6twS4AhLJ3icfz/QLMfawaRVj5PHDWRrcYv/OVZQ3WM06J3r/wOrBsmyyYnzOv
4T+yYK6C4eY909wjkUSJdLa+rgEJ3NEgMlGFZbz9Bd27MP7zz3HDIdhnFgcKc7Y82w4vXuo0TaEp
4KsI8dzrFpLy3YanrHcW0xzJoFh3EDETzRISdAlggP0u1tCExu1DuQ+C10yTMiyYNkN5kZjy6B4k
D29NHj4uEBGln+RPHj8uNYqG5Po/RbnvdfJnAWAMXV5GulTjrgVx6OtopgbkVx7rSPj8d1pkrRaD
5iHugKtsjxwIDDJQSIiqmQhnEy4i1f1xOZNwPV1DmaWIOwoHGszhovZD5rB6IksjvpIKY+izvqRO
sDZB1VR0nGqM7U3CTA6qEURr6VwRM8RG/ct1tCbraYHHG4/V7HI25ICWTXQ7edh1grldnn+giyah
9Wy+E36RQ6EwzBgndsykrmVbjMCBwJGv0SXTcbVCf9Fms4Ugk43L0VNyXw719m96pZa7y7Oi8b2N
Ko4MqUgJA+2XCuMlF4l4pRWIoxvcnFfKmJCWe+HDAJRjfIapAQnkTXziNqU4VkHZVJzqbUt/VeOs
emjOefz75ja1MhjYBiq5WlOI41UdgjVC0rG5+X2Uinw0VcxoAIXeOIuB0dB25MsDhzbyT6dZb7PT
T3jRhjpivJkovoKnE5FGCuj6Opdr5khe1cL1KW1kFWh3qg20EP5RL0Sq6pPqFeZWW3BHhtSFvEST
4KrVQFAMwxu1F00LseMeA7iDgCI8E5RbVZot3LIg54I0flUlqrGUNKAbiEn3ND2gw6qboqr8eaxC
FatXp2LVrL3oI7BA9PSP0zBp6dFQ/8UJTl+JXr5KCFNy90ncwuyuu3f8Wlgsivk48BXDzN990whe
NIPHMfNh0vlhKC1ObQyXFBA4CFuIj3AeRdI5OHWfc0N1d0rkbPStbjeziZgKUnFTsdGSCGdfX0eV
rt3PgDpN4HtZeSjJ5E1/vrsV03xbBLVcc/hxF4sGJ1Z5M2MiNSmXV8uX7/vmgG3Wt9NOcWCYrmy6
71Ft3x+X6S5EY8MKGFjK+WDvA8yqqLj7Dre1EQL7UmMin6zjNfmc5+VFu/x6HPiOSspPBR3zzVpl
X7OQUX0KwtDkJ3NH5evHl17ldkHBMNXh6oysnBUARPZLZnTlZSs/3KBQwzyiFz2n9EB25t5pCeCQ
dhu6LpdmsKUZ4yo1DCt2RN2RZ4i8GJU5YGBNUI3r9NrpkBEmpUXU8jYbEurIXl3+IfT/NUTIpplg
GnXKWYfAGS0KyPAFR/Zb2OfasB3rc2/6uN+M4duIV5aGUgf1XW80keQxmzc8nwKeVGf6fPRXTvs8
IhoOAyK1VNzRt00Er53HEHOntYA1QPTqxgOMmw6nee91ojVRi94+yElVpg1vZ3s9DhkLBaseLdU2
YYyp2DQhFYvuG/KT9VI1zPdQyxw+Foll5OxfrPaQQ8oRC4jcFCpscVnbLqxv02f+REjzVaZNlnRm
XxB+9RnL73dHFVxBvnaJRBY9o8HMvZJaEPEBZBdgCyPM5HbcSFfNiji9cdYjXGqyRoIayUln/aZy
YAw8dnO7w9+fNZs0TZhZnKGHi3MtehtAPbu+qMhClWv388QDBO3On4N9qA+eO35r06P9/wGT9dpW
9SYZchhMskSpooWwWuRz1mZZGiWowdTPy2kOfIsgJ91sSqKH62ixMApUjm+ttsi8Qvk0UqYGUxFH
J1VXPe4kpEnyspeFTNjPUkmTi8tOWPwy3bdwBHXdfuc8QbFfz9PdPabiGOJIMPsQJiTQucvOmtN6
25SF7SBmsgzxfvHYvu6E1z9eqe1i6wsm91Po9f1wuuuGWY/YWY7ZXH95/HzZNnPChNMhW10AjDX8
Sjaxv0Tdl8f9uO27+AIIApj7XK+lHa48Ff4iP8zad4gS8O39EyZ0B1Lj3xekTdTxmMu07tLURyLc
OVC3lTPjnnb0mLx1MK6HPEmbB+oBymv1FOnDZbUhGD/9v384bEDENtimiVVafEia8kVGXXiy6/Vp
3GNW59hvdtCoRJJMh+hJLUvoQoeiMmFu9LabqOMs21lPtn1BURoz/Aft12MKcRGHGvj9z+racMxS
Csdz4cK4lys4TRY/oislFb1VOAfTOz1JcA7G3qbdMv0qGSRZkzUYwfG01JGdqrFyAb0vOSldWpyE
OwBN3pnuqrqIkhgeW1f87qF+KJ8kSLKUIxpCYpjb7zpL2pVrh+/UgMEkd4omYnHy0DAQTJbtdUw1
zdWENo7QlbIQCKZBk5jjIy5IV4Y+JYmANcT0BqaJXppbEOf2w6lrbpXe7FX06ZdAbwl1hih9QNOP
RDScLgnAn8h5C/81Y4U0kNS1QpQ+R3ZReD0G8Fz/prkS5DXo53rZpTxraZZdId7coK+GpsUeaN/s
cCOg8aknt1jnT5LtbidKG0VpRcfNObbLahXyqoKyVpSqSHRI/gKRPk+LN8y3EYhHl55OZB92wZUp
arLphBq5NDanSFh0gHvrGh7nobGEnoqz20M54uHo4m1J2mHIxQFLAj0uR2XOAj6MeTc5tpA2kcC9
bvG7cGRpGHbjmJ6x5vzlLg2jMz4enaRyU/OG+LJsrm+e8nFIjMW0JxeTsRULF6PXFMKOUy49zD9V
spNXUkYYkfehs0hqO5+I+ZBfW0ke5XnR8ym6EPdCKxYPVaVBuk4CJIGtikDHzNDjIFtCdW1U8uDl
0dEfKJtw6rK2exMJKlJC9EV6NvPP3gHwvmmhklBgaXxso1QPqvS447Z5bg1ZZhd/IMWPOmiX01Gm
PTOVsbIv/zKFc2fG1O5AyPSrsR5WQA6Tb0pQ/sQ0kx0Sv5L7mxOOD2IMEdsFCL4+klzrlPQSds81
l19N/GCv0UUi5g6lSxcXqEbe8DZBka41PPqXjNniORiocGuDVDyHdgVqFxOD4bXevLznwlvIeCHP
cqJiGwVkjwiwPZTi7yUeTrCaLQtczz8UC8/heY95uqsUtBEQUV7ASmLIP65gkbWISaxo4LaBq/KD
Z2yfh8xSVGmDHtKsr+FYYlmm1B2yAS5vQlBivW9AdjdqboJYf8Obt/IE6As1AE5waAgy2WkwZSGt
qkDtufZGN8V9A2ooUUpwnM0eAInS5JhGMFq3VhlyeTgZSc8Oh+ygfFZo436ojSmIOI36EWopb7fx
oBbRAUx2cnw/WkO2VqBG+HSGa6W5x2KYuQV10VPrzKDL26EaeuKsR+4IFdDHXRAUJKNeZrXWmNfr
vZiFmptwicvX0k+wElp/wDs7dbVOnIP0FOaZIaS4MBStBQ2sREGbRziSgip4naUhske+wcYLlzoK
e6UIOFHKJmbWA0/fJdfy8jADN6RA5/yXEThB4vNRahDWn875t6g3+Ot7riuWVaTUeTVKatZ1WnhT
UMTn3nOs9A6qcQMCrSVrKF46xdIZsymhRyUNencfzEruCeOp4BnoQNUIWoL1SGtjFVfdUWKs8o1N
PGFXbzBxCvNcVaZKhhFLO09w1GRmeiFR3TWf9VoyoCQFhl3WfeXVGu/tu42euHo6CmLfejOUk0Yt
7nEOGs3z8riLYcu/aBIweUau/raS/Qwu1dj1/FN84CyRa9UqgMKs3n7Fqzt4vKsyJBepL9rEn3ME
a+ft6BxOaF0GCRXooKcudp1CrBzD645Qdcid4dPmDhaM70gVcjHsrHxtKiSltP+kfKRWyDrnXi/I
op07PNCaPE1GYT9+YB8sBKjTpxH80oCF3jglKx5Lx3IZ3Ff09sXK0S1lzf2D/3D1yd99CHI2FiGv
ed7Xzia3Bgpr2OXyyDlT+rvDsXZK4exc3L5C+H6OP1+fKNNLmEdCjbX9/woLry3fYgbvqvRRFWVG
C+BzHcj/l1AgasBsfZdb0XvXBoLbUjzkp1b4CWc2RjsS2XqVxUtbRZXaQe71BD9QDdfgkzFnIL3v
t87TK8qtH2TxL78SZT/Lo89TR/YXGks6IY2UwqDJTUc3u2ra9XwAtmc5PoEW68JX5kJU0yl3n2sp
Aad0kMvfw3lk32+fvCnCxtgVbgXW5aKk4AjEf6yWKO8+SK2JAl3ts/tEHio8vuZ8ybO+xupgQk7a
cJ8piy8J5TB281J5VHKuI9Xkm5jupttb/KF7zfo2s6/RQUEVMz5xfNWoxfFqbe51QCsGloJXVEdK
NIhYAnS/A+MahWb9nwp2QgEKnJWNVY0ViMP+X+StBAmMYZYk37Kt4zW5adAkmYBPqT3+3AwMx664
YELc6qNuy3n7CweOOf0ljo08uPs+kF+7E+zjckgbKF46e+LrGbD/f8rj03VrMXbrmpfBHNAACyJ2
7AyU/jPNBmYFVugjrhNC4HzytRNKYB1kRbUZBwg9V29hn9MBBmmrlVJwgAJDxxcvT8cnPDO6i8mq
F6/68mSq7dGfHUyzC8ikweoD0hFbPYP7vVjt6kpI2WFStplbdbF3teW+cPGRFrcz7GyiXGec/kwQ
03Te90NSloTfcXzgwM3wpMx0bx3xs1+mC04rNMLR0BzD3f93bEXV1HgImpBW75gfO0hhipNhtXJr
eOeYK2pFfarYYKpr8NO2iWXRIG56FpB+MLaLKWy7FmMTbuu44L5F0WKnXpdrqyAuz33/gLRfP0fh
ZRFoLG6lmLoWZxo7YrwX7L0UgtsF8XaF04KawOgrPDDCZja4asi3jucn9zDooQ5cxUeH4ZnQGkTR
LP3jlZmShIM26wxv9TaEr55ifUEIx9GwRW+99MQxfRkZ2zIxSOW3vOIeYQXff7g8ceFKyejivHI1
L3FU47Ij2rlUHchjT6p1POKzZJkYqLI5un+vuPftjiZ45vDy8W4t8s9S6FaaNVYa1utHnhFfMV5y
NgOv5bHXTzwC3lJcBd7E+AQZe6ZevNYo4OjSbWjLAxa8D32RliRBdueaUH/0h3du6ZaVO/gWXhMK
OpaABOW0AP08n3QuMZZfu+kTyoHG+MyofXjh63idJE70NrSqom48RCnmivkicb31l3emk5j7Y7H3
hVuDM/UCyvxMmnypGfzwhzi0zthLTjt4daO07m+fAy9ghbDgrFDdUWX7rvSBTYZalp2E0W+Pa8wE
wIM1UX5zBI4WByK9DyzMPnOTyEXDPf7g48YcpPB+2Hg+opfaCorWClhf3XpC9GdPSTxGXTN0gH8A
T3AbN+xnnqnDNcSuu4eiHNUVnIp28omM4sKsTgCIs+5Mh4XopVqEaU4CTN7+zQlBZyg0u5CDZUXx
CnSK7D9VUXfbf/YnuyKsivpzOIbH+QihaN72zMIO4nLH6+PSNLov7IP3DPco2wYYj22Qu3mFFiVx
Y2sshNjyDUH8LivT8BteAy33RwPP38yEmllsCIud9oEKN8OvCaGoBd0mrfZhhgssJNFgVPIq1Ua5
S7Z4k0BNW4NYnKELDJkD+zkJ5ZGFRc7lurivUzGqIslPGVmX0rdx/nZ2NwDltKJR72gv/MWQ0f2U
vZmc3IAg1vxhwmqC8x/bQysP35C0ObDgBD41uNM5eH0hqQqYLVx8YMiYFovkKwe+MOPEPpFptcP9
tSzi6YgUSBZDPoePn5KZmKjgyTT2xs8GiZRvkITMqKQOQ1ulZnB3vWBV1sL7rFB0JtkYVMk3Igfe
gbDC50In2nYBEExOGxjp3Ne96vRNt7YjMC8DvXzavk52+JEKxQRsMDfj4jzSI02cA9HOaGrCYlqG
Q2imBLikn0PWBn6HdiC2z89bGFP3iRNRXlNgX67lySnuhqKeVCXgvpWafdYySoxy8fD14z8TVogH
YnvqDS4OGa7oCF3VmJVKCJQx8zPsLe8q9BBtcdtvndEl1kUnT07lwkHGEEecYwYPOESL0njXqObg
6J+FnLooqBi3PoNtgti83HkPhqy0qeKV5GSzX/GWNpymtwaz6BED6NcyUZeQWZYwX5kN9Vw4ERZH
NikDFpKrThCT6pT1U1hpLrL5z7NqON2Hc4NdLAWh7PYky2VyvZzfzLGyMQCbzdvP4CdrR1BEHxnO
yjor+Jm1QO6VwGLpHjISWcauh5dKLcMXS1g5sD2fBngLs8z53x+Yf39GRV42B62Etn0aj8B4y3dT
HZiVwbiaMsPZnb7mdOLgvtT5rIe/oazF58AoncS6v7cF6xSPlzrwplulUby/wFVaOMWviai53jwK
o7dVQvr5Q0q0EIuIcAxbK1GOMO597GIEoSOmHE2/9zHEGik0LoVsj/kPh0p6iUYqnboy8hAaZcEy
1CqyY4xSYtDr7HOazSeRivXi87Et5h7iekemx59tfzO1x/nNTlPGdZpiuul12laEv9yCSSJLCI2v
kQYMcuLmb46acZmVL5gHnMqkZD3A0B71m7U8ZXqEcBgMIQBs+3VoW72TmJHKtTIFvNqH0VXAWJv+
88N1N9KkHcjC6GzU5jW0VVqsYRPSoVrSV+4JRBL8xc8y3262+PE1Mtaz+nnjjH3ta4ldHvrPcBAC
4C5qBv6agj170A9QYFinkiidmKHR0pdFQWDp+jVJ16hguvq/D9jsC5vnKiFpVfPIMTSkDQHnF/gG
8eh8+s26ND341e0hv9XsjrFCWEP8W0O4eNaBObuDq2ekcWcpofmHqCJWz3MGa8NmcbR74m69ctRD
eVQpoSaMuzTtFa/0IbCXVwZV6HCDUO8q7nEKx2zy7Gq5fj+/GKtdM9H68e56KRm/y3NwNZcOQclM
oDkfwiICtDuSQIN7GgQ8FuemLeh5HDbTGr8/g3VBqDvHig54a9fN7xDNe1HZIA+d9Kfmnvf2zXAs
YKz7NvPMTPUH7emIAqzsWNLl//PyvGAYgGdZDIxHsJPh3yCcXHZHS5WqRkQ91q8iZ74EhRQnn4pj
J60qw0AdWAEnFYVrfptpGjPAAVNtEmdE+/mmFZ9aBiOrKYWAMflc2l2mTOG8Yy8EwraLd3btlvpB
b9YHZpBymxm5DE2l+exzYg7NnV5flGXfAv8VpQpwTZB07dI34oH5XLKsARgDWjK7sI/u0GHGo/qv
Hv0fkwIU/x8l5ogE/Sf/G8bpXoON2boAlo4fsh/ZX92zfTeu7TSCbVuFFFDbQ2+9vSynAN6CT1fV
FhqjKnsmaWd1SqFcKD8mA8u3Kk4y98RFLvzcxRgBumJ6BCLJ8ryevg2fasliQtBQBQdbJGWDonn6
SlNbmcf0AOcub4s0kUiEbPTvHXHVXrp3XVFN2ZuyVfIgGtCLlol43+9oFdglhoyK82XM7VbVDzJb
Y2bieVqiMbkJP07bT1vhpkYaqUtT9xM7ef/wJvHawtZfVCuiZEfv4NIDdiez591w4xZXOk+4nrZ4
Hopypq8/ei3MCKz0XVzpN96soFd1/mC14eSetdsLh7pHFFc5FCnicCoQkARJpM+ocW3Uwa/lG4ht
zmWKfR2MeOflsj+nZzn+9V17I0HSJMP9c+/gZTHPiEaPNFVWhM4wOf4KPBTRlOS0O/kqGvV5ZKwg
++tKRQVxZV4ydEoeR4qBOT3l7CcZPdd6YL6M+IP5tSIXMXHfLE+DZ7tLC4x+b2Vb0cQPV4MFhyZ9
LqKgbT27QwBya7wVjIEEWrxmj/2wWvyJo/0YfhV4K3pNSr8Ybj0ho+Xl+V/tlCVf98yv/KxNf7Fd
E2fUw41rb7drr9pirjOvgGgB7HFMWF0zJoYwRUz86n5+9ToIFM0U1vo5WcNrO90cPdxi7Lnx5mP4
459nFQub+MDJ0IiMV2rJO+FDSrlrF+P7Y0E27HrR57WxVr2/73VfQIh8gNAZ1wFbuv4L6oz36cze
i4D+51faklm/M0F9CIvUsZ1TzMh662H1+RNOaDTt9iSfOHVyJiYRGsWOCNar+fxhAsOIPyIS12il
zVS65IMM/06R9Pejc1SlK+qAylAJel5nFYv+zscpBncrdSZytqujh9jqTdUloiBuci2DKlDRUokP
6EHIPeXMY1WuTTIACSST6X2eBY0KnpFowJqlqUnu+nccpnwIIyIQttDnOVFAcZe6I8JnZshAtyOk
ubmMy3cOdYFzwv+CuSU3Z4hnxMs0x+asQMV82vqy/K8b9dOtwTSyiwAn1OQ+lb5ZxUZHzn7x/M4Z
4p6b5ifNKTQzjqbxcMs4VIjHBXLm0vkPQsUXxqCdOwV3GbWF2pfk7aPTMi+MymvdDEkNE9R9hbWL
n93tjoFyxsCdPGJCmW3WVzILrUh36hQW/cwhYzPqKWI1N+ereVCyr7jDvZecbbrL1y4JzKOr8z1X
7W6s5jGxNG0rhN0vNT50g+J/I49Ew6mdT6blgFlafI4zZV7bLNwMSB7FqoNuMl4ladCt7MmoN6JS
rUM7MmEJQyF7Z9Ibi2/UDcayb+diA+rs83V9DqhgKxep8PCeMw8xg17eGYWHSmJquJuJVWrn1t2o
xsOjVXclAe5BMqhdZX2IY2BioswoNpuuf6HuYZN/qzTcRGcADmL0j7pAIZCCxsMyPBJtKtUI6KEd
QiP13csz+iQmr/Hm09gZp4hUyMdI2fSMM3CkzI+s1O3mM5F8Z+b8Jd3j1ODWpyRRTZjjHqN/tkav
StjzP6Dwhv54p7S86DtxnOB1KtXOLnL0/izML4iAlbJHDcMqMoUZ11yVtGZtjGj+z8/eNCbjSGoL
Nl+qp+zf0R6fZ5BpPceMqMtmERIFVcb66buEqxkYNRJj2ilDuYeLwOE0Gj0r9Bs8FbFF5P439Mt5
sXUnahUO1Wqr9g9z5IQpMsxQrBK64w7x3srmkd/oDEOiC23Gi/1+nemSL0uJ3Ah34w0UZCtV6kOS
Bl57QsQmeoOQ3XWZgI3YZa4Y2o8XTBAoLmlVG6+j161nJt+b4BHKrUq72TpdIDoLCSDEpKNxKtxT
cgfPmPdQbS7U7u8LViEKWYNR3LJ0Ebc4/B+3MbZHe7w3kxSpBT/U6Q4M7pDroUor+pp5gSyaUX3n
bIb6uU/ZmiHPQlcniI9JPuePnOzNwJUIoge67fVtHtDbD3MNqbZ37Jb4CYYWQyfM/LF1tZDO72p2
DBPND20RmoUD6WUnGz6wCmpyQyevwqM7RycN5h6sM+XJMLu13oUqAibgOs+kYqRxs+gXKa8cI7Ae
A68K8fz7VXmccI34Lpez6revsjNzD3kvwCJrdUREqqAbHBg+y/GPo81eitSzOn82n04FmCr2UsaC
TKPJkwwCBkV8l7ETiGg5GxKD5/fCQx6WMy5xGI7+U9hWaKMHGzYgQ9HqynnWKm+DgPaQzW3k9uu1
evh1N9Sljd6VuF5R/mbfjYWAy5sInO4dugMCmjcihKZGT4r7gFp97VqAKhhtjsp7Ssn/I9jYUn1d
CSYPfBZ7Y9twTbGQNnK8GjfO6L3YppdBALig5M5MK25ZOnbUq958DodEOJ22GztbBYbeOY5PBfq6
ZILntfd3MzvHrXi2STh+4CGalz82xLWr5jsQUmElMqEaVrJLgvTVZQLTS6DqZGXIW5Jz47kAz61Q
5iWeSO1erGqcWhYcd9CuIwHGx1WWMz44BasT87I05WpWw4Rg7HSKdH2aZIMNWgaQ+oczuhKKwii2
YCeU0n90mcM/qtEjnt4km2CvBKO7Sk4vjgHCaMNwNfSFfdfvLlVH6VmRKxzPXZ/2qJrmSM0YLLwF
ydu3hV+qsHhmQYurv67CW022favTqVYDYfvO0CX9gejc0C/kFp/dhVdKSiL0qjRMaFKJFwfIxbNW
Za23solSOcnKWoJXs9KWthHr6RckIUZbMFr0sfrE2FCLYRFNKT0tcSXC7MvA8etbFxAAvXHSIJ6a
ZHZs7ZdYA7S2mqDFS7oAZUr32IFlKIRUlTIjdOOh2t2lEv7xd66y5v7yoZamokYKDawikBtXwd0h
IkwcXpo8H8pGyETXbY9/mj1I4gR54WWWT1sVilB249zXvrEeDYAS2Ij19BgP4Lb+pqnOiFzQFqYl
B98ICEjs310j6jVFg/DTxvP+yw8IqjWcUbpPEzJW8Jt309YEv5mdDfysqJnwb8+OwnisRouaF8wQ
3hMHcpIGXMEBS9BA3x/JxAvpmTU6JurlPBI1CtpbI7Bn7UcvNUmzKAWgNNwqM0mJVLlubgOKJsLc
IAdnbOjxGZFXoOmsowcLu2cpjcq/lCBN5p//94qJ4iN5dLIBP6sZYaU/qFCRGSQwnO/4QlaKZG4x
I7TJeIgg1I2u0BsVJKNPyUT+WFRWjAq+XaCBdzVMj1MaVaagU8D5wHgqS9BkUNuIH0Ie+rGvId4Q
dtyarFeU80C7VZRvlCjWcXZJuYuhbotnqp1ysJNQHzZ55RWMjCXuSCReXoLbZw43ZVWULnsaHKC6
J98DWhJJB8eSU8/Fvc43X/oB4CfGV0PiLPqhv/a4GK9YHkNe79YtWrDgj2LWt08jYK992gCSCuK8
8dkuc+eKVS1h+r1FSzzPJdObSiY0sWdvBbKp8EijrqidyiZfusjYKFLmKKi0ccxRVFA1Zd7x/1r4
PoL4dTUXcjMgsX717AHPWIqjzMcwR4Z5zGA6gYpUaFPb+AnAb+P61JTuEpC8bLAE3uD3j2VkXw4q
kWXYXBb2zJc3wItIFUJLJlU76duGvcbd1Nc03QIfS1FJuQhMdfD04sn5bA3S16kRl8stqdlrwERi
cxOEgyX6fENJcpZKcmqcs1JYn+jqV28mN1SxiDc0CO3mFR/mOxswT0cZ3lCD7u1YwnEMH9gy4ZvK
+63pUetPvehxtCKGNMR9Xhl/SHo/eN901yrao2dRBHURHoj5ILqQU9q6nSjcGR4khFliZHuCbtCm
9wlXcbOmEimxP8gQC1Plhs9kx5GmhCxFG8N2vmP9u1Y94ICx8wMJiHR5+H2SGV2IPHPTVYRL4WwT
UEpMsXia0S7tORJC2P3s384UbZyaFaPv698NVjrxXF04A8VhMp/y/J87/JlwZu3RSZ6TwzqLytKw
Va//2WxYAWE3DY6SVprAWk7U8dUeLuaIrpcrudgU2W3dj9Vyb2YuWvAwWQxfZBBIYLRe0qfDs+vw
PylT5/gqrQ5gdE4jyTHxEGrt3MR7bzNaSxPl/zo2ahdtsCx8YIj50iPGqyPiqoHLwk6UVynbdGH+
U5ubDA6Vvm77FoKUYcNv8m3Kq8M5zMaQxcq1Iu969JqwL1DFPqiH7WjilS4IAiK/c+xNUTXC3QEH
R3Lq3v0eQAMZkKLRCK4RtLCoepnY6jjwReZdgzVdPZVrflESr/v+rZgVzFhME8ap4ZQ5x/+jxiMm
2lWc8Qn1igmw0Z9IGFEzpCqDJC2Zz3KRQXS5yy06PNAtQTWX5iirmnfyj6KZyRm0VjT5IE18eKZK
aqw6sDvFPdGrUnmXzn2FwVyNHiZ+nyJTsoXjM4YxA75KVW71Vz7C+94HwH2MrtSgX8oqybJ1dceU
lv+GJ3mxLmfQiU6WGtdDv4YLYGs1LKtfQgWyLpR9kTe5Uh41eGve0CKPaAR56RG4R85V4Lmn7aZV
EZ8EiY9L8cZqG2POfwzE0lN+UCzlP7CkHvxAR245zPt4CjeRoB7Sp1AX9ojaMG7KRzJfwkYlhWIn
ADGskmmEdByYQHXaUZzIYMIs1p9+zWPznDIdLPTx5Ifwoah+C3hRNaRW/JxCV9r6nFqTPp3/O8n2
UgH7s1Rcc3DWajadEbby2iV1CrdZiH7Evu5foLVYzcMc+uuBW8Av82uBM+q2LOJV/T7FMGT2oY57
HUj81a39+UKa7v+ZOMoybsMax0qFoxEw5UxhCP5bUMsRL+bmCwY3/uWKIoAyJ9158wfvBKGl01T+
AQJeWpTQ5cOt65i4OLx5llzFsG9K+62B7AM6wsKbNagKC1NWQ2r5DCUVpXk1vJ2BCXXFYZvzvFtL
l7gyY92usjlFITH/nvy9Ld200Z15OqPY/2YjmUahKJ8t3drrN79R9k9PJviFWHh+T9ph/VF7LCMf
wmlEIugaklpryGI8jfMNaUUM/1ijgenVVnisMYfbME/9g+7SxehfLkea3ArPs6moKYBkoVqLKgxM
FNyrgu5QfCY4aWBcQ6eWEe9cHA1E20ChuxhclMi2hFeSOzagiLuES6KW3HN4hmSI5DvCjIj3aES6
DF8k4gA9P8GxPyxNMltd8W4P9d8HYb4nLXM22+PgxIa5YAowLnSBFFbk2lVhGWkvihQi75cGGP6B
jWoUZmV5cCEFxWNJuS27AptIK6g/CbyW3GURPS4F/+/L7tw0ATbvjmQA0FLcmZ/pY0FY3gyhHac2
6hSyoH2b9P9DwaoSBK1tuz3Wzgn+NE57pNp1QFD9KADYnZMiISHPGbX+yIIbSL7Js7uHSNobF7DI
znh5W1/DH/GQsLZ/W9Q2Fr7OcsAUZnFUJyjzVvRiDGYzONbphPhBXPxbc53NZe9/uUp/dLsBQqX9
BLERX7W+QlAE0wNWuEi31a1G8RLCEC5NKkrT2hw6uB74MjaqFOW8lxRxj6nhbaMiDMEg8zDnE6Z3
sILRE/qjZMnPR4DQ0dgD4oCDobeMo5pQQq9ZcJz6slDXbAz1Lz8PjFLhL4tHftAE+NYC3y7ndbyz
lNnNGKoLzmjrn/BC5eExCnZ9WruT0rioD9upQLf33A3x36z9L1ZHZUHuiueYZaCXRL0uY2qPEsjE
WLgvAcIdOtCB72PPoE0ZRLJyXBQUgyb2Co3hpfK7Gh1mDIycgCJ0hWDPgZDcIn8ADxxt/RWkWgFd
X7gqF3J+HHr0w8Fgjj4GIDp+H9iMJVv5Pf2M5+bPD8yt9xLhwNHsPEOQWaOMFs2py8fLcnhAkfY2
dYYuHBgQ9L8DQL3adXGPIVlHYcabM9Wad3cZ8dFlYJUZqWTRUsWM7fUcmc5WwMobP9ZKyideNXI3
M/XNqQQugoJUnbm3+gCoaNyfXQSCVqmeM09zqO3wu5nNHlgVVKfL5LxwXz23dqjvZt4jkLmZW2QM
4J+XAnBU4nCeRle4bVLG/cM81R/mhF4+A/ABUgK7fQQDFoE+7qkzE2kPBf1lHhTy2AxGUWzQ3an4
nXHZUTnxCEM/C1uT9fO6dmM1/BTv0otEvSVUMeU7AD7wTGXH1wIVRKjH7VQDtOWbUkpxzrjUJ1Sv
fTLqRc2NByhFhieRBrJvT4pybEgPtaUOll82ogmMRvbE1YmP3nzX0nUrxNSah5KXx74Fhjb0jtZF
ro9q4lOARstwissYbenwHvTPF2PA3tWXGcndIYXkg94aB8TknBcOv7GywODpeR0TuZ4P0KFek3an
HQDDmkZ9M8IIA5VP2ZM0aWjYwZfrkhN/cDC7rkoOOC6pUDmvzFfR72Ic+rGTCwH43i4UTNeCNddG
z++kg05lz0YxL4Ut++y1hvG0brFNsEZ5n8geVOljSey5jRKmMApW67aaIiaqPLuqY8f14wWq0183
f1SylkjvpyUfUqFXaQPPK8PlMKcvc6mUTCzLhC2OBe6p4779qUkdLn+EO9Dub6KfADSi/3Y3fHSQ
YDix0+dV+UxgQoXYnBejRd1h45Xx7YYsdMl78xcEcrpsB5c1Sgc5WuemU80m8QXBwK1ndF6ojTZu
+EXNwlrFLXeUj0+5LwOKWERphXfzRzeZCzgdRXXeR5cOfo0FrPj7QqSBkQpbNGFTpstsWOYf3u/b
BMMhsWdZXqOWXLarhdjn7g8fh1ATSafxF5XYvTRrwkIyAM3wvK97+BsAkl91mV3FsoJY/OjAZjFJ
2m3m83qQeK+zRQqxwht1GaN2JSFW2MuTF5EovGtFMF4LhbRkU09M3eDBUE09iE8uGtyTyZBp2PkV
PbDMokBT5BjZIqyB6q2zMm+Vj3fzz13si1W2Df+JjMR7VS7HuEYaS06Dk1bsv/kEPujVl1SYWaqm
nE3cVylkP2d9UMKDeaUW+v8/tuNGPcx8ZfJZQSrPRuvYBRGog8yiOOLqhmRSHWjA4YSap0g/VI+C
ElSmKPEnCfJ7veDIuIpFsWtnajc3Aa7WNMNZbV3bwKG6MThxR5AL2lCJV77qxpdyoBJroUPzQyAh
38tvhpJ2YpOTfubiJwHDbB8NzzXBLBjSyVwdXWpvNnZPp2r2y65VKWlCXn/Stx3QWNO8XEM4VwXf
ECFUXqeRm7fn5FBGPCd/Ld8zYgaOntWLjkmwNbXZ5954hCNxhxKtUve34oSuEhEc6vNJwUUuOQjh
dtVmcj3aKho0OqD4wuHlAYOeUqcr2gulO0uuaN1yj+0fMw6NqJW/P8u6GG8nzQuP0Hix3Ma1szSv
N6YsSrIm4ykAvdXhQ4Wp9cIiDWTiUmPymsuTJ6ip021KRhlbg5ubbRqrFt8MQpun3nR6DfhcYnYj
9uO5vikkMjwMgunGW01T7H3QWfyf7lyUd69ssVGXdLdv7br2InDTdlopukfYeE3we9n173cwDHLu
ke30qFekZgR9418kjBMCdL/W3Gzwybv21i7en3wRgCEq3wAJHCJgKTOvdwj4NMQ8oDy8h79h70yv
r7fnoR50Y8JYEDPs971MFHcXEBapd1BK8/0qEECvDyfOXgBpPYMnbHhBozkn3rGPNYFi+rrc0Ifk
4HrBXSr/8PYGpsTeCTevQDOtDMtRontzZMH8R2WYvGgrNK/E6oorhBXskMJ2nZU04V8r97pAvmDM
x6T6DFGt/XmTpYLQX6iVZB3VOc/py0lTs6ct3/pm5l8fMQggajOzw8UAhk8FvlKd0s8N7KPWRrHR
9hjG5Kda0Cp3ioxy0wN5qK/cshTnu++pnsPsYMLsqlrGEN8pNnSJUcAROzW9hLyC9q8lSp0JhBfQ
HafbADFYYLTzLAtSiKKn1OxswLUY7x+e+f/sYq3Qf09O9ZdB82Mq0HrdPlV6EwdsRV1VElbZHeOU
SadwCNYdfiYf/5umAS0riIpdYswnpGjJRCjOyjKrcRvvdays0fb9lmeWJ+eUfJbENtL31rbqwHVp
5PkGrKvwcAdTy89UZ29ZRzwxGobyNkVFHgDq2JPa5NKDsqp3mlvVwozLvW4uaq47tekcp1tnID83
wShS0+v14jKxHCyhmiwkQ6iqmBQeRZ/lnSnB/whb1wQiXb17jA6ILVNh7GCoWifZX+LxcK0U4hg3
VnsHjEGRJwamBrGEzlc2E/LfQOISJcfjMKC7Q0G8BBwBikgZa8sK2+cF58pdMCIx3hZX+ZyZKKd/
mCP7O5mL1t2roCmXkLCHM2m0s0oWDsByV7+w+g/FOe3gtdmzYbsJjjZqfMw2fUS2KPCdow4GES/B
4IpEcZqZzAarm9gKWLNK7DZiCfhzCmBku5LJdfJejD2hwxTyAxX6zoSnGyQWU2m8cK3ePyElfeZf
yP34q/N0NEhqj34Wf7J/msuxF6+R/czipgHzDpnFZ2I3GC0pP2HQLDFn8JC4GgwByhTtbrmUxqHS
IArm96rPWalLCCoHzesCpX0rTKyU0f2L0t9cUZ3oY7A4gQXpRzagYXc2ODJ3TBQvtUW20cHFjiHA
K5dOsk8V9VWXFkdtXNNUEIqaXe/tulL2yWjjokzG4aA1wXoXv/RLisxhUZD3HK0Az1xZ7Wm0oIk6
6HRg047SflkOv5Ga2+x55KzTfGp+8D+tEoW9pSsyb5Z1ZZ0yOO43ng9LewE2opbFwv07JIefIX5T
7A77ocMwTZfUyEzz4qk/g63pqF5aW6SHYEBvJIXuo2TiulA9QYOGkZSIDs0I4mb0e1ILvdEUYtXD
al3HeoydtE4RAunmwKYCQ8Xues/MsJiohVfxlZ5xUONNUlTQVoZA/YoTJaH+ZWu3mGyItoKrwJsN
yxq+MwjYvC0FBDdeWtn1Banp3hKoKlJ5B9MQ06XdPk4hSPCeycI7asQnR/UHR3S4tvCX/mEUDd4q
w23V1UdjVlEMlxDW8rvRpVlP1yOT41ozzt7FHhcVfHfSBoZfH6V53l4mGknhKzCD3uP4Efftt8m3
n0IbzWBNFpk0fFuZAFJlmC6nUHePB/T7K2k+/JLxlhSd1CRLRYQDMygkxLXP39nKU8WhNPlqTWAc
i7JL1bGXUbut6OPgp3vPRgcpVYX5Fxq0X52UcQWgoOTgtCtU0O28Xqhe0iaJn8i410cIyEsZsr1j
GDmxHN5ve4lUGbSmt8X/BVIlM5Px9BZNRnJtZUQjpCoOV/kx2lhOJCYqrCqH4N3zK1i3Bf+9pHAn
83TTzqWzEsn0MB4qy1t1oxwaAZ2n5CijL0i9cycbM4NM0WBXwc4RtoO1MMuBPSX5Sh6Lq7UpdsSG
oRLorFBQAPPOQp42F7m82ImD0HO8PUBhw2p+C8AFdenpmoh2MthEn+GmJvsd/A9a29M267gVmY2r
MGbSzlOwbBpmjzKbUYIdERn/FpxbtExlwXE8PZfY0xJJuS0VgleRAyo0U+ItN1s1fiSqoWv2mIup
H/TUexmo1foqXBWYjLHNyo1TzDiB4iboVI4n79o8ze8qYL1WJrdQTU+jp4IkB9/xteRs2vBIf1+u
r2Vne1Sfgp8uHIAHK8L+wqytEusPQOH3ze/NEU9f59n0zUwrmVvlq5e7hvW4NxeTnS10lhBy+B7T
DzvsQfYXmZsQdIhxlApvlpLvhh7XxXoJg4+PtniV0k+5mLV9kRXw00AqvTZsuNNbQIQ98HCLOGL/
/Hums2mRnu5IOlZtq9PwgCOzW0Q0HpldxD2xEFV5sH+4/DSR3rggql0EY5buiRTkTIiM28jTMl9I
YPC9fALZ4+J6tEZRAqrOvlXxlRMa8mHciladRsY3k+213tB7wERCi72rxW+QrzdbCHzLr431gWpB
gFY42EitRKIqthpqLrpNMUkMlV0Gbf6ivWNDKh44S2GB59DmYU25EpKfzs+7GIi7wrGfm0OEBtRd
zKWSvla+6vhfaPhqy8hzfmhHQL8b0JngGvQGkjyLONMYHKeHP6LOfAs5w2LLkffW1qqCvgUYGyXl
Q7ZMjYKNaZ4eXAbBV7UR2Vbc6rGXRYLtfcG11FpfJaaFULaLlAu6pGYnx3jQEF0l1oGaBfZ/uxZI
3yn6XzeQbLC/XQcQszr2HlxrDbxm53i+UpHo2SnH+6sl1mSSDtLF1QP0yghMRaWtT2Ari7/P93pO
JHO5CY7P9iZHtHKnh7g4U/qNk+Pv3kTYOG4Fxjf+caJ7vdaB804xsXonCq9btuE6orS1FTr2ebWK
pYEjjMjkysCvapolPNv3BwDCTx2NdjuXJsvc3+TfkNH5QEDYqf5poOV/46y4nry6NepX64/p91Ji
A6rzlWTiw4TCSMfyV+JSxkaNsc1kWDzSNvcKWConQVmzu3l61/u8ue7RyRf9RPQ4wrt3dWKY1mJN
6T3edAwSpOmLmsjBoDdnZ5W4+W05d6LxDpzOTAyJa/BXSRyh1cr6wAJZobnVUIsQ/whlaK0+4S/E
4y0iSdkEZZTggAgRky29Q3NXobUTzaFlTLA3GkErLQeGcL1PB6i+aAkayYZtFTiiLWVguBIXwWUK
b8NzPbYBTR8vhtLs9Lnl/HCWlf6qOsyVFrXyKBstAusQJeF2PxpqqzP19VANHDyX0sMsi7C4Mc3P
baCKyBdErg8ekq5rxynnJCfyUAqx4oeacxEAQfyDhpkBOEKQMf4KWaFaKKyQWAUG6ROpCmGFlCMj
YGG3szV4oo2NSrWn+ZbmOk6MkA0/5Ab+FBdELUnSOGh1HfBvvTSnHBA/j65p4Z9W7UWUPXIERk+K
tSjkcuslF9O+FTv/+2e8EMiTAsa6LTgoL73+oKlEQ5d5Zho0g7rc4sXRV2LLCjVdhVJovalNwayX
H5yoSHVaoQq+VHoLCi0UHGs4Xuq3zglF/bctl+aZEZn4g9NQOv/TEjPljMdpvi/l3vlJAXSfH4r2
19o4M7gpEAxXAKkJtfpVtAdlHHqcrMPfy9JRvf4Xk3xu4Mjpk+0C4PQ0PC5ELSvE6jOeVGu9qa8O
lLuPqdepg0dJ/hWd6Osey6dyldVbY7Jrr+YnqxZzKVDqI7svhi5LoEU8nb2ziMNYjkFn8SgMGiAF
fCUu9I7ZPSn/Otn/5ijznYN8I+mgnnJx90aH27kFaCG1KQJIfYMxr2EmXzRkbKqRXUNiFBdShfH3
7MxBqh7q045wUNO0oAd2WUgRAal1xyvsTHfucheSc3/x0X21ldr90REDci10JOfn9cFSJuCF6Bzw
lTj8bODFbSupIZ3U1PM+4Zt8GLtrhoTsJQw2+K52dYS1J7PRc38C7KYYhp8eBlObfHuvG/vNLrGo
vy6oVKy8SaIUhqpDJX96zgHAFxFcm66BiyW6v77I39ZJ84IcjsevYqVkK7Jnlyi+o6C0tayuUTG5
ZuwDb1HRHKQihkI01nq9phD3L/039SF/51dKArZLNK5FdX+bZByLS8N3acwuKP+29E795X4w+Mmm
vgWPbRLv9zyIAfiEK4X/7qcKoQWGtm3DFaT5iCQamF6/L8Kshyf/3wjYjuelBVONfrayQTb/JYVu
u6Su5I/bFhAxvcicGSQnON6tPhh5I7fOQOyTwUlKGqSHZkPLuYcvx+1BKWZWN9IUuVrtmM9pkcTt
PsgSV4EyTwsBJvp+9GjZNKDil6J+LWhe+adA3gpU3oQt3WamQX0pDB2P4xfb7TcWQrHDOtM9qOe1
CsmAvFlG9th1aSDixncwsEqh7um9xqV+kwC3eSJ/x2dZ2JkHD/4cWkBiJGigKjk3+ql4OkOvRk2a
PLTgPi47O8URm1khbwsMiazHJR3M6wW+sT4Ft7Vl8RAsN8pZJ09Kye3CgmZyeyxMZ4ajQXk9kUGw
fm3lsLLnUqhzGRE/9I4YZ968Fvii0sN0vvJE6B66b8/DbpXtTw5a1zEboSIXL70qVyGiDPkHlnT7
ftUXravPwf+DBrohusK0waYBX1QsB0hT6eJCuWVvhcrAl3V4NLSzMFFUT0XhltP3mV7uSIb6/X7Z
UiX+0igz/KpzqiZjgPCewMpH/LTL32rAbBiNlWuQtYhc+XvX+mJOrAY/Pqz1UPuuvUg/Brr3yCSM
DqAf4HhdHExHkoSqT3Q1hSgA0TRJkwkf6Z+dWfIiHK4lTozyTVeEqAnNXjklNnx5a1nY1V/4EcWT
RCuZY4fyXyl63dOg9Y5mtC6KWziD580ApXbVDUcPZc6Y+t0UHn/dE8qHXHAlpb8PS9isEBA+FAGa
HXeaLCsDpM1OqY8CRBgxszuZGlOv4OITfhGEt+srOgbI1LvSW8Nd1Vg/I2MH3vk5H7tkxR3e3s+W
ldHEeU08sA71s2vczLH9uFjuL8+qGtmjBsGjhBpDnVDZbZitxsIBCCmlrO1lYcaRR7x4WQX1qRei
WuwPQ3daobdcVlfLKK2fYx/w08N72HxSHbzX+elcEqNwLvihIXN3Pj11M5F0y8Tk9DGLXXI+j9NA
YoKlQs2auZ0fY9QSE937w8Ljk3laF/URS+4+0zhTdj9WQ+0pU4PT8qzZrbguDp6hVjhEbfnPlkqm
bWY5DNr8UBHt7tclmZ6+/jglzMPnJIP0RWrQeEiJ1asSwnPsk+1xDzVJO4XCnFZNRsXSVp+MeDTN
FxMerT7D7fZrkZAsf6ji2mgFQdt3gAnNainUl8cuIX+Wc2NKVeOyBSoiqCEJPlI/2jEpQEwKIERT
F1ZCPlzyr6Wt0Lq/NNCEti/CLW4T4ppoK8ybJ8W7m673KV3xSjE46hTMB5H+H8362oy9L1ohsysr
HLnYqy+7V8Je3U3ZKijGBoRs4dn1RXj5RJ8m2XDg1qYCWJgRbl9wSuEQptTUjGkbW3AWUD4ZAisi
A3JznzFYIpl/ce4E7Mm0dhjinGxv3+Fc68GpjquVHrOVlP3NQNAcm55HYf/1DRtyemrZ+Xml7e04
Y6Jy2l0btGjfuX5nryLGDPF73cRr+bvaHI2gXAxw7i9WBqxm3ZzTBPzU9r0S/+yO8jdZZEhj8FDz
Vo4o6ZQ+0E2ilEisXq7QAYGJcpQJf8iwi20z9ioTWU3LPnxEnlMiWslb+6ABvvIPUCiuX8YpBJKF
kJBQsymWxgHG/zv62WADq362k+/NnkWq9+5q3FhMKNGhqeyLSg++tXMVKbTbDa6FdSjQhhjjg3xW
AI/j654s1SYmwXBmpyQ6fembCx/4/asqzRnQ1ITmxNzu0nijpyUSFoe2us1u01NhsQOSohNo+s5a
5iZmFXVwNXkhpcMYzDV0zfMLpYBzUehwg/7088xvsk6x+mXeXt9MM653OPdF8/maglbwrVY5fzN1
wIcB2ZM1Vsp1i1t/qcb8HFB8/KwwCumRAQgpozT3iqJJ6uRnAYO9WZZ7Ambv5GlSFgLrRsGRKsfq
EiaYo/RRxRV8VIuifYUMWylW27jVjb6NTdS7ZXmNDEVzVGR7szzI1h4OgGrND32oBfB9WU5o8L9Y
ExANBYnnD9/aI4DQK398rXyhr32fhjDYFneUkUUQa9INaFiJ4kNX72j/UMax2/ajZYKnqr+pXupS
vJet4byotyRu5gGfDZYwywWyoPVr9BkldY1TDlZsfZqAviV8CZ8FfknF26dS3C6rTlcNTGz34IXE
m6Ka2Wyvuer9OTcGBp+ciiHQyhxFSzaDmfpoDjsGr5BS9pykfLoBjBd5y3Oy1IfFfg/or8TEHwiW
Df7SAXCg4YBmhfefZ7fGSBY7WqkhDsDMPLl4k+MwnrJKGk66LrDpbLJAoGg0fLtjRpDZgVR/Cahh
F7JOuULv2C5QPDLpzfMwM6wIQLM0bvH3hOge1nzrWSg0OZ/TMNZICn9sAMJynYSZ1HFz/sW34uU0
wixd9LZarjmg/hjMrxw33c1E/J/W5HjBOIG+YWRPjEaAohIMLX+EUja+Wz1dqlWHFBxUs0GGTvUo
Br9FF65MD+63fidUnAciFDIlXiKuNjBeTLiuxbIgFV4bznuVpEM2NQeTIX3nACWV0I+wf78rXGur
KgXXSBJyay7iPr68KpKf2S7YLw1vZ46SpTRhhll6OYVpeL9SF8X6mknHqGlYkxrvsPLCww9jLhgj
662qa7ZSH4b3UQ5n+pbADl9fn/aazlJdWLz+YbHJWAXcsKtydEgT1Ry4+FvMa08OCpB1o/G6vOlx
9lYdIHr0SKTgR3yyIbjuf4CZD4lWb8U9XiZ+Y2/fZaUyWVzaZW8tLkZbHf89daLDKmmtEIEsldFi
foocCUQ2/095h4hpoQepjPEuN/JIWPGNqwlkdqCixkMXNwFwC/DKZbSoL3RqlWKHWbq0rCHTalTy
eo74zMuUmHGFt135gEWJXeXyZ88kVLOSuudx25YUE5fL2EJxgUet8aEWfxIrQYRqpipaFDm+t6tg
UPoyhwASp2qMy8OhOctriUYjqNIANqLQ2WY9Np3Qw7+dhipOZsDhYx1oqiCPvs2HwqeGbnh4IDY1
rd7IlzzkPWHwr/ARAZBplvfvUvaZvqg3RTt5iFdVYspmlvwsJvN6zrsDL6fuK4MU7o8PSZcjeqnk
hcCIU+els2Y1EPXsEn+cX0kw89aWVNro6QGL0WWX79vKkltiEuPNISYk0hoxr3+FoJlbjSi32feV
DvQf/FezilTUYqY5rrjwN47QHJrV5s91f3I5tV/1IYCNKJYvViuZo0Jx4W1tSfSjben//rMJeIAr
jxi6gcqvCKTkD8OzrXGoAJ0QCvEc5nGgVF3TNZmkQfJREtKZ3PILJLVOiAyRN1hvuoujvBPIgtZ9
5pdOA/n/dGw5i1v7kHcBPsv2ytNavk7kC86VYhYeQKmNitiKtQKdqRjH+Zi9YlCXzmspXoD815DH
Sf57IBgqDiTe9XRtPHQqBIhdhu6Al1HEaqyAo4UKVrjsvDRb+v5T8p5qY+K8PwdTCv+iseG9TWCG
vbUgeQFyONj2dQTKzScHMZR9QnAQfVWEM9Ha0RxUMtOz7xhc3gBhkU2WP0dd7wkfA76SCIlNAWax
HHTB/YKQB50FPh4AAjbMq+a4DUr6rrGxopPdVeFSjix+4ICtjQN3TxbSQ+DTNIbQiKBwd/2jbgjs
MVfkXYUihP4Jw3d8KnT2mOT1Ss4jhCuEQqUl8ObURaXfsfHMeckQIWjnblox8CATcX3vVbVukCEp
xXufNmOHo85xYozk6bOOqn2SAbOSWifoel2mSWt95ELSutaaniy86BSjblTTRQ9gVM1q/x0xosvN
Y4rQELPzdXOprvr5g+YvS07Ezmsfme8KSsovJ+PHpJgKSFekhABk4Zt9Dbf2JTlB4QWStndlz9RM
NfG1WFqmjrFdhcI+joLQ3Z8bR/qxk/OfvxfK/WA+bCj+iJL2Uu0G7P/05XEGyjzRTDcsL1IwQaqA
TMBcGuAhozPwVqOHpNyaiQUfh7f+JfTBtvnWzAv+B6qXTx6FsWoOuR9iGRuHQZem7jfb7QEStIcL
ta/LkqkKx+tuKXd3Jo+OdfKHBFDeY58jcRqwK326eiGDalbDh/aR7YKBZLhGY2sj5e/hefHFIcDn
8WMTpNg5q9P/KC+nsG71b6qrAnAuaMkcIqgA44o1BxT3c77COQkLrhWS8KN3QbaQxXFkE2d2FPB6
suw8tIlCCpQ+z/4GCgfF7spMBkmiwz4nIOuE4v7rJxvBZj/Dqf4EI0S3Rfp/03mrd8rbcEOl4Z+G
VLmJhanaJkqoR3m6NjnRATkmD1DV8CMeJ5B3huejNSpMlQ0JAk6ATq9kDeHOAL99QmZ+0n18Pfj0
lS7/WSROsBj6njwWOl5A1Rc3TfExk36zIAqqDL6Odvs59GQEGEygqyHb2Bw2VfnmBhnhEY0mwjdN
DrH+oKHVscqRN7cjcIU920ZQhJJLdcYKKGn1KDLEdlCTYpaegGxzzt2qTvlnFtvNwr0MP+AWhh20
UZh9hLCryIhE8hwwZBddsPEpdFdAE//IgtdOwtYKQ9voRpJHlnVi+gj4Oia/QeP6lHkqtbbs5ZXO
8XEQrEgSDK7FqHt9XvMT1aMhBsqN15sRI7fAPjEzcwhBFS+W7zm+DVz9CacrO7anaBs72l2QgycD
2BuS6L+IOv0xiUpIDbAbIWlGnTSc9n+HJ3XOzYS2IKTnD1xDbLI43o6eKqTChJG5w9bbyS9qarG3
kdVA9s6hLJd3wcxs4KD1Ci9Cz/h1X2oHYpWVOnYDM/m50b+697p0P30Q2lolGNuig2mXNW3PsCdH
/DXQ3MuKo4nOOsbOLiEdx0nVR+y5jGEa7f0YLwol7KslcIjyCFDB/93HQT6AmmQf1OV9+73kPxaq
pdU0BJO0KaAVOMoqfqBRq4GT7eDr5wkhx8+lNj69dlqvOJCfiwTvdeJrYyzNK/G3fuhTExlBxPG2
2uCoEb8Vcyv3//sSsRsTGRqp4DuXJdpsLEIokiEI3oG9Ui4j200tH2XxD06Pm+SWG+9b2j4ZOu/7
x2ECCA7ybE17o/r/IFYdEgeI0A4lKUOJlhe4YXglYObw6XIXnWoZb1USPzzF8DFgTgbje1pfr76W
+gdlsv132Bsha8jvTyzmiqu0E0L3CjYH/3G423HV+QsQiONksD/Rn4PN6jgfu5lLjDvDJZM9pfxb
QFeCdQOa5eR0yYfSUBwp7CWe9sHHkROZAnihUPzNoLJWU2xt4F95GEK5UNqYDk0sY0a9G1LUJaTs
VSXbwjLr4SU5O8pQbCMCJ/0l+sIYdN7P7xw4pcdQ3hX++BBHEdO3KMTNQzjqpGWPZqEWQeHZD4OB
gpXbcsYaYwMREJDyYQkd0/6Ct2jJWVW7aHqGjWT13YRCg7SnsJUmEaqr9W+kFdiOL0JsIGXKarZo
I28eCH9aEVtPeDnf2zeabxfTKNkI/t7e2oxAkdwOG64VhL1kCKWtSaElH6L4yqOV9GEcD4i7U+uL
gHj3f18FElkNg/nxc4bMyouerKogbENAtHLxKSiGCfGK1YV14cZKplxdVTuU93UaQGnb7wzrxFU3
E1RzqaWmuyBVrF4CJTfEXINwinVdRHfYtGYtxO2Y07TANqz8vKWWIb1iFgdEQV2bOeJWEUk4bOFx
ZIDTw0G8jMM3ogLUTcycXfi2fCLECEbqP/TmAAPt6EW4urav9v3eg6pfYmOdFLao4Bc4gQot80Em
KMalzrdoLSK1oVJzQpjvZWLQWURK/imj7pJ2rEG0WFec+1huoK/UkizNrebL2r+srjjnbnwihNS0
W480S37mqwCybuX3q13P1uhdsE/1RO1aYXdE2a/KXnbbptnx9W4TmXVq+SegNhOC4BdTDTz212Fv
HltHANIdjVAxqe3SR7QFtQOzyMoq06u+0ggnrNqsj80MSEW2PDLt2zsLA9v636G35tafMM1zWw1K
v8FNJ73eC4zaG2yiQXmqTCa4nmoys6h2FWMS+AB6BW31Bh+bU2c7rntrnve/Vsgk0MYC9V4l3N4o
YF4Qi7+Ot6FWGCQdF7sNbB6b8hQyPGEnaRTnTCMCQsBrutQ/brxUpoBtf6Ax13ptc6SsZurz4/ld
PbJJu/BQ3CQqNeQ0QzRX0bxrjnuljYpvKi4s9GHHwZgsvKEhih1+iprArIyWTNcbp/SiXAP4h4VZ
3yxhelwPQn47zmFpGgj4yYBcbkpCHBqzIyhUh30uMC5RTHZyZ7JA9p2LhMTTRaXwkkFSoXynATy5
dng8goqjvoyT4SgdDkgNWcErkoaX04cY823WKn1Emof5P3zfX4vYSut8ba1YVM2METFmLuhC5crh
AMESwDcQQToZVTbv1LO7MbjcLOhtH2nZBlkZCYAyxMN44uvtw2jSAyOInmL1afWLZLBA2tsIm51N
HKGCww84yW+28Du6IgucTM1cR2pW4ltczmJbPiIw1afL+EPDUIA7/JiNmTpSm/ocwVI6wq1n+ucI
9bdp4n2+zboVFX04fHKVdFShsP6LJWqvzHMLx0+3WOmeE99VH5k5AFrxVLP7R/o0woFhH61bx4Gf
8b27wcUkUBqZxTKJNqruQl2e24C/KR1fo95u9XJCByC1PQccDqIEjQ+9O8uAPznmxZr9e8eXC90k
Db7hZwnFATakPrLeiaRk+LKoNBc8NGid/aTxzwtHt+cs/uhmdlvaMuWArRHS0EIpgR1de8yidK81
4nAufJGjbgvz9gUTEuSiDdEm1VrxDCqwNYVsL/gVM6cuwiqQ8EGPeYmsZjLfdH9FbA1AC/F4HliY
UM2Hk5Xv+clbLYTH/ktuYW3KKdbTXQFivet/ZXFW+4Ua/6tKDHhjtrkMvDsiaOqU3Fm5fwMMVYxS
spL0t2X/SVvH4RXOEhxvPWRjqSelA0gwPWXoIjZEgHR7RQraS1tjeD2ime32N/wYqWCv5YAdGIGV
QCz5D7ne7Ur/nzdVnNHFj7Sb/qwdg08Xi5M4tMWAAivE3r0VKk4zd1gRDqbC+MOz06tueoincJf2
qE78hNIDMMKt0cfsJA3PMwYZf03qpxuYzVOxyI4RLiYSIJLnSSARhQqF8sekUPNSXvPEq6qIq+bn
jza4P6+ZbDTAFk3RVEOs72MxQzduM0h68ZZeVEeJ6AFYigy/wODSEVy88lmGlbYKq4ezdQRej26U
vNczNahq/5eFLZsYAfje9vLPMjAbw94mTcnaAWAJcZ36pO8slAzqpalP+x+cuqB2SH6HVBQh+ujK
MmPW8ai5Rvaby+nTbp2zMhcWCa//jYxrpJPN+liCyb7Bj7167wHUWOJH2UnAi+SnCMC94WnAcUFI
VpPCGibn8EhQOY8s+WGHwhRrjm4kFikOJZYP0DR7Bht/WQuVeHKO+wWQfQy4KnQzq7cTH1+7zGLw
NPxFCVB6LcOmRlvT3KXYP78OJAOLeSZHIuwmviwbu7g9xU808kUf4KlvqjjbxarjCz5a48Pp/h8J
kJ//bADgHXrkm6kmg5ovsgDr+65AQylVa0m94SxE6Q62ZKMhn5Lg8o6PrPLABUFs2fuF2XSS7lbw
YNQ/UiYz//6xlZixilAX9n/I2hN2Bt3yVQvpBuTDEPyacwq/WmaR4ya8ExSyrUZxOy+Qw3kSCVFd
zC3WSqSRr0XS2kkrqkSEEp1Ysr6giiTcFAOzBTEaVEm4Pfqtu2a0gTWu4eyh41xurjn+oprkuXue
0G50670orbKRo7ovup85GhP42SdkZP4Fkai74myWNATJArbCIzijJ8TshpHu68Hqe5JAf0sT5pIw
33+lOTSpQs2RpdBnUMkxnvi6ZpLd7Jkmuoeho6zWYm9iKJyFdyLr/BuEgGr7BeaRKoXFPUQy2XBy
sJmBkz3MI5nK1TeP683SWaqdJCTHeMH4pmVBr0LPpv0LaE1yp13WBwEpNUE6lDqqvadRr7Q4zXHh
uVkvPqHKSSLB4JrcZQvfck/fXcdFwUgefoXz+ROQephdf/3WBazBx5d0lZkW+fwjg7YVGPmokhv6
4aGXQgZVmWNXBGlJnMbFkKoMiwXvPzIEj34M8HO/0f3a5KT5LcenRt0tklmzDSf7Z5yqFlHhdBpV
DlUWhAGHizx+pbJ08gD4jw+NntaFqmi/HyS/ssDT6UVP97OgetQfLy813ejy/7KicaEQz7L2HVgQ
XzwqTzsjFsqbCs592qU/fNyTjoeXh/6E90SVq8yrU4yDf1MKRyKAowHlX3FkAvIx8Jzn3Afc6NpG
wING+PDQIi0W9N6lzSRajroeDG2OlxmX/onwdLx4Dae097D40Pd5zIZZ3fE27i4kNCdyQh5WjPkH
bS375B9jK6GzjZhKRR5wLbbyCjf5y4oeEcGq9+CxZowxa2JlYQF4TS06ia6asHBXmMcG1vFV/jcY
bP15QS03IXdOHg/rWky5U1QVAQAUVFwiDWxy3dWIbL+aLoKPXmikpehyCpIVdQXmTFQXUSPwz1A9
vqW75QlyPs5v5RFdNDIPYeZ2aw856ta3rF12SO1u3yvTvudXzkB9GL8TW+Qho982gWKDybGgjcv9
tA3gvqiP700yoi1yhPt2X2IG7/irrk6GYG/Lw+6uT4sU/CPLZvDFsVguf0Adfytgw4YescvcPOFq
QnCjOdaQdZrbCu4RrcgPZzF7O9pP64oz3SSzs32kutm1iZ0fBsPBXYp6Hc8y1+VVANWH0Hz9p2V/
qNnbMPYFw+4mMqAsUWHlgYvtjOWHXLXZY8+4gN+OirlyEEXo7KCdpAFmsZv/+HKyynTcTWTNEWez
Zrt93CxrDORCae2iRA6vXNITzrPHumAG8rsw0w/EqxLtu6VLghqzbleDQNbbzEIAjCotu1//9apq
Mtdigrsi9HtbUb5aln26PadGp9oAKoA/hm8ckZ51P9e7LPABL222i62fWDCWYpNzPxxCX8aszv+h
pQY7DYE1uOrNZQsEI4OoAHxp9TsbKshWHrSCvAViq3/eO34f4ho9R+vSGrDUUYICPTmFKVEj2ttP
8QW1+EF98oFUWYU1UZ5hsf8Wk635UtZWH+RZnwyZOFz8q3jaHkydf2I9QoB8QXNSVKcFe/JhdOIi
9uqUQ3z5po+n9bRRGXQeXNCSyu+GUn3MaRcIz20Hjs8VR3s0b1CZ2aM3oVD6AFX8jeB9w1/HRyOH
lDpP56B+RdgwMKXnQifOK0dmpBK8j32lthRi7TZC/ZDn0p5RCZCFQ+ekunP2BjTdT7nzFAr38s8u
90Ufls2z/94yOyd8NIJkvmN5FPZF9asi0ottLf6d4X1TxDMfOEPVb0XLP2w9i91VBkkhwNmzZ0uQ
aPY4ewBG3Rldx3FAJcqa4E7nmtyfX0YO8vsAkO4nz8zFE2jGND+qX9bYvR/jJH9sIjEYwl7vobi4
m86NkjVFXfvjHHhvfN3p8TyEDlUJbTVN8CwL3myxKdeDUVk+4D03p8nB3zZDRjHD5JBsCKgRi4ss
jwZBeRgVFHI6Fky6Ol3eNAX3IquLyVbPeljrP3tHpl75cK8mFjpa/BKzktl1YadM8D8Ayt0+swbW
B6g5BCyyTRRMQ6TkC+u3oQfughYvef4TbwQ5ZWobMlTZVfgycddmpx42ka11Q838C3MOgoptJWs6
kWY6yxCugEK9+jzNliH2doZJx2moaCOwSczjMCEvHhq7TqRKpBQ6Dmj5KcZzbhwFPx2jsXYK4M6v
jjvW2wwi7e7fT9MTL+rJx2v3G6NTTIFuZh3/oUrI5t5zuURfUWKX32chDlLrZIjn2QzmGTrxwxBj
iVF3gqsw3Z3mXOGPEJViv7tAKiZe3v3cDYt6HVLvMlucaLtETIC2trYdEEyhPGpznJw2MxZoMhtY
QluRepJcJRVoVHtKNEH00DzATUNtqfohORq2eYjvpVWmDazUeoI5RpB7UXBYB1C5aX9+5sPAXM/E
JVH6y7whwp546TzUhMQuS7yi9W5TUl9GHdhNFn5mGCCfyzKyKwQvfMcPm8dmkgZjJ9jbres/d6RY
2k2FPzDyglbUFqX+6qWYE1cA6croMY980Mw/h8gR6eUjZGTY1bidGPLaGHded2KJngaido5IasDn
9G5ormDXkehQxRJ3gEAbLTnScwKET+wi9ktW2HtDC3hGVdDSgIFlYQeiwTNa5BWj5wqAcNh7WGX+
Z5NjmIkP9ZG3ck2IvrJ/c1CfM6lmKX19u2mNr4AdaQ2k35vohdQh1kLDBDp1rJ1eFyMScPk12N0n
oKY+Jo+fS93ydM5AZMxugp/VLLkcuz1tdnh43SKt+SywvrTzKRnJHj9k3eyON6cSps/qnQp210+a
IL8EfWwKKqgbtYp3SIWPLOdL3VjtgSRVXnJkkZozyyZXi/6V9P3+edT+8kyfGqY33OKpxeyjq+GS
T2PYXCA0V3qjtHNI0kzF6KORyzzKx4zPHbB+9nYfaIxAZqRxTPbtfWSGjI8Ht099FItrvbSW75Ux
VBqQhDTJzIP3OF1pdpcGmNIRTaVZ0yNCNcVV5lsaO5dpoS2zszU+PL5pEWArCdWNBiUKNRFBbNSk
LIXBkgJAkA2SUJPKhlenkuODSzKQTMIpBsYcDs0HdY+VdwstRY4V0F7EujDQqk+jA/JnZ1NjNfzW
VKj52BP1O/ifD9TsGhe9dBsukuklquzdA7d8KjiGhga85GlYBHZ7GMWmM48ICMoBgbfW8Sj+Zq+v
8Vno3yMMc1zfu6RDjnWT5eoK+066Gd8ZBLaEDPyuY3vYNLnOQN57wu/14xoU0F2NRGcJDeA9Wns1
18UsKUeXzunjghEpUMo8p1ylgkRvZiqTzRV29Nf2e1788wWM2VBVYJh/ZAJHM5hZpiPVOnXuMXw3
7hcEecNSZoJDt4BpHbdGIq+fW5LLC7fXn+8rxF2o5EJAixv54Pgyz7V0bZ2V78cSaACZDen2nx7A
H/a1xgl1Ucu9U43KW6hfipSr1oQse51L+tmFr0aYsH28ALFVnLe7OkHClrQKY2lDEyHCHD+CCJqa
xlyr6sapNaHavbkbFebSuItGUOGgjCdyGuj2OWbi1WgaVhHcY3IQ8Oi0m5M8ixtgk9EQUMabCDAo
cpqqpkVWzpDk2JaCgokp5wMkqgvPonyc1l0zR6jIxUX6gUjVjIqsAGhgeC7ijQIHBRUHMp2TNtaA
RFUo1PgmsvWY5DY/36vl8/eC9T/EawJ5yhCMeew2tbZj6yIwelZJmp0BrTOtSIRY7CPW9O5zeEmL
0zDGXl2xDwiNS7w95e5YOkJ9UMLZ0J5C/EsXxJa1GbrJsoBkqgXrQVrMfwdsYHy7JI0UsfFFX7Xe
AOhlEYmeDI1fk7inVihjyEpfBn5oiJ5rHvOdczHWwBWw4cTEwb9CZlwkeWH6NLJiTLIGg9rKL0S1
TJhAUBLQAPzNgKUrdCHSNwiXH0dJlukUo68++vWa44uAIheR0SoO1mD6arm9hidByFh4EZyRyTrV
8B+Ut5hRWjjrVovWykvCKYy/FnLDdBaIv2QLOOUL5INKyRxpDzuT0eyVmj+XXcfrdtvjns6gFit6
YmRDYGk5dMuBMhAg6OhU4AHOXii19QYxtTbDY53yePhu1s+yR+2oAUhmjIgymBz/77mhKM6e1QGW
OZPPIvoip3AvmI36mQJFiPnmakOM8BZWUqjRC6pEQm2FZFnd4WiVcJBJKV1tj+KfCFdG9cr3qqCA
by0seo5KeX7XNQsKFJ4S64uRB+n/4ne+D0T/TvhWJoc+eOMCnHCLKAk0GDpRs3YS7PHrV4FTob9n
oV7tO0asvXyv5Bz055tYax4y7GNGdct9c8/l+1Y8mes87JgijvqKGhyq3ryGH24pzhtUjtGSEezd
DAcs85cRo7X04uOEDuR06yuhKS2HNS+6FSaqUvgShz74mu1yultP87Kgenn8GTW5mZ+pW+UuT1kb
gMjw2NADlQElZBXfaYfmFOaJBRPQ9iQvfCHoO4LC/L3GSp+Pn6YO4kP5Z0vIu8qByvcwIcRBBBh8
H8G9okZBqeNGcld+esjwZ8helix6Ok0fJ/Hd5p3QrCqQUGHJfhwOOW8Myhf0RKn+6ivNiNH3H01k
j6nV2TuJcQ+lbt1h5EPG9Ec+rqvGiAggGpcXJkFk5XCjOuPIHRXRiYNKReJh+MlW4OZSXkU1gGAj
keJBQPl+ghEcxFLB2+r4qHAC/aPeziRov/FazI7W7U5/0jsiI6OLzbKT8fisG1eoW9XAdXIuzTFM
VXHlOzNmTj7WflEu2XAMdOkfHAjPAs+yXZLuZ94ISZa9v1bn8vXGJyqSKzlcp/UO2I5rkVxTaK6+
GBO8DzCSmVcqFPjupTXitaxPfEGy2cMCxkafFM+j88kcXcSEQTLgQB7hc69DRzpZv5mYsRjBiUTw
Wrq2ZeXMs6y2RIRwb5VtTo32fXqLU1vzhGhSE8MlVv3BuhMk482d1Q91COPTii8oGJDngRtI0Yso
qPQ1AMd5QF99sDNjRQt3tX6/auZ8EX7p+qcSLqQYSnUwUl7Sdkt5lbIf53Cdc+bM8cSm72ii5wOU
MUC0xpaIo6zfdMVCCbCXFATGpDNx2/0P1KVsRvZVs/a9nSyCiaC53TtbTLG2CgdR2fQ1SzmGj6VG
zcTZRSLQKk1pfgQpQPEYn2iO4eio0kLDpACQQm8+LbVhZD1fENE//d8AHx+Jy+oDeI3id1+rCBWB
4Pkj+dUEERN1HJD/GVvIcwDanGCGTixLAb5k31LRviqAQggOv0gGl7FyuFzuiK7/UjfDhgzfWFw5
tM0Ge0iEaklCQp93IrUjvuAxAME/2oOZR6tuM9JHx0KOe+vWEJUPSSh+XXR3JCmR5w0eyQN/bAGp
me+BymNs5vYN2rXz3KiF+oehMgapB78Yc/ZVrBklbxF1PYN5wupdZkpjhjUT/EreNy7YzadHS4PC
g9nGj/T7OyFld0wckCI4XmIxm78Gqf15WKkOGIjpiPcpyz93cDcWu8PAukH45CJsSzJ2YKl0Dkmw
tLKAQIYZppDvIQpmlVL+gxRoHIp+VPUKYbOXMB8yDv0kakIg/jB2Alw9+4aKeA3djSBdXwqRyM3N
mPWwQkpO1CnhsLEVrnxxco9Ne7dbjhkw8fyyjDHdGoPlq35HUj97d7wSQEs/dJD5Vv7QdiPhCYH3
V0FisymPTbPFLZEffTGqr2nEpQ4YnvqqMpM+Eas4ZArV7Hy8UN7YUGlmuh/c0WQlylUuwbdJIdJj
Oe8clzNSGmd1y3bAccIx1BKs22B32psF9f0M6kNCgAMQhX8c0nHT3XpbK9eKrUgwOctDG9vBCanR
OHF25wkZ4sesuHarSNiqKg6irbnTa1nJsmw+Ud+sYKh4ct/KTng8vQ6mkSnQhgyGYSAL6hxQzSvF
ERX/x2JgleMwR3BGeZvudXoMBQn677LXRCVKSpWOAauZ6nnTNymvuarLhAQUTQ3zyGMp5YnAJvH6
a5qWRQ5MA6VHJWvIkArFjy7zsgLYYY1M6MsaPR4DO8YmKq2DDz48w77W7wPs62QSKLK5HI4j/xh9
GABoYvVqMShMKPazVPBaXEtL0Odo1WupchKqUtqMraynRwWI1b1FZuR8zltClumEZRxNxKNd1o5O
7AOF0qTWV+9BtO2SgqQBdOcOitesFmtWQBqyOZ4eywB/Uc/NAzEvJJvKXX7b9tZYWshcOip8x854
AFvwRP7vZb7yMbo9gY8d+bWBkLpRnuDjH6FBhm5rNgoc4zu7gouSZ62XYpKCpWbJuDu6IcFuz3nl
mq00YyJC9ToOoGvL48d6HpW9z/hHfHnPmpD+6eKyjc3UtdcN6S6TUZyOMUd38UgoeBxHZOSfhRcJ
zp7QMxG4WnkjuKPh2nNuEWoEgNET/49p7W4DdqLumdPl8DTaVL8OGMlMH9sz16G3u9vK+obYgfvy
wEEo3CKvISTYH+2YApdBeVJBNd2IbtK+1gcDpkHybvIvyoFWp/uuy8Q8foavHhimh6j43n8luF+6
ZgmS4Kf5cX7QY8ITVHYxCkSHFX/Z44VYtF4Cix/1VEEIfKX821ViPf9Rqfu2XZb6s3Zmq34J4r5T
z8DnzvYAGqH3E+nDL4JVDizphMoHvmtAwJ/64E6zG2OG2heojRWgJPh3gazjRQmkkrDTgk6+ONjC
9cHOET1nI6qQ00hPz6dlrGCA/zHSYObkDwxaz65OiQrgraSXADlaw2uevFyr3uNEjrC9+LIRmBLI
KGqK932/lerQXXHXAyeG51K497CZhKMHNK65rrKHSTHh26+KV/Q7n0KhvgLy33R6kEpj/wFo5aur
PzrmVg/ANjZdTfUqZOcM2YvHMGOpaffaChwSoXNrP1VLC2SB7YqAlDkhMRcg94xmllUkwjqzWSHW
Y4P0riTApAPQvCqedAhLcyLpMrjSg7Hlh6Cksa1iNanCfsHodtmyI1U63NdeRhmyN9bfILS1uYQz
qcodibX51O5kiCPoCa7yFWDhrPmcRARXweFAYqIxbBB65rd3u2TARBpgn7HCPqaD53YOmx77ZJFz
ySlUZqc+2Q+dQnzghReML0gBsI7zg1jRaIKdR0HUMbRNVnVtvxLy5gHsNJ1gh4AosEFM9zLYN54Z
diPTwaOFQgVPXLfv8sJOPaUSLP/8vtM5SIiCuiz0oz8qQDGzCfWYQQ5PJVCz5JzNYH5UhqLK/9ka
yv63zrU0hjYpKhmQwHyGCB+pJ72ZxNwHhvo73tEy2xY2LWQjBG9DV0WhgldbL19I7p3XVtCf0z/q
Ox6ekzlsbqb6UBS42x9bgcq+5uq91AqsiOR0xIzm9NWYZ8Cr2eo8rJEh+apzrkg1ZT9NsQQVUn4l
fHrg6gKd7vtaFoYeJFdoe/iu2Us5dWtJr7DpDF4M2wnraaGBFdiZuJW5HG1hALoPTEQKocEybUX9
wxldRJW+DxnHiQMqkOnvSrK/p3AWEerQq5TQJbSS4f/bIXHm8MUJ9bjGQdfYxkqyrHd81neBTu3g
yuhUxNkJG6XfPebLyJQpxlO9+8+2XV66kRp8EB07GUl2+DfjL1bnW9CHSH0JenCmAKLb0/iL2E+4
/tfJPLI5qrSg6XannjonLyHm2ADoKOvwQaUo73u1eOIi7iKrxp0t/eKmLp4zN2g5lq8BQMBeT7k/
jjjhu07ZR7OUm7iX8jivO4fhBBLaP0j6TDks0nSPUCy7TYGpKanUOPwKw+pgqvtC2heMomE6/FpE
3SgVyAFKGk6SC7Cp5giot8DtmeIItGrnj7vM9/VPQMJr+RSboaFas8zXBVaH7ZXbH3cKn3mBdiv0
/cVJrTxfRAr2JnidDOrbIRIcPJ1E+Sg6AN/ZLo1SPXnawkek7WJ3ten37JBjZBhwUDzZ1waaKTVV
RCuRk2t5nAW7JWpBLx44DovsrKJAV3Z4ZQLJ2Lr+do3grscVMmtCxNs8UlRH19b4pG6tYwt4C74C
H9qBI2vLJMxsaSvWvSdsWLoIn5iKaknaOivpaC/Xy/mF8Tq4rXfo6akEBUoM9CeIETlzTthKgFNQ
oFbYefOVoHq51qennNXSe3GhYRAJJe8F4NREmBWc2sK6vVOB64X+X3cS3NTH45K7TAsTVY/cx7Il
QMZb284VcY7xFsaTxmRKhtxfSVqqbnIKtmLIXqidLz7oBc0dY1GnqtbgTkGmo89MWXD5lCfDAsvF
Wivuqg5Q5Yz9H6cxEL3aFbbhjnqO7CGIR+/XMAwTKTr+uq+VM/doKukgMR1scRy3avVNr4MXpOXy
qa2jTnpu0nQyZ1KLWk/eIoIJBxptRmkLlbCc5ZYMYlCafXzpxPezCGF6bEIEtFyJ6wma63iFj5Q+
+5w/ZOoBWGerhysRSuXv5YSY3LHpSZBCQvkjUs3gdYY8p/A11jG6yNZkGo8pPT/VJmzL/63yeptc
Ri80ZWm1U8oFwSGtswj5AsjO+bKinhf7d1ZJX87fgtFtwfqzFYVkYHMufVm1+V0iCYfF5sAitS7i
6PpzarpaZ+qfpzHI0FN4F4+hdCBZnHtaPPI5uc2eGC7ILlG4642hmNkj4gQVowoC3An563XnYIML
KH/Bm5oIl+RpyHKauJX9Wz532Uc0kRMA2kGsuWQKbRyHZvqNM3PYPp4dev+5kM0l68tHeciRiE7q
50ghREdju0Sb9bvS1XK3HK4xR7gwK4p6eb4c0sR0wUTiIXx3ncAe++lMYWd4CedpPf5lVo5CBSP8
mRfx9WxUUZa5oJ6HkMGUKoCpjtjM0xjKEanLabs3yVekmBFmnv5L1nf51I5J4usG1/WhlFQjZbL0
yD7bXUoAgdaBrT4mFQGZFqm1mJnOmwf/XM3+G8Hbf5ndz4uYuIj3JX8os2tET8xG30+IjBsE139v
JDiIJZo6vHB3eKlKAFVq5hQ7fZEYLcwJ6CI16p/SkzDPmb1/lqQ/0K3ViCq5KvuA3UzADnwLNPZP
7ir8lRb+w4UUP2eBg8dJlWO4W9MaJIKPBqrL9TPe8Yvd4JMePM6f85mflP/30++xNlUlMEJIV4GG
+KeVTTLZs4LMbvHknY2qLAaBt3FXlolYyqEZckqFhT8Div1sl5ydRL6ZX5pvb+F5ubQHTP2I/bMN
G7bi0ykM/LCBXZLdVSDeBNy2Fod/4Qm5C/3QenMki4iePGHkZ++Z90hxgCaOTXCrkqe1l7h+/RMP
p+rswNLjyk9xAZcHE5DHdu9axsi/v4bkODPnSatMrff/pTp9YRgUNcCUuL/xpsqnTLxvoY6lR5go
oPVw8hC2VyCtU/rKgPtYPd5fkQZi0R/pTAdmRQU+QKkQzB+1USD8HwW1qdrBSUyrJegxMSrQUtN3
mK7teTU3w5IJyKaWBlnqqt6FvOh6kdqt/sftaS7UHDGYo4qRGHOqs0QwNuv3tIpZWDeRJIdhS7VL
A54F8XGhKD28h9W5YX/4MAgheN0gCQIyaNK+3LX2t1SNMzR81ZbpZ7/0B+VjrcB4zVR0O3cX3kiy
iguhOO6jTj+RaeDfIOqos7948bMyZho4o71RqPJ5G3u51eUz9p+14SDKlLxNPTq2PxmKIRzAefJO
VltydZ38PUTIDS/8r5MGRVAHuZuHNI57j6gWOJVri/oEkJ+VTNoWz3AOcmtck+RDCuyiOCvIlra8
go0UM7plLIS2bcY6OQroCN39nTFuPEL6kD4FTve808fhe9Qv0d0uUvNPn5An5cDVPGVkNLNk4rlY
gUwbduHYw2M0YtqF+W/HSdYKE1Ym9fDqfjQ2/GVEKo6FekOk8KCp+DCtGOCC8eoiFKuoURYvOrnk
VNkWJKBrwqAO6vQLj6HmdfCBHTqwygFLoOGrpytFlUcHtOsnwuaGok5tyM6yaIP56rXZU0axpLsi
U5aGazNnNeMttoDk8ChwOp/dyuSWV1Bsx9RITer3beGGn0ONsafqrG1Jm0mrQujxPe71FJMk42S1
s7oLkYAf1CKga8Gjsq5uKaSYm6rgZtJtOXk05wIm1PwQGfHs4j8D1Rhh3PSwhEkCsoVjkdv9ecib
AghCxMVgnTyyxeEduEr18h2Z/kQRrE7lqiMDFRYw+iWFgOOvkFvXbHj2x+LxvDBhteVdow4Rcjy2
UNaYird0mBCBPJyUr4AsoAAdmMMRFj1SefAUM0ej4ncyd9CjcijDYcCQLZTlwx8KhHQuqcntYeeN
QPg75++fOwt/xLg9IajUzaI0gbY0tu7MtnOFa38l2qULFA0w41B/PYwcgY6WBtHb+CfTwEPIqSVL
lxBGNonifmI0W03OFLA100tCSURnH9YP9cRlufEQwfKJu/vSRXjtwXMFAIYvIjP3S3yA7nYlljK+
19LOuvz4nHwFRCOpmX3HugElHm/WU+WKNzjPk7siGbles2/6WdBy0VdmtisCK/Npg2jlMbW/xDFK
IuWgjeN2BR+bUnLlD3FVd3ckq2/Kzp7o5wOlHshyojhIYu735VUE4Nw991VchEoxTySOjF/3o7ri
rOCC5qgkXJP8Qr9iQKQ/luKiIwF/emP9PzOwb3EE/qtJtJIInyiwgnqeCK9HqIvX2Mao9ugp/aqS
D4IMjl3VlCaB+mbpPK530Tbch8gnvbzVg45yUr541JHxt/NTgkjGizL99xHGCC2zBq5IxVls4ufg
YfzmEFiqVyPgl7V1XI49nFnnQkqO3XgohNVEO7KLS9WOPwRXcDkxxvzgRPCzVWsI6nImixUH/aEL
3Bo5XoDG/1mCI5y02JdJMxGGge/wnF8dwtdQzP+aqCWQskz+U++P7+M90P/qQvpvseCTjNiJs65S
3/RNeEZC3poL18898ZknJzY+s42i83bRiu/PHGjB6Xa0uQVFrFvN8aSFM9FUAZxKtrRBLM0ThVrt
cpF+wbwQ3fld26IjmY1aVTGRzl4fHULTQSzAFvrXcmMubIJkDB08KgD2r5Vo8Em0DVq8eumvPmwy
9TTpYwaMM1vpAzAmqvtdAHAVOGoKALr94gAyKq0jrJOXAAJqGbAVp9vrI+1oc0pMqyWpQnad1o1q
smKwO9SAAs92KADNnygzZZjdIFxKgJSPkMqdhi1fKEX/B1hMS26uw0729l93p8LvYGpCnh4HrTA5
CNWQPNXfesPzB12/1EY5G4UQS1ysjXHUqfEiNc2LfBrAAFD1Zs2wsUZHj7n8oxlm1+e8imkczwhL
sE0k1TFnEqaLat+IK441aOR5h0q5LDkKB7aR722wpPVFuuiX+XYQ95K2Glm2rzaqIBm+0c0yDKpr
siAIPysrZwEcMA56B4UXiUJk6f1OPOhpAxB+OYrHiSLh9/QkGcaQp8D9RqmVDkvB5VCnhyygCCXD
o7ezZHW5ztW6at1BKufYDGdQk5o3+pwba94KygnBB34/pVEj0I2AO7Q+hRparGUqq+LuBovmTE2o
6bVcCTPKicHFkncr9noGhB8yYlhL70zhZRyNR72VtP99U6sBbKMD2uSlkG+7k9Dqq7VnV0kGWSWA
+sQn1csn3xMUT8GR7/t63hl2AH/U61VMAzZOC+jyrjdQahPP+5SE5w7Yhr9g2s4k81tO6wN2tPOV
dUJuNE1PbCRgU+/OVDwNF02BjoJtMZwx4CG6IF728cvobojqSh1o5Alsy3pkMsjIn/Iq9w+MH1On
QaKjjJwuAFW2kvKi4cinRAYZgmLzR71oxZHUaeEarxR1xhVMl+5eF0kPyCP4vzIIedfYSV93OpJA
HX5/MWLHMjktaunnNsZxZgicDRteqm8VhXJbF7iqkStgzenk/GJqZnlEPPuwHplpmlegD8lnlLqE
BzPLLWO2wzOXGV4+3t6SZ+FF6F3NUKvOURzSjzwZdyJGCvVaPOTB8fmB+5BHQ6kFEFXOWg/Oj78f
3KYgZs+BrPY+M/GptDAexVCCgWuwAUqhqGxQm6TuqHJrI77KtMtBXQq8SOe4//i2KtrTp6vV8Gyf
qU7Vco9kAV0B/igKCUuxeUx+zDDc4XBzc6apqs+2aoscWG70r3XuBcxDNNaU6FJD1h+TviUOq0Gw
4KauQNMtmRztUhjiywUY1jazc3Mc36PTaWipBZsSQMtv+l/nSTy0UJG653ukaZGz1a+hJM49gXMB
eaR3sx2azryqyCEOp9yg9X9asEUg3TxQ2hgnmS5fVNNnQn5KK8iQGV9uCBdNvYgKR9sjzJWqMmRm
Hf0bG4Zz+Lgr+M1BprxX7yyV5QibQiTJ0v9YlY7Uo3dgNgqKZyBWJ7ptrdqeWFPDI8kP1QkBqvQP
l5L9wNygbPZ+1RhtomrW2ZGZWLJD0RtF4T5orw7ZxNtGTnkXg3KHG01osYi65q3pm6lDQu7zUJEs
MMQ/OtKAQUDNv4ARGUjZfHWGHkcUme9ByehSh7S/TpBTNkmPQCcocWeX6GmrSRY6dk4OgEgljorG
oygCYPzdZYa7uo/u9bmUj4hvVg+9jsyG4GTneQqAykaQDjylNQWA634AvXCega4xpnx6pOPw8x8x
+MLuYDdSZJcyl5ufhgxbL26lrs0pHOUSVFi/yGGRcmgfRlTTYpc9WWBO0zTNRnH0YqlRv6G8DQHl
GfEZsnKCY1wrjtgVtacSstfyOqWxbX7UR9u7h+nIveMg7DkuyvuEWqh0jXUnNxh+3QyVAMt36N5C
aRPUeSHGBBUCqc+sRHB6U2pOlQp3ZH0K4KB/cEUm+FwCqPEO85+ekvXHBRUIYW1kcEyNKwvoSRWI
0OYd1yyI4pCdGOVx9RP6sb1o/q7fKfwi9r196DFmHPZI8QQatS1BxxlbanKHfX1EenhkSKBZfx2m
s4R21qY+W906ceHSFAZr/xHumnTgcDb0DrUFEa81GGjy1ce+XZjrXfvDyVlZhjXH/BZWxslGDVPY
GZYLMjkvEj8lcy17EtJa4nwvQJ7Ey//PLY7XoGgcn8S00yG2F0j/dV+XKPqs5fVnK+ZSZhDB53//
yvDs3FaQLWyJfQdb0xWUINLATlH04kU1A5lWnFHRGWpD9xA/Zme6VLP/8cX4gWBx4RzIW0uAo+MG
zFoqMW9v9MFA31txbWcstJz6uOuMW4FcqORSXoLau6SweLf6NM4WB9D1yJ+gmcm2GKY6YCValnat
m33qTWY+Qfhvdl0yDu2ipGIAHk6pmK2yN2wM/TDVCTo6vBQsI6vZEqT2ccK1EP/+54Q5HMDFh6yk
GTMACThjv8jfDbsJDVBEN+CHI2MXufXSQ+hl6H3/k+4a03xtDi3fQQF4c3BBa0AdBaGjxy6YufGD
WKXR3XQnXxY/9VSxquB7IrfF20OYt4TOKiaoAtGOyr12bBJqdp19ehARaO6DhU1NG7h9etYWgNRh
w4nHNjCmVVmfXyeWCXP+OfjavOkymQiokbD332L+Ht+knTfHbclFD0PYui4iROTputLwTUeG6yda
nHKxnfuxxT0fJ0Sf9DGZj8d+XvSJtM/XynzLxJy7Rj/LqwvIBNwjHlvElVSiEiMUYNOaFv0LtJln
HdO6rtMmxWn70oyxDYVj5ynUdK9ORnXfnaEIKMy1S99Sp6URPZKTxAM97CdoW1zoNqmWisVfZLe8
Nvg2adRVSkzhRudbwq6ebg//SPRtOS8e2L8Za1/2Unwld1DvycuEGPNBDlMEAypSAxDEXCYzMO4B
MSdg6KVjUAzJlWXWrgm4VWU2aIkwXjv5lvvcU50Pk1cN4Q1QD0vLg8tgC7hCShjmhnu9o/C1J8kt
d+tQzn5JM/KniYVJxcDYLttED1tdctHQVKLxrNZOIUjyTsF7duVMRR0cUwpSG94Xw51D50NYtsA/
q58TdAIWZxUQaSegJtSZmijqeCGIfCn1MiI9HFz+LmFtjXL1vPPFYrSWMz3PPqkYrqJJYUPVYlFa
0nPurJXEghU6cCsNSGriEDQJaivLo4yQUFj7U8q6obBgqXDpwQGF4jwOB8MxpdfRWlZuwsyvINk6
3f4uZ1JXUvMNttuLY4tb0iMYg7i5BmuTcez2oe+5ptnU6AIRKxLCtVuGKPVHIAWoTkJMbHXltJ9c
2zLx0XMa6SD/Gw6t7BzFNk7faVOyZNsFiwa3ad+zHOcxfX+jSXcMHyHJ8B4eKwX70Zeae7pJBRjW
Oh3dCuws2JHWuWYr/QVHiSLzSZRs+xHSVmiBCizOOkJ5qVFz3ecjq2CskRn0vY4cOcPR5OcyJ5cQ
Q9HvVijphSlXkTC2GV7vFWl1STlH5Ttc0jlM0C7Lotfx0gh3VuoosejZLAx8qwW7CzECpSzbSA1s
iA6eS71QPlB29/r3odCSsvfBUjBD6u1jZXGPJfHsGfwn80GZj2kWMvJeMBEiV2vbqeJglM0PiFrm
onYaebPahnBpT52MjtVWyGjbOesH8x6dvln2ZBpHS5goP7wkwRaykDazxoLgVm9FqKYETRqS8duj
QXv0w3+O+C7L59P8ipUxPmeBePpTtzAOKIWKggIihNILY6GK127FG3OWEtnbk5NMwMIOvZ3TsnTi
+DXwq3wvLtBVxrO65s35dUsBS6H/rwY/CVI5tkzEwPcnIUfAW+tmobSfD+odFEcQtbGrFK6G5f1s
ijbp44o/qmzTJT3Rjuv7QDlUmfN+XPvoKMyX9qi/L1VcQ+6WZmodCsf7wtSNuh3/W1JP19PecLn3
aR9e2Ie3Xy6iXLBhKX4mlN4RfGkM7PbTQ21auNsZwGVd4ETfasbHBjZpf3SzMOSqHUYHw0UV0ccU
GK/QMaoeklYQGJVqJs/16Q8Kz2yvDF9qU8bvv0HA92+FtQ19Bs11ozkRoJw4WhsVdNXEC3mS5jrK
KGpUsSG6BZF98/SMGxsb7YaVoLbSkprL8whjCirjKrqXxtOngXCtmScbqcitffgyJ3jN6z9vdlTL
Xg034ijnXbR+Mxhr5WfQ6j4ziKXwjUrjDH/ZdYX8bOhmp14EFqg0HHcjbKq9ZLA1rRmN2uFHfYrW
q+agXaYF5QeK1iMXz098WC0uxnaBETs+TW868rk+7I01q/G73VgbXdE/ObmtV0Xb+yv1eIb35gXc
SwILrTpizkiHBzTbo1Vp+trYzcEsNHaf0JeW6o1r6MvEm2puiYHJ4qyDSNMgNzVqvMDBSSdzHI0+
f+LL5dEIAs/TPZkpixmEt4aW+SKQPATVL8kI7am9b/2sm3tFIaRGAw8tnw43peLqh89e/WhglpmV
emPdN6g18p7b8YzJvtoCcvl6PyB/6BaUkh/+b6PPjIe8PIbDIonAtXVUcWWu+unwAm3fxofyPeFM
c3o+TkQh0ZeZ++3kWvh/DIZPMci2om4gHOljTkH4kT+LrJXSilLKuH/s3RWo20bWB4Ipr0NVwjKr
HI2MBH8G70YGEuxzdlTIE9gLw4vvRhYXr+aFi1e0cqX8dFKg1Y/azu+mH65Q6VeFeMm4IBVSpJcy
0Nj/GyTVTc4ImfK5LGtIFhMGMsVE49v+QtFU+dpyGve2Omm5mFx2iDqGxZzqy65UGvzpb86VMhEj
40e5eepifLBHnAZsTkOrLin2lBbkTMWg85bJSCiLVALEsCedRg/VtLtnEvSExuOrqy3JN5DzQiWK
iawU4+px5Qx7E7ZcvAEw1rT0jho9uISh6yZiF4WMqIb1jC7LOI5Ye3sU6jPzygiHZdqkXpQU9D3q
1O897J/SMEbSCjR5bl3yw48pAyI2nceOl+SKksFAjlWX6IqhdeS9Qa+OgrniYQnkUCo9BEOguuVe
2x0m7MABtArdtpM85WumXJIqQKVwnd1CjJVg03y8yLCusOsCj7y6SVceqYOMUlgYnjEtyxtwmu+C
E+DbfcYks5Bil4/vll3d9zQQiZ7IT8MWWhiKbGoAruDAmgRrcT6E0TmlZY88UZXV2f5HXEV0iBgq
q6617cIEVmOgARFZx218mZnRdbTcWEkvLM+gY+WheJ9gfyefrg0PaY6Eeu0WR76cGJh/PQkTU+Du
lBjsxnW6cFtgH0ELzjKdSUjIf3aLyTY8o3WLuBDRDIxXSaNJSx2v9UTny1sVzqtKda3yO8cSoHSb
tZ0YnYufob5qYTUGtkypzxmvGv1H5Q8wxWR0j8FHcd3gVX2FB1XMX585nP4xYaPcNvCAKAzqKq0b
NQQ1HTz7ALO5zTTNrjWUY+wFN6jkfS/OyPhZ1/yqQCHVGOUA0Id7i3RveOtTY80WZBzQzMpebsBq
9HvovzTrp7adZMQTC/PTGTkCuQOkX+KVQ2N3/6IU0rphTyby+5OIpk2IxdgvYkSFRBdn5gGLgRqJ
SLgRkkVNihdSkpjkcsV9ZVFwqlAiP8NznqoEmNtou2tlpYmVjXt7h/NnvB9MvYeNYT9E7mzO/8wV
zplY+Ib/A94JsRtn6iPLjrrTjxyyhjfRZSOGUkT/n3v1qacKD4fkeNygMyY2CTgQTxolZDDFl/uo
nPJoUGOxvuhaAv7EqEjCskAfNSPZ7S2bbzIFeFOAZP/i0KvVUMBSR1qSJLtDPt9RtuEqs0zRCbsX
AOTBUAfc6uWXcV/h6fKn+rV9jgRJuixlVgj4FFoRjq+jKB3WfStqyfgq12qRX5GIadR6L+ri4DFR
BL+jE8tJG+UzVnGCNul9K8tfoDq3sMC5B3O1SMEOg4CtjY/jF2UGVS8TLUhVDbA76uZ+0biLfoua
KmT3U/JWm0RkcWuwBhPSdJ4Wb70wLIbyn9/aJHieXGx99zlhf/Q98iLCInLUcNhAPEhw5VgKPsVn
7sGXMzXxSjkdhl3lYHNoIWGv63UVOaas57pur2Eqahjq5EUb0hRGc425Nut+FAdqPkfb2pfKefHd
lhhYhYt4U2Df2JtCS0ANZetyzRaOWNqegdtCoEq/bPJ5HCvTyJzVbsZlmYCX555LS/yf5rxuTjoG
WCVLiG0L2zZMGlC219+GmR4sr6FJ7mBwQoz7Qn8Uf/G4OmvoMn0eKsWA3SVhKIBzpEFJIOFy0CVz
2GfAfP/L5FiUC/tOgRJx7R5dwJTj4LfhgiLRn5hZYPKRex2aDsb1+bc4amZcgFt6RU4OcTY1kjVy
1qSwVcBRmAIzrnBIuvXWBlM5ryQtgTk7kDUYSIy626JdSAPAJzw9vY5uuTJfNopaPTcLOLt7U7P5
baqZfbyQC59jAnk2vvIsuRw+BH7nuxdeqlv7IUV6aJZlw+OmeNfI9A1NfPfmSs4HiUtSqfoxPIQy
/HFur+U/6shzZ9y7AdHBKgBxKhVY8vWmoelIYdYNm+4t6KRPejJV03ihD3KwnsGbsZNDrGLQb6/j
wRuB5aWXME6IslPD5QXiH+Ep3bKjdsGv0c3Kezm4DWNG06C3+JVa5jbs2dsT2ry7jtnlzf2caFR7
RScez2QJ7drxzWXIQuHsM7mFFiGaZNYAE/uuPrWpLsQ5mVtZJ+CtGkpEuAfVIfE0WSBzyuy39pdB
BWUGk78UM5uCdUByQDkwWRj4VsyST3MPZMkxmoPXzm1Mt98NTvlgJ8vJPxLZ8NaTUR5FdW/r65aj
GeQoxJ4lj8+k+0IJqhP5QjtXtngDq6eHHEseOxfmjRekQaGucxNWMs7SGbqAbtsWt+A+t4NoIJpW
UuiScDjSIdyPHRCIHfQMGRb/KTsentBg4RZk4CeLBQXKnX3TCceETgAv1RcBdHkDVxEgyz37r1ML
Glv4Mn/PxOUg36oSQ9sArG6qb9XE1g2hDwY8XO+Vep0JATWpl675CQ/VBu8jrpvZzaihFVpgrfE8
SwA1PMlkL9zFFWzlsJbYNALYuDe0yLW+KRjy5659AberwPNRg9wNxMY85AysXP6hOYb2IEZP79XZ
Qy4BU11hre2UIOJtiiIbUWNgckiFXtQBAXVynQ6qpyuF0gW9HEP/3ZIfTcYs81W3MJPUElGZ+5ie
Gg1TtArBjWyUMcgl255BEbYaXSBNm0FZ7hvddhXggoi1zXgBZE2k8zzB6JcCbDNGWYiFsXd5QN4q
5/R8mCGrkBt3o3LzauWOgfcv3celiTl0TwtmxkL5KFfXymBlLD0phOSTspllAOSxjpQ3d/lWicrP
494GLyPt1wIBWuoCtfsv4Y9fYur+l0wi8hTXTdTAAhDZX7AKnlgo7dkjDALHb23DgEMBMcBsiU/6
uoiqTCqioTWhnIqyyzYM2rbLrjOFzBse2JdfV88EKPYLxWUqRRYwhX3Efi5MO7cU3USOyx9XT73U
XTc/bnP2f6hGXMId689Fcl5hlwwc8T7aZT/F41jmc9d8j+Tue62Uq3Zpui5Kd9bom2ibvIATfj4s
EERCYk3cZW5zZgOH2h+yE5kFtwc7oSMnO2Mg8jXxFIcAV+FYsGr9I5xnGQfFJdqVanGHCkJ1wOre
cXaKPbyiZpM58vF53iUaMqC+ZHgI/TJtHOZzJtmzJybrvropJfxaq/YsbgR4GCo6kHrVf+pBLPT9
rJDMXTNl5WZnvNquo1Ld0/WxGXZxALtY9qyEx4QmHmOpMXSbKsMkSOwiRu4mBZKIkZlRBgutaqJj
UhCCEUxPQARD5jl72+P0gF7udIhJ0WP3JVdWbzjEP275JQoC7T4PA1ZJEqsF5mJm/zt8L5JQCD4F
6+rAQicvd5jxSmvdbDJ9nA9KG7AKYrSZ2TBSUvVOq1uo38JXOE5DRmBfsm9DaIuLiOZIUQbEfusi
bPEjw4aLCF/9OuNsb8nkxpzMxdPUgJ25ThV3kBZx78ShPlevnc4bJVZbXsBPFczdlyDP3IawklxV
HR1L767lmO7cBlPdUHxa4Z4wUJ2SjVRaH5qPARnMXzQGl7QVRH+1yR+xJggVwyQVnJPXApY8UU8g
vMSR6LXxE2EkkA8wYMRh/TlenJdSakMoehwBlTvBt4qcTamvxBMH6ngt+VUC4NWyM6T8xH3wOwT2
tNKzkzpK3iV58ytwn3XLlhsBKMf6ob7gDeWAwpVJZnnE+aJSqw7v8X0tsgapFmlLrPAyLZ6ELc6x
eeuST4qoR6EuSw3KPkxom5j+pwELEXAu3bw/ZM+73tlCbqppB40sutoPhLyaZ8+Dsg11D1UfgWZl
hRuPb7fIvwbtIf8OiDGgaxYt1zMziCDB4vjTUGOaOol+0YOqnrkA/qF8WZ0M3JQnfCarugpsJo2/
SBFuVhKz2DSGCmAUEtjQrMx0dj8KRw58jnGXZiKqwu4UkmcnLNEPOlVV5VB+isCXk74h/jbtVPty
yvmOSrH4961phLs5WmwH0ZjJE/bDw+69ZmT7IljTkwj0DN6e4l+8mOhrujjcYbdVpbVexOmGjs/5
UPblrMNeIqhFIhm8mLaQP6RNrl8dOxsF0Lopnz0AwCRFnEBYAT4AqnFDJKOG9/22V93Vk7+U9ruz
2rHQqPSDsGzhEyJMqBd6rnUp2In93bBSSb1OwLZSVuSXaee04dlqvXrXVqSmudjcw4AbUsRwVh7Q
v+oTOA+dZYAVQ1AeBU/PCGfTY60MYE9BHvMlzqVwXHu7tIMbe6KAUWArMw2mQ9ieMFWktSP9ikKp
drEAstZMIUealU5YKClQN9u+hqliTJvxY9qM/yt3vM+qrslvywnpZ9CMHYi4nFgEqOvbHxYNIGhS
jlKwhdvi1zdRdnFBPkI8PZvcV9XWglxyelr9aPO1wTBLKHQLxDIljd+vUtjeVEy2lpH15H+YamFA
ktxqi44AiD8BBfz3vLXN56qWKbl4RWeRYR4h/eiwPCJrRSxT15Ac/epcfdIBVzCzFqVjZefTJ3dn
sN4YQhG2mQEHIuN0c0+p8TKBYzDJ1JjKMrODgr9uir2Wq5IblGPshSdyQXzArTcATJZsD7mC3GE/
EUuljakxwhAZYUAnZ0JiUxV0EwzYa/gKCdtcIgOm5tgpYiy4zj3R5alA6CH7o5BMJtdYfa+VQ4tz
FvZDHFu0QlyycslG9klghllT1epwMrUYMdU+0oZiWkirFCzocrkMTAwPsvCBKIz5bhD7/0PWADCF
ombdtCkaGOsoRkj8xQQgRkaoc/bBTpOWCl5sufC1JN0mqc+NZbvfU7h7JNMODhJAMbaWwK5cBpVD
ANwRWXvB4K07lJodcxBENF65X9gnAlYgrutmjX45Y/xzg6LUDDoiTFy4UXJmZ/xrF2rYHphaGW4J
XxdL6gWUC+CrqOVt5oqVuK4uqAfzUS2oxLP9L37z8epp1fafz4xC1u2JI2wF6q8RzsF0HxgLsiP9
XKtNTsuMY9+6Jxmx3zAnajWhBhQXLndq7lTUlg9yzk8e4HlNv1/Pzcq7/qsGMHw/Areq0vaNUa1z
YwWfGcOLyiqvc/2RhE3lJp3ZZJNgV9ZnirsgxvEwMhj/rHG/tqaVsM5JDvWOAIxiQx6v1/cQUJa2
WfTXzkdy+E7Kyf9NiohTkeRJ0PjHUXeC6Lfrr8tyaYjV+t784ljvs6joE9gg2xeJ+B5MpUKJIbYw
VprVf4BKBguf0+zLCtnB+0IGIxWjzAJ9crMRO7YQk2iuALlnydk0l4pyH4Pv3kbBfUfZFsi3N0/y
0D/UB/US2aeHICyXqGRH8K3rr1iUYX7n3skQ/qKbUoRPMThbB9IWbs+NyZNhsTO97BjaV4NS6dJz
I+9K9BZXNt5oi3oX/MmuSN+jN7Oi5eJrRXM2v7g83oG6wQtmYei9YkR2mRtXdnvs544rrzVyo1b+
B9XiBS/RmASU3ZNvKU6QS+DmPdyJ9FcKAfVFZwShv2LoxCiU/sBkO+W7peb6AzCJim87y0ShpTUt
Nc8pb/KVL/pUB6FYfizes5UrOGOsSB/2cVc6ujSnr5iNY3w++tL+0lJFoLmQPFcIr9sJaTl0zWM2
stMUrHb1NRGgnYuEAAkhREbguZVfI7T3BI9dA+/QTJiOQYjnvXAdw4Lce6SiW4WN+81hHf3/a0Wx
25VVc8ByFckFBx7HKdLJL4i1DSztNIdE06LU87pSw1sDh21GAWHIiHFG+9tAQVW4UEh09wxUwqZs
ErFuJOkHevBpMPK2q1BlTkp2q/gJAonpNNIhBR8ckGciGChAGBUtYJIIvPnwVH/ct3I4V9djRhPu
3Khw59nVI7gXWq+6nSNWYRp0eznYjvxTvGAwemHNUQ/EBOAT/JmLtFT4wZOOXxf+RC9m89Fge4DK
n8AxJ13eZhO7BD+t2sLYDJ7gvi9BsESunmBa2dXzO1uuUN0k80YgbRxh6pX2H0AssweCMaEjNiY6
Fu9Er0VgfpISfp/3FmwBqwjzaJL/p66aV5B57UA9k8ya84hUp93+0rGHm0ZmfseDC2M47h38e3W+
RMzhr1vWXIpxHdc90xJL57vSSdcXQZURo+RzYKOE/6atSrVdRckyVgZL+3fxTKfdKf7ZZOGZ9RNu
YMTTv9+zKRZgEbwdg6SIap8EZVL8nkyfIDpX0fG/XUBcjzkD9BTKNIe7JfOVqUsYzulPkUsEPDTg
JrcfByKWrWhU7piJFbsHi8Hku5a40AI+VxU/3Jnxq2hLHOPapLRxJxpUa7ogVTl3iH44BEYHK6iz
1CnCz+i4efRSg8LNwZQWk0qdHd8sdYANPRpxFH598nNom7dxBJipOynQsvJjI6RFL4fZeXZu9zNi
prHfpEIj7H1Jz2OsYSmMhQDm2HbdS32LlxK6Ts+mSenWk5RdLdvYT4Av0Y+NLc0fjBcj4lZqUGeu
Zg8xD8xyT0q66f1fxH+4OesLyZpkQ6sWR+vbl5eFJrBMDFBXiFY6QV83g7qXjYAm+2HfsaOWJl9H
FKOB/z/RBmINM9OOvw9/f+z5m/w+srkpY/MqvR3W4bGwBMNuVJfNfMekYD+sfFubVM5Xhdry9WQ1
u5c0cO5VbxaiwxT5drPyAainVDyWKcP0zgKDOJHEoJSn1hgKu+jPcx57GXZy9J1blw2u8n+5O/l+
gSriCGXpTwDkG6yO7Jx/zdUc8WAOyMHJ6TRyd9NyBjHAIAdKysiPgKxKIi4uuPoDpSe0hQ6HTSCz
hKqnMmdr+k90vRbBaxk19dCY84Ym3+9/rJBvVHVQmuYGq/gWXrdOD1itQQuKorKXIYTeoKzia89i
oRnHesIkHDMQ2u8TU8iRIoZMtj7TXs9l+GZ78kUZvZSmdTGNu9kOBVyiycyTGWOc/2C5zLXQivSs
hKuYJsueunv+45lqYGKRcHhDr+WkEUSZZJPquH0c1IZm5PjBcnuK1ZKnTWGwOlzCSQQl0LwfDMOn
ejldK8+GCu2EBJ/aoFJefCwDr4krbsYirORRUQ8zsNiVUK7L2WIPYsxfTz4rP82evOJX8tOu9shm
OnNKFxCdl6d8Naw6cbmefJWQ+xeE+BTSddhcDBeY9pQy9fyMx8TfkPcueNxi9Cf5GwVrvBqXUWKN
R5EBmlrJOrJBXngmjZRqY3CaQ2ibX8Zai0OqQzGSgQ6hHLrwUNuS6nZH1YLiw5MrYo3knj7uz8DZ
DF2lGTfxZLJ6h40rU3S6v+R2xwOkY5u4NFf2IgcXl6WsJl8uZ3QxhnJCj4VSuchFvJd4trEO7wKR
3SL4s+S/ewBYWfOj4kTRFCCpiN0ARqW1frdZa7wuNa31Vs9wdRoFcNaItOS7y+NrfUs8GTQXBjKJ
Epf56RedbFI9wYNnHJuWtQnEDNeEEPKTTLHZRnvT3vNCNyTey3yrEuI4fVLg4ZAWjqIiYJZXM32X
Ltib7hlGVc+smLHxELGYIT7LV9lHym8PBSNBWFvdc4bRC4QMAHkxXLB28IRCYLvdvJjRboTbspb/
IUOP+jEOg88JP7p6qWfdaHihUYOSrTGkv6J9Rr8IB5dAq0g/oeS/VVI6drr19M5VLOcTDTsyeYKr
Hd2Y9vVvAo7IOnRPBB7mhwS4q5aED64OL48+E1hMJjoi2oTopFwsDxBXNhX1L+N7nSnQaIz4onEX
G81yF03P3oxBAm3oyObwdtLfW7Ol7CrGj76S+ou5AEW9UIrZryuF8qKRGODQ/aARjj2GfcCNwwi8
7qNhwycRXuY3Meib3pmD4Iol+xJrp01qNg+qLhJF5J1zkm69b1kZeSdTGNsD19HGDH7KBwNlKLOD
gjO44xOqZQmVpCrXSKUL4gZUwlE84UH6IAXt/6jlkZhGSiwnQNJ7NPs85H9jmtmVfZlpOOc/15QV
03NlsevIkV1jC/i3G7FbL95ZHuXlXPFhnhNcxjwjWqfR00edzWoPEomZ7BAX1ehMjMONMP/OCb9T
r8w2rTSJX8n7pJFudrmHFQF/lHC2PNXea7X3Fhs7wtuwkqazDCpjSgpL3IexgEn0byBdeUu45Fih
NbvDr9pKl/7up4xq5TcDEuYrVrhb4gD45+Erp3BnwrXmLJXSZFJzt4arNziPKpecDXTsf7wEFmTQ
cIRoAafbHsxArL09qneNVbphyMITWCvn0Wya2nvZhBsBDRvqdzK8cKOEFHo/bVvOHc1LALG0V9U5
ecdq8augz8/tjwW7NDT9uoO4uY+MsSWm294v4kp0wGw3mwGPnb4xc+3vJu6/HAoRXAfp0luGU55v
NKC6NSmXa5O/42LfH/7Hh/BOByfg2KIsw/3mcoHtwFnFllK+m756xPSFjvfZ5SxjfB8HvDHnk3OA
k6XmA3kUQ6yoGYBMacWayII2Tv9PBTWs49fSkxOBcnN3l+1dv7LqfJaRAPWvI2TlHTyF21hseJor
np9KR4JfUIJA6oyLdkea2CmP5TPB4Irh8l4vn8bwyp963/TZ1w8ub4Ipj7FbNP+NI/zgQktYM9qd
UilqKOCtP+dw/H6xpfgVJ6QVDbo6V2imopUtN4z+V1hSHe7yRo4yFKzq/dngssLhjr3y6Od+FUPk
QSZ8DB2Kn+41glju2wpbRl6wH/+nxcFUArCgXZjzKe0xf9lzLeX1iIjeuYxEJWuo5hZiJRjUOtGu
7fONy704I/GlreY4FqgpFUob6do9G+FNugLB7iY5qOc/rsrPl1jXZ8JG/8ZDjFxryUkpyET3s0+T
fdMBjalwDPuSyURT3vhX9igSDacHhJgbqaycdCjeS+pWvRK8fPcI08i2p7MgUSENujRt2IFbqCzZ
0WS79NheV2CKlcbkPt109WhhChGI79SRUj0HBS23QgVDunYV49ZRYGjLDPPFzw7m3ZQCRQXfZWCv
iGKTb9N5bDi6pvmNE5MfT/ZZjXJls0hWx/imLEzsJdZR8qG95XHZPWKOYCG2a/Aah8UZp+SW1GGp
ykbnaCBkivIANVb+WmZBauanL9x88Z2y1JqbUnGcHLuqvcxNYIAiaqMeHVMBzgrS6JG4hOm8FZQ+
SYHrRddzalQSfDAGyxBViQGszKDZLOR2Za/6ZUq/O/JSg3TXkOjLD+BOfEWma9WoPrfj0yUBsZzM
in2glQrlFGOoWAvQIE4tWlOQMd7UEFOULUS0vNQcc0MvngAYOhm1iqk58sKtQhnyCZ+MP5amQGJ/
997igoSptNhRy/0A0mKz6EpDbe+mYE7weEecR3Ca5oapH64hPSk0OIPYMyHkwQt7hTXwjItzpry7
JN35vNrVNFukIXMsY0HKNYdq1wxmv8tntFDyDXQD3/EHk3pwdbPInlSkxYSJsI/tu8CXt5G6qw0e
aBeLanuLfgGKUSH4qQ6h4bcCMBKZ1BChHdEFgXTi7SImWStdtXaS6A+ffqndXUi6Um2J5bn6GWeW
6GBufnN9Hr96c5DhrSOeczLOaRF2xUQvHGC4yhZCODIGR/mgmxKgiDc10NzmC8G4PNgiTphbhWy3
69jUq+d1OAygwq5aaB6eiuLl3IK5usGMEovE/0AsQFSDUHetaNNbcPWz7hOpnw8jVvtpMlE7DyJG
3vo+AdZoWec7Fzrtqyk3s5aJNFpGFnRti7NvkPtkKcgLX6yCADjBDoScjXq4lQ1L9pQJr3T5aNpp
9Sz17yFuQZpq0B3dktO368EgvUWHIOLAPhDH2mw3ozVm+xKpQ8u59RMU5OkA4rxTuCfXl3m5gRvW
1C/85XOvD39gBLg3qEAjcTu0C5DOPG1EQNr5FGRolDm8JgyplShD3Fo5eRRz/tP0dzg0Dxcxpdl+
UcdqYWwnAlRt67QIGUm6LPau5XEeshONIkam2FK6TBxT0vTOohT4qsZGknFN0QlhhjQLIfDdTyBm
QnTQ+eeD+Z170KYd7L/XWYm4vdMgk3DCv3sb0AUDiT2jMqM10T4Q31uMxUu8Uj1+hG9envlk91Re
Ok1pfGufunn0VFr1eggQwciR7JKwo1r2osqYvI7XlKPgFE+NapLymHu/0lV6OO1levsCQGoWgR4n
5I8RIQaEM/H/tGd7bzGLeKnY1VBihFn03J2/Yy1N4lkivo9eTKJfFi/BWAFiLHrSi+cjzgbHmZHd
nEPCC2IGMNgRHJlNEcH8Pj1sldN2OnvjFKXqvUvXNLJM8kuMT0qIPTVqObiO4g6i+oGxCzBBmo/A
MVMg85kpWeEVVbdh5zrrtltfpWl8jonenMafss8bD+h+5L0whM0UaxCC1lNfT8L6mrP3PB00vzZm
HLzAjx4vuFdfSto6KMR3PNX9gPNgpj0TOn5HaPfMqZ04h0wyhxZKlb0seKm1sUEtlrOpLBZuT0K6
lGERv8q4gXi2XaqUBcfJiYKwUei8n4zFjipzPaK1ItCf16ma84G20GcEkERP1FHs2YASmymNqx4j
AcDKK8Sf/DP6zTSqS1SYQzHlpkBXE9ITNaBHIPZUvLBlVS+fH+ldWce8asOckv1UGbCbkRsEbnnb
EHzaoqIn2e3n0O3A+WteauShbd/p8Ak5AGnDyXdgVmoDJ7+QjtF1wYZhM2hlmZKv/kZCuIHIyiru
T8HJSVN87UkZPzmsUmNCw4oNUXKyhxennYMAdiaGLOop2gKJu1RuKeXeMALqHl9GdtD8/k7J/kft
k9q1dfKB5WQe/+GseeBejI71pyfyviYBYzakO4S/q/s1qTAH9Fe5ciEUgPkzM5nj6pDe9edRgw77
uTsjsEcT7IgFFB9JbXqfrl57H2Z0upSoTltu4hpreT0JvfOrlQWC++tLj+bsVzZPfuHrpvJ6JqNa
PcPhxjq/qVkra704gnLvn3yiS8C9FGccM9eKkPrULUjjsEghteKBqn7p3GV2F6rq3UYIU5V3W1aA
cx8+caGVxaC9mqkKlEnVDXY7qfUj59V79bTCxAPZSg5Xot96MMIO0K+GR+XftixXppjcAhXWn4/W
aP/YC6GkexHRPCH8NAZN/ensiyGegZZXN1owejCWVHZWWyeJtpSSqZsLySBoHewlsUXYosOimzgz
Cv+d07p/spC6eI1DWCvDe1+uiSJJbFFnfOYTjPlG1xz6GavFf82EGs1ljpq6cL7T58nkhXqOq/5f
SGLGmTTf20WtRpvL8sxees7opYH3TEkYxCWDA9kMz300ItvqnTqxgoKJShkL7MtaLncYdXHc//MO
oBcAVdJDMdlh6a3jmAEGjXxF+ozhNLgZq+OzgRh/2wPpkOUJPnxdCnZ10hvXlA3rz76acUNpNwYM
uQLVDs3TsjpxI2W1GKC0JaghsP8/bmGu+5sC1qX3xMs4V0Rv7m6RYKni+KnKyVyvekctIfl87Ojd
2teWZlLhQFtRoazrbyKbuBNjKPZRUQNvOG/5afEF1AUbYxSuBPOcD6iA99lZE+uoP0foBlf9LCWK
xCQIqC7R5Zs7xZnmEBmG+qb00CPf77gVpHHfpF3lJezJU4OqDdZUALVSNu75fbLwUxyb8yDOpO8T
ObhK2bZFbuPZ1mafyaq591bbEayK8g0pj/COo3UAh2bxwgXC3ifExbclRhXKekB679H4b6uLec1y
fsGZ8XmPUKisXKPdtS/z2BtmIIOh8UgJ/iU2VY3vwXHsPojgGR9nl67ZXTevu9ZN9xDtZ1c6VzsV
7iJ/4U+iKdWe7N7EbtBJoFtOD9kPUNaUJUWd0YtC7HQBJLfyjki2tqcdxLPF+4o7dDGEyNICH8TP
Zo2DwGY7p0KReQ/CUMEmPO1RkrHbelAdvN1eAUFD2P6WK/y47YOU4f6r4eHTry9/N06MqwPJOjM7
a2iu9pcQRfDoQLwTaQGDLmaZRYnxcyF2bwIriNb62k5IsefxaUWIC3cPhCU2DMoU31Bwq9/tATy4
uD1wjCw1Jb0yuNE5wcACwmeFRSS0QxnmRdamG2wZa1yhy4tof5FMdrMqFJ2KTEe2Fo1Fwr8XrakX
+OguYrKmyoRwVnvPQqbXcrwakCbE1a7dS2dUH7EGJPndDUzU22vKjyCspl1dUHmI52vwYjWYrpYK
Jk6+fWMJJbRxWoVlHh/grTPBXX4cFYTP/pcufBuG24As9WCgPxasxAiRGZqUtL1VnaC4orHZ3Uyp
nSNi9U4PT1tEe7sYiI2UeziNwxvPw5anK5bBhBp+CJUmjjoHB19d9/LxzqZaUD9BPqbF9K3/cCru
5hupdmGdXhlp1BoZm1mp6Gtq4u7zhdxzutfw4InoclRXkoZVNBGgsm9Jrf4xhHYE+LLCS4QR/BIB
4Y6hsIp3+LN7aaTXLm5oUDBgGUYvewod2Ldnd8IRhA68pw7LK16AsJgkS7Wi9Y5qE79PvmNEIxzA
pLt6RmklpQzXsZKVwrUtLeacQ38C2VZUqjC3iWseITU5oOlNJrYe7tSdudaB8NOZrp4Nsis1oyJN
GhlYnMeDabk003YlaA67Ff2A96vaEt40w8a2/RGpj7XBqQn/6EGqDH/UD8qduZhLihlCQVbYEcE/
fNRx2PUNCLktpF7y/mSTkJ0oAsQ5MmMgl845C22ThNRgYvFHUwVRu+0kvamvzTajdYWEM0jzjt91
wUsJFrtaaN/FkdGyZwH5Xo/kTa6UR0AMyqF/GAR4cK1wWo1AmGvVIj0PfSVBoQlRz194FYb3SdWm
JDVyZg/Qdwpv0nVqR7z9Gqb2glHfFi51X3xhEsAOddXBf3EKUmbjY7moAWazmd2v74V6g+s+qTQ2
x2Im/r4knKQH/ws3NHfib3M98VmQFY2dBUDRqMxnAh94c36laK0kpVTTM5XA/oOUsRdktKGy1xzy
gz/vKIujtNCs1MPBjyjswOabJ6+1d0hamNFp45vuNTWRVXX3b5J0hf0c+S3F9I2zqcjFOsTBwpRg
dvCXYZsqt+a9lY2AtnSwmWKHnGzSOwhLx8oLzJiS2VAPQS6Pdhyv4rZJ7+vAwYY/OrZfGAQJokhe
SnE9Wl/Uzz9ecjE7rCTo73eFE0w6oX0UAepWw5DlrC7fEBN6lpFSjbWme+RJMUzSEpe5Op4gcvNv
P8HKVuBnozAFVlE1YSDodaXoNcNs7sjsUFP3Dut9tVjt0t1y4xzLw+bryZkhhYe1j2arDtth1IBd
ypIVez2EC6qMOUGhYose/L+a77AWj7QC9Aosx1XMU5p2mEsgqRp2QrQxI30e9g8wFl1qHs6TX1pX
dNd31sMLqmbzcL90EI1nxBtq+m1Skdd5M2/2V2igy9I8+0E0Nfgat9rMdat68+opuSBAVlWiair7
41YNhcOMEmixWvWCXmB2yMFdwEst0AqTJdc4T4ABhCreXku0sHnQTQoQAu3MYlVWCTTygyfr5yeB
zjO0Jk8FpSyYWLZNiUEDT+48XC0azKPnd5OVB5J+Acxz5xCl81Gw6QsMeirR63fVpECO7yS1p8SJ
LTavE2Zklagf21C8tBVZ7dq3YeA4UBGwstANqHYe03Bs14S29XYI1C+VoV1oayrck6LsbIkots0b
j/E1uWyb3FcoUlyVQgUCyyKkoJr6Ji3P6cMqPevFqyNEHdmNUfy8gWxXXGXwfhRiKTKo+ee2eONo
EwBTifhFg2uaXs66JRy7es4QH/hsWNFrGP+99HsYFXjH9wLY2Wko+2UbFi3zFs3F8kGPhE7rv5Jx
u/tPqpGIYRkGZsd6PZgIQcrmJjqCU9zq+S4KAWxT6px7nV0hn6gTIIr7OiEYM70EylqHylkb+LE7
14BTQLN0x0T934CDJnMROCJa8vRDCE1rfFlM2vBy2RxucoT2LVCaFE+d55fDp0+bihIynPLRTmAi
mDCzxCyIoWrVBxNZnNYOrNdUMJvLmVMb4C24Yiw0+s90ATt7khUMnrxmjdrLSIb0L3L6SkSLDf3d
SJCU7N/BPphnemIukZABcmlt67cNQayFdCU8XP8pdEwkz5hcDGRzNXrbdJb7synYU9L3RZlCb/0t
su0p6VhpcaeiNjKVLxdcGLyNH2XyGmvBQbQfl5+l+ETX7NT90mEkwCSM3AdrLWYh7eHKydQi/AN0
mfCOHat5OpPG0jRA9dRnjqqIzXofEyy9Rig1FETK7bsbgE9wVUlnamNkylJIlrHprdQ1ssvYuA7I
t8/tRmw0kTcSuol4N7sPhC/JEbSmm4sDzRJ9aEs/TizUk+llAV6OnSvezPr4ZPz32IBxS9USWLF5
/An8EkMC//U/UEKaowoaEB7jBQ3Rx1LL9pnMFYKuoC8IpTU51TxEfoKsdkBJco3KU1fcFTVDbFej
EQfrP4AGo4XD+lNVX4YV10GXiLh4MOl0MLJ1Kvkb6ItbBgSXPN4oOkV78OQNrEtKncNsvJDTq/xs
6ANpnj0rN/eFOXz+fb68kIiKEMWBXhw2PRZxHs69D96OI3byguy6f7p+3p65QnLlUwWWBuIOrMtQ
mdgk7X7/zHqgHHzq1XU1fw7+RQTVDQnjCXdSXyjCmfU7uAnl25nrf1vGrzEP/BymrbM+x4wEqGzn
uIVP1Tk0C+yD1ohI1PK1u4+ypOT7arTFUO3oQFgi1kR73oXxE0svdHFfGT4n6nKi9LTiHQ2Sxw6W
9ZJMYGNm542g7Nn/XXTAw+5xHRGPYHq6zdbEc3VRXA16wKrGfUeULpy6hf1YaQHj7Rgj6M4gQzVH
1aBX8SQncGODWMz4SiZT0DXb2ax3LLkUd2mSwyeP2mMCyGj0HFhQD4R5wV+fvVWwjjWqYnjmshdd
TD/vxOhcG33PpOfJ4AJx+VXQh/JGNDkpBPOWwoZjBO0o/21sOo3QDsaQt5jr51jGQqbKwGgG85A0
wkBYTn91NYMyaLcxoYPaSsRQB+DB5IdChhN8oh3LtyfUnqZ4qC8RrlI6Zbk6G2NcJRMRx+X8dPgl
WehDoqiW+86ZZTnAA6IqTgOopCs2Y7Bc46DSqvA4YBGA7ScQpPhuOCz6BrD+BkmFHr/nWryDwsKX
rhdl/dOs6PK0/7RuEed/VxeWTUZo3ybDjWHLtcYBQY0ozSBhDll39eijjVOdkXyZCNXRZBrHenxl
DZgJp0NB8JvBBWToYHRclimH5wMwnsZ4OmRc5rrosV8KUs+36nkvrORGJgYQGn0QROlFbaYAFdnQ
JhJav+K3xvyXTozZVoO/0/etGqTdAuEJsPirTkfv6/E877vKNa3yJ87oPr6ecUCuK1JMSNj/2l34
OmSOo7QIbnrl8YuKKDJDKwNXgvRa6rNIOmZgL0jVXhFiqU0i8V+Sn0wlVKpRsV8bdowkzRzAd7Q7
xDv3L++Vj8VmTHwR4UeSuDuGGaAEXc53doLBPNsDuKK58qdNqaL692ZpqI/YllrmTdt3GbtLYgnr
IHNgpVBDbMdEE8cSet7/rAuQsAuPILBRzqrn4fsm5y3I0Ice8OwKRLzhZi2+FfZoMnRVl+lvlPaV
lwLpvoA5kr7aKqjuqxBfrWoXcMdyksfurBMGIu8kKwK+zEQHzVeXAxyntG1H3hlNcrb8wAtRYisM
LE1l5e8t28AG4ZUwki0e0Dw5/gj94Om7VMQbwsOgQGDX8qrBRQLhSlDQvEDKpKV1X3OCmy0kpJTu
c1NKL0qHgW6pJvyWleQePeplX41IbDT4/KbnNTpUhLMUpDp0ekJbtjNPUWB5zWFwGxz9Pf4Zo50A
oOriZV6kC7dNxwHmMxb/yGs2iW344PRpWuR0Yq8qwxLfkcPwWgnwsJLBYKjpCsLJt0QkJviEHZyj
9qOoPMrsDQpx5tx/iJLvV6OtDdyjND25x46sbKTYfzV8yPyNNZt4Hsxk8ywgiJysp8mCv1EBSJuD
TfnRoxk3dX8NgjtLClPzC0MudmexuybuQhVE5kYwYRY6vt/JH+hm7wY12oTsJNVqBl2mysDqCX7w
Jn/fHR35RdjfMe1XI3FYcwL/FCesQpuTDei28ks8DqcpNk4P4PwtpLp1nIqFre3YU+em/9afFzqy
Fh+eVlPFZB3HeoFVO6RNphJCHQdOWD+VtHNyt/tfvADW7mei8NW9fIwdSEAHJHk6zsHMwf+rQiDJ
rbzmGFGERfq0V1QoqFzd+snCvfO8aw+ycJgm3B//BBdAk5UHikXS4SPXGN60hFnmVWOi+H7blB3t
vz9qdHoWu7FmMEzcLlAXyU5cW6tDjrL9cFppAAgxNGvzGRo51qgHz+Ho/ay4mZBil6n1I7OozWfv
bcoI0XqlMXlK3QeHm7yLdTJn8GaoxKff8//5F01iIf32ilWGf27+oDjbZX8ZFs6/sCmfCGZaSS2m
/nD4NfTutFl0T8FDC3j7FoT2EbVO4XAZwWO9CpeCvnNkYUOmPy3qb6isvNNj6Fx5xM9/Ck23YPyU
LKQbSmKAs98EHMcsNF6vCgTOwxUvMR4tWJ3Rpbhe6Q/H1XxDrMcCLJ8H1BrmMU0N+V2O6lTtfBjN
r95u925ACobMb0ibplSG5ko4GhZb2qtTEY2YGIowZM6/0JhOkbB5/GZ6hvLa/BN3qfeFqeVavXH+
EFRXCilIL+mfamotK6o8HQJOSXJH2d/nNaPs8hbLdU4A9d2YHRPQpM8kcoqvKNAtxMBTky9gmz6/
cypf/JeFGDH4g0+4yFKM/PJ0fy8CG1dIGPjYaU0u0lO0SjjakXoRnhVAZfPjFp88eS8OK+sJu9tM
c27TYDqRwuoTNofZejGOCnW6/NPvi/uiIZtO8JNdVbM4yZ1RTd2HMfk7QF4iwWCjxyYvMWWyzjV5
9wJ18KjLAhhX9Z7FwAyGP+wJD/T/c5H046qILmX+dngz0Miy2Iwfwd08uMRMEgm5m1oYe5NCHMlU
t/Of5RyPfefSn10GhcWfoub0wh5xyico2FaqFxxVAetknQvm+qPVY147hLWZpp3S70zv+KkxGDv0
jSXNzSKhiMRUDNEosmMV6PE1V2ylehM0BpUtQ7FZOUhL6GVUurzAiOmL8GkAr15C59l10GK88oCc
wv3dBXQln9K55JXJeZGGqVQwilk7YYxMxk3ctUvFOXkVpaOC2pcyP17KxL4gGnCgHF9CWUcVAkgi
EvFJ4vmnJWmh548fd2VYKzh9G8/0UJwceUvoBZuWIjngtEs9EDPYAOrQhhQt6/VKah83fmy3/3DL
wlb29bas5AzTZJlAUxeDLaFN4hGRl780VvnA5iK0hR5+izTKGdlHHj3lLSFE0/ScvTyN4bLLQwnY
9RkZATmAHKm7yiQ/Qr80sZ2AnTPMAAJXBNr+9I1YHpV5yfuMWwcqToj281EJb5ZRRemONG7PfcIn
SZqL1UsI/7/dkaDpD///KSkSy1je6j8MXh3F8dlNXVQR+s/fHwsFHXD71JXbYr9NFjf6qOCtDG+4
BMthy4NROIIkF1vfESycTZpPydJj4/p/xfPhyqBbUZGaISe4qfX45XvEslB07MALmqXOOCEf7ckv
l3p31ekdu0WK+quWxA4gUIbLcBe79gmJBV8yv5dGejyEP2Me52UkD4kXdj4amVkictSuMnnYtiLO
w3nBjWjCpipa4kvsSXEThWyQL1PI4sQxOOf/ZcMlb2dR4zeEPglvvHbtfknkwQqS1DP8MNC2QhJi
VZhI2YCbuyUOYPtWkEu5ec6WgrXkmaapjQdBNZOC4M4j7ESAouziD2AR2wg5ay2Dtw0bAuZ0WIHc
IoOcS1UWRjK3g50wv796I7ykU94cw0SREaAjRAqDxIN+rX9Hb+Yt3TmNwKdHAGIpuh8qa2hmyCB8
9PiUgT2Trcrz/4VFw3mzb/BGKHCuLaah1+xcqAPWSiW9aihyTLEdkEtAPXdsKMJhNlIPLcWQfebN
ZVZoocCOPb5Bx944YKu3+cmh34zSvQtpXrbSCejallDOV1UFaE+z/hnbdT8LHgcSDDLl6Kc2ERQa
C1GWF3TkBOQGYodGOpuIAK+Ch730nJ+F18+mNRDIyzRvQuI7OJwyHEXbM2jON2m0Y5nNlfDyNhvc
4Ji/urCCg0gT1vXQrE+CPP8N1b6JLz5/ts3YOSNXXpoTmgz5l3Y0v4SM3DuReYX/Wl7apoJ9YnV+
thcp6r3gBqLcg5waxGk6thaf4gRICSAxdh49kNC94m4U0tafEHGVXEooiJWjYiISnGB1JERYp3uV
OQSJQzjRQ4gKZzYBPFvcaAGm9kVVlNlpdMDE4g/wKIy2/lhkbFyWKNr0fTzutRkng2pLw1Lca9uv
oFdUS0bpiHsHLPvu7I+6NbKAlf671TnAA3kSiU/h+xAEFgY5zYaZCnrvkVbY8MnG5EUEHtjOuEzM
RzpuMxpf/DLOJJ0XphrF26sH7sDjzOumkFJuK0tzrr0Kh0iUz/9if0F+6OQZYRwSfVjFJW09binj
f6mrn3rnLLd4VprZAsfbVn2c/i0x1CERFygdrKPhuuT6uGNVQfIigmt4zoh9pZhmXdY+LBspxuyf
uASIwi9V3UuSQgHSlK9KK4KU5Tl3Mo1sMJ0ZnYULv81KuETDhjx2Bw71R1pIiVsOf/3CInzgzfUC
9YwPbKxjZbAQqEpOkb14nvbF9StccczDsoTnrvmKOgm6KJqO/vy8qtYvKl2kNsK9DV6yJjO/oKnc
hSCGM59vApDk6d38ACpeo5XBFLNtNwj8jZRhnbkh0Jy1YQU9Amp5FJXSwdcXgrLQiMB6Ryfmq0sW
x0PP7RgO1TOvrX2G/zRHFNR7m0qBozHNyeZQcJfbz9nEYLuk3nyVsfNY8zGQYt8Hh2pofWItNq/1
QIYxcuBB/4vwBs0VbKNsjBSiVrVXhF5MN2ikD+FTQ8cwAgu7cTjCTQePWXI7tWWy2Udo+Lqvunv1
hJv3y+TULA/EFxVE61RH+fRnZ7+8d9J1JS/qZMTtVjuH092gUl9H0qSM2eWdczkN2S3pAlQG0Xuj
/aS9HkU1X6C0n08Wp5W+nN7WCzYn5VzOFs9F9/vkM+C8f4LxB8AZQSw7UyjLrB0KIX5EcnBVcRIS
SdtDY26lKPoZnDl591+I72eJvee+sjqrlupNrT7uV9wKuqCty82o/b4JNQNqVrCVagz3N42GyOq/
SMLkRAYm3FtS2UJjwEtl1am2ALRfc1g/U6IqOydiKSNWtt2Z3pblhdmIlct6zECacBiSg8F5t7/g
mv/HnuQNrzIGQoiqt9ARso0JyDrq/bwouxcFoMdUIOIrxWFzzrQ6JWHAn8zKqfbasj4Z9fdWzMsl
+eufPoe6UvxAIl0fCdRUmtX16/T+4u7OjyNeR+CUHZo60RRiM9izNl4hcFLN1Aniz13DhDLtKsrY
KWlEWKRqxex2YxrtAob8oYSE3xt6wUvz8vyah2/sRZaw719JeyyL99jpJWg89kxQM16vMBnqOOaD
uP8bI5X/XqsPv2O1zw1i1m0MXpp1VV648ztN/g54JxxVcUJ66nl6C0MbHFH4cFQPAe3MFZT6BKrL
geHB52vP43sXA1tRSglG5wTwuJaDPPbFtsUIwscN7NOcUzHg5Ukz3u1Ns5t4+Z985mwGFGgtCjqn
p1xmEa3VII8u/k3pcJiGmN3W3mi5enYNP6pDEp9foutfZC4Cy5j4tKeAq2CIFTgEKRZ3gYemFrl+
UwJo6MbZ86yFDdKjL/T2XG8FE5XDJqjMaklwZT19Xaaj26rgqGtW+eJQzD6Zf++RRpnkKd+DNnMi
ZSVM0B5BpHapFG95cFvgZX6E6JOLXl+Ta9JqUzGmXRngZ5pxer75RE+m1SkpZGBNPk6cbOBg1kpq
Qypys+CjTefMOHIYlQNxIH4NLB57pU71h+6+IHdq6HLxuJ+zg+yp+Us8vBZ3ofnxgzqB4QbQZ/W+
sdNsTiv75o8kpAp1nzb2+CFkC5iqXST5FY3seOZtP6348ATjlfD92xKO6XbpM3Abt/okYfIoMJlg
CSN3gEDQTx8pgzmyfdDVH8kx7Xe1Al/eCtSRfVPHKnM4pZRZnn/Ri4apru0AdDhp4TjQLh2ncViF
jn4LxfWP9kqPAhENQGdPngNnrvkEWJps8yL9dMRne7Vp7WCTSXfSZ8YpjIsFMeQKvOx4TcumU1Yk
uqSLukI/mSCKXpHpoYi6+IIw6UePN26mOeX7ChgE5m6g7esVymTBpXzIqLYk4XtnVCwIM5n25SFN
xTcMbZmQoN9oUX3Baqk+AQnUn/5DfLecK6c7zB4YK38jayxr7zKn9jJakBHt4JZDau2NrcCtiVud
irF6GGO89GO4yGICm9vP15b20aHrFIkxIsmEH6ec6Pn8QOykPv8x5J4Z+t18tXEEePWHwdD6Jyx8
GRPzISxpP9CIOi2SrNFfm0EVofA2nwSWemPeGpWJePWrzd34+KZxZYAdHZfTih2JeY9LJ3IDpI9Q
bNQUj/YGfp8hjit4PKpkpjsG4MNhoRQub5nR8Q2YLoGq0l4hpYvvG25lhgYAx1mZCs6sg2evIWi9
Q6E4QguRDES0jCwmnxCh+QXNjIxfliWglGUpeZjoYHj1xZFHT/wUFO22Fqs/0WYBvbdX8QXxQkFM
8+9buds2raPctGvq/5ygB4r+pEH7h7XCZ9us7MB20Cee1DjVR2wVuuU5hAGP3B9qzQz6mgQMDZrg
0CSG+mtmVT7AP1/UOKFdkTdStRZnmShaFPI3V4C9bUFmCzUF+V4RHgHPyXFsADK4XiWtyOdJkrFq
74YQAB+lWIt+xiSEfvWxJRqA2bfp+OvCZxOmw9d1lZELbKLFbxlofGLf2bLp2ilXAwNtbfUE3QF7
7rLpIpi2xBI2R0Yl26znJSfykgzGuRTtsHcqIbIu4fXL+8yCQQPp4i4OuQZ6EEXDANcFPsdCTTal
7jqbsCY0fKmiU0D7j+6O4BW9T6upzhu2h3nnIr09UlsdNQSWrBLYBjgyoPzKquLs3L1xHCbdqL9V
Nd00UWTtHeL4I48knGmKwEtzAK/xko/hdJeOA6Ss6gWDubw/cy3nrhd5SyO7PZBGDB4y33KIMIMc
bpihoPSV/39PNtpT91JzlEZMnBpHjiwOZyGLi3kPGaTU7WPlFB2gG/vgNcbvTHLhh6sNFtaems21
wn56d0+Qgy6tuxVPnqZQeULIqajtNetR6TsPRCSTjn+y2QOOOnG93jNRoT81BhD5lp1ic6MPnLZN
hCUWSM7Y9Fl2zjVg04RTs0CmHrdK+fdxw0bUulspGMldLeUwBa9XFSHl7vEcip0bDWwsFHCqSbqy
JK9VIOdib9K2AnB2BCIOFonQ5tYC9W4ZPy6RzzcN+xkSDhPnoCWAUeRBF31Qs5bECS4KivNTBzaJ
HAAPudIYK8M0OSaQkh9Uc8eq0t8pR3BJ0NmjKgrSetNXDS9tzLItJM3BYckn8eETmBXYaEirONpq
KdJ2xEHpsCRdboiT56jykv+lUNimcEfC4WEMZ24oaQcmm10k/zB29iAq7H6av4lLBY3gZU59Bglb
EyK+sVVE6oOeB2NVP2n+i4wP+fY4wAIcZyhXppoAJqvB2v4MiQujShrOJRalxCEIF4TN3f5U1hl8
NarRKMCMLHu90+rQZbYdssr4fhpzD1yUbd/UUczBcV1K0GFXvjG5UlbbC2u90yxt8gDuiTOfNhz/
dc3vfbHli8FiCISQlUhSghJ0qawEu+qaVuNsbmQ4mcVbCEfpwnH/gjEBX5fKWMUvQRPZfSSr2ire
d6CUw8zQH6jRus80kIFsW1nhHrx7CIZuvOdRkYP2ulFEyADSOjhHLtO+BAiK87idSsTGJVHgyKGu
mmv00Zyt2duaiB2Du2EBcIVbr5yqqhUUuK3ISn3A5jcXgAUCysntmGGiVs3DJ6ARVxAAPB+1UMeu
Tbf2GdUGcgZvGjwDBsjTzRENWFMG7rpEuirp1yNIs/x6nXOdUP6XLW03Q91kDIzVzW6F/2D2Thie
cf4vLoYnAnfoLNtITjBKZ/bSkUZIIfJVf0ol8e70gX3/lY8xeX9MwnLufUy+r6YR+7F/H0bViGSs
f+b6yJYkIo5YHscm3HfgRemBXhQVaPncjtPuPl+10mdMw6j0+O3wjQAIOCqFFGTVxqD9FAzGg0RL
BiADZkItyRpa0cvz0oxgXjSLY0LlU18NGZ9ttBAYYXF7snS61vWV3s/JzojCtWYfGo9YWa7P+2Hb
hxQbZ9luE/ZyaVI7n5tjsHqO4nx1Oh5BpBi6ZREsswGSEARrzPs6VC0dxAMoj+WeYsFXLrsjNQ95
n2RlvdhyBwvH6glnowpDAJ1OhiylCQFy/nizwYEGwu01YZOs+uQV7Ewjfopi947+S9LTYs2FdqKt
cRFNupqimENdd9kI3A6sN1xptv2OM2XKEhEHXfNkxiBqU1PKpWSisCIR2YYcZKDUVA5E6NwAu1Hk
oCU0ruwhlQG5njfDAxPyTSlrWl1bn9FbgKoUSvsJzZ3OYy5FYZB8GQyZiFuhbaZGQs/c/fcf9vX5
ayXvka2KHz5eP1On48HiOhHSnKob5NzFxQUtEMoPisA+MMd/erj6DHOq2WJ1XdXil25GH6eX5sXf
Fm3gJorXf0U6gBGhqpGpXjLGh128ALZsem/e4tRBNWfSNv+Tt15p/QzcKi9dbR8f1Y4B1Q1Pq1c6
5SeUPp1OBQcqjfwhE781QyMakbJxTQZFx3vqeuxDG/RKNmUUyq3XpD16HAyeG/maqxcx5CJO1EIu
lQ3KKx9GI/59IX3bdyBwTF6UotKgfhWj1QK6PpKe1fKkonSvHaLW9wfwCP+jBzaV1LCiapk8L21o
7Y5E1Et8xknXtppWpf0xY0dbBuuc7rJukAMfUuyYhStJ0+JFDCleK28ZSleKZnO2MSOvN7ktqy7S
13AEegcaOQEkU9RV45CzKjflgODURpCJ1bTsN1Zjrq7zovR3e3v27uDGz7F9wS1zSVsArLXaD0Ci
5xxZ0xpATU/tyJioOPpXWAEzG3p6bd7jl432iDD73zOWQi1Q0OIjMstBQMAiHCBo/NtbeL/HxgdO
PlYHmz1lHePNo/yv6uJjRMcVEsZjM88M2QZxZiech2SaHtyhVGhzQYsGSE+tBDyOksw/OPH0oimD
unTVSS2aj0e7xVrdKfjMTwVL5WXK7QdTbcQK2SNELi2eFWrm+SVr0ULvDvWkxEttGz5TDTBUxV5C
yssXeYS3IBMN/KK+HwqAI+R0ficulRdmz4CrOcdvtewOm5sh+ZFhPKWvStyB3z7O9w1gIjkmhhNf
C76YitT61CGFRZO/gmQagBl5FkR9kuG7D69KzjTPT548RDjh4v/cuuM4J7V2J/yfB2xnyvh0nehO
kYhCLz/PGMaElJhO+ZM/6dvJNpb3HWHmkhXnmO7yNZw01jABq+vKyy9XJQLMzKDCaXMMLrKX6Ndb
Lc2SpB2qSLtizyOhXA87ZX7cymq+XY6CYpbV2B0/RSLCxSG+epbwIY4Bia7Ui8t5jtKouhdVO8lY
BsBq3+ZOrVW3z95kgDX+6uweDspSCoKqmtheyWIXfdf3gQ2zbFCgMcIyybrK5VOkcDara2aZA3IP
dBOAhXogpHO1LISU+oFooyA38aEU/5oItTlWligtljA34JohC0bw4cR7kcLhmX5KBE26jOJtYPA5
BqWdmsHDbO2DXFlC7vA9voENvZysVRJP3/QP4shuWVFdJvhfZMQ1NzWJ3FgbDvThWmwVjQBvg0MJ
6ahlFeXgcMKiREc+F5jT6gHCfIRGcdcD+MBC4SGS5MXQ3btImRixs9/nQX5JTWhPFIqawazcsxAM
vFMfvj/htAhSdfEqG0q8D1xgnJfDSmB5CuJlAb8TinGnOAR7IDgIR4z2H24Y1st2RERJfOwdYw5e
O+tiOqh4TdlsJUpHjwg63vmpzhPGN5KN9LuWyFRCuvsVOe6t6hji1JTwCfEyOQfvy1hNuHimr9FZ
6CYH382872rNi19EwCk3zid19YsumVb39judqxWE6cxJ6xpTG4LrjN85HqqvpdtglOTz8MNwnnaP
d2H98ls2mUnY+VE+gTA3Vj6UQzVVR6Tcu36tovrG47mnZT7CT6L9fcGO51a0gymHrG93JrJxkKlK
nxy+CivmIzeFOs/gzRdMv7fENP7dxKYhgzFzYz48j6OgSbzQEEmlviIHTLtEPGm0kMTw2T948xtB
v7h+PocKSU4u/d3nFd8eiwCyXP3vb72XZWsxuaqevnqaHJssrIzKwPe7vHOi+YlRTWQG42YmEwxF
zuJf8PcG3Bf8k4N1VObn/AvkEd4suyrq0vh8JsdFWuM/8oxQcfa9sTQ2mzskcAlQVTGfDdai+NBB
be/AGdQ/cGcg/nxViNRl0Fr09un7SsfHE8YZTLoQO7FsDFMbN4HUzqOmZxXaUe3jO94+SZ1I1nkO
Xiz2rAfizDvg4kvlNVx7nr1/dVFky9CFOODMwHPmfVmbwxzvv5q6T8Z/8FLSMqcuWX6Kv3U0HEQf
DOmb4UJwctt0b8haDm9LSCG6weS4xw4YshIp6hlCfooi/kv3/eD/1GzbOaMvOEk0ymYq8ixjTGrc
hDA5nSrAwBdi8ripMYZmyQi2gUsSIEUDbHkb3og+j7tG7IDMQ5t1sNMyGGnGA5FRH+r+wcnuc0uM
BhHP3rKPZk323s6bBoscOO3dtIktyxGCC7u2mIQ8Ox3a4VLutzVZV10K+MQ40/dtt0P3dcly1rjL
rP50T78dcbgtdgo4THelIqU0X156dou4BEBt2OGV+LaSnTVS301abYLYcJNVwrgQ2mj5lKvSsUOo
A+VgTZMvrDAeFhUObiZAgphnx84/wlu/2UNAqxBh0rTgdtHbsqgKMfCwZvXQNXib/eKsJTkYqS8g
nejHpIi3wFsc9eJVjMvQWMNg0+TDoPT+Sc0xbV+j6VP8E9WYYCGXCmgrp4WnAW1a0KbTwMh+wVzI
yDoGqWGjR6mNB90tH9Tqnmv13/z+F8zESEFvbhJj/P+7Bkj2o+HomICfM2r6RrppR8GCEeu4KHqD
p9NbldLL03+JhYIATlBy4oGgsSQq/CQRkT9+KLLFCWj/yWmUXx1HfmifPS/2Gjc8DdQgfo5u57vx
LTjkZmdDYTyJfXDntLaOeyDRP5hl0BZgKfibBJUNLpbboOdnDwnOMSSTN3Zk4MFg+cM3a/6O/G6V
Li+1kGzqmLBO0d02yDidcW7glWmvwxqGA9wXBl9N1pfIxb9I8hGjbOOkQi7WYRB4KIJ1DNLZ3R/t
19kNRw8IXGN1PXgyLuV12oN/hgUogbJOdOjbpPMVboWilKGZrGmEP5HjEFPhQQiUxi1URo4cKoqC
UKgY6lbETUH3z/mn1DdRj0EviNSfXMJrgv14rQHdYIiRb0s1DspDscwGUJ51qCii9xIiBZ+VT2X1
tZm8sHOOronse7dPTtbBHNs7F7/pxmI2hJJ1nd0AmtWqvPua6aEvbVMFOfzM98rKbQvU+rOwYTvr
zio33i7PWmBowCV5YUINAa2iG31XV8oWyfpFpQgvTM3MdsbG6QbazEtyLaujGqQiSBHDQJqHcScd
48Fq4Cl9bWYbMxKQpZgdr4gCK/UVUiN5t93RSoMB4nYgINswqfNrSSiKyZLDwfGO3MXuP7VAfecF
BCVnFvijVHa37s53op+XeYgubPO/E45TH55YlTLk4QJsAtTnhRrvjpdopc40uiwVVB5tgLsrtk8c
AboDp1UtiZwNKC9jO0ofZkB4u922iSsm20cNYE4ayQg9upMW6xYhQc+ev29NWhYszevxbZFsgAse
ArtUMwHOOBLR+rDq0GvSkdKgwNt8SbPwUUFNQSkc9ik+BJ+rx19hHTCtyDIWdhjvFFkJDur6Z0GL
mZJvoX3Y+wymLgSJyeGEhpe04pKpgoA+eE3P3HRMWnG4zHqSryBq6qHsBknqPcx3BkJQtKNkeYZp
c/BeikTkOHatqp4QsbuifSzYlrESrRv9LrlP3AwZ625GQhnlAfisoa9+BPUiOeEHVuzHrK9PUZWI
pv1U+3ldq2K/sW5w0I6dYjGgbcGORnv3kQvtvoWfJUoZETTd1Z7LuAR1MPpXMrHcOxv/GmzF8TVa
zD75k4eF43wbV3iXOB1lR58sA2N21839FQmnA676nJ2oTDM/mDeCIEORaDRlj/EB+1x7vydN4jSq
TFDi0le0VCHHiGuD3Ch84h6q755WYumYgPCyrQyv+9ooIsWzLukf2JSBH/Q8nBsVQ0klAcpyd6ix
nyvJ0Uz3CJcj9sC4e0sJDQGdQIJK6OBgmz9o3gktJXbmAjt/0zvTXdbW3VYEj0VtiiywM/fim1IE
+xj9Zy/uVvMRTb+O9BgWoyW/0wZjD2Kk6vLWZXjVWBirqhXSLzlQ4CCu7vhUXQDPpp9I7W4kRTF8
LV63pfzXyjJG4UACMGO4AoGCa5gcCYI2Vu02Ji+y/w4KosWNKqM3zOUB99uwUBwfMqnKuYKnwFos
9GAAkuVi72Ynpet/pa3WeGzIkxr9DbU2vF1KYbv4yCPLQc5au8Rr6G5KFQrdUyKbUQX8DKv8AGEs
wYDZSIkGYTyhA/GQfyXnhLzujkR7g5T3E/koLSTVcdwTMKvIRn+iqgCStJ0Th2pLKiX30Aav8RqG
L6aq558IG00ichVIMNYKSpGbzmJ4hJTj4pla+K1PhMvWh4uLa2L8pugT1ddtTmM2ISkOoqKCaMFj
jgOY0AYF7Q3CeVNpk0sFRpYNMnd2qLAdInHbe6PCFkqxfBA+BOmZ6/dH7lffnqc8hKgmUDzjlMxN
A4vMIAKxZacM3RUZh6TzIPDXKSRXC0s0brA1J3U++xCJtT8ILyH+X3NBZ0E9Vcgdqmrg3/c4JGTy
7SZ2VoBXdZQHFVvFkkbsywm9ZxSQCm0aIzfpIGDDs44ktTfhGG6YPR2wfuUW5vnXkMWnUJwuZurq
JyrlA+lAiIY9Ejp1R/dp22aPyL32MN4UR1DkcG7ILi77c80w9Nu8LKnLaxSOCsJzlYHXzo4LqPnm
IMNU5yyn7q4E85vbWc2x+xisPvz2vwB2PPDJV1hgMnG6EbtoL1aapoF3VHyK9CfZGR5ydkWNEIWs
sl9DKYfoP89+YqPqnkFBMzNy/XJKykUnoCg6boRGlLyvyhnxhzld6j7OWmeo9JZS8jvrjLw7Yn1X
geeG0m+omgqwiP8XtZOf04W627kJBfT4j7C3Im12UzF50zhxOHuTKt+HR9+slpvZY8ZYlkPSMrbD
boo8g0rmcNCgqMqIIoWd/SnB957Jhx77Allbh5xi7G7Pfz4xO6/UIBjDOfm3UfcjmiMky916tDbr
/JsUL6OHJ2Dqc0hMEAsK/yLaSPP8m3M+wl2Ne8a2AFw12kw2OusoecZB0NUUcUjWu2o4hjOyO9wB
dDe+XOIMmDXUqvokNp21gxGNlF6FPfOH4RT+V0LLePtRnarKZi4MV5bL5C+6+GlC/I3ur2GL6Viv
0E4o6YNIENdJTIsboIRUtDkYGKUZgrZZe5VyfEg4pk6tJ0IkDO2Q1vQhqEtNO7+SHtW+fGUVoOhL
XHnDNTfcbZgWQcTrPs77K1vZs+pAwWb+gyr8im4prFn5ApN9BDNzqSyKwpFQhieU21ewh1Zrkv/k
CVMfosmnoKkLlbDtRIETgPTnOuX8crlRGIwzRmFw8zwR2HzcnMsWm+S6A5E6qPNxv0MDrB0HnkV4
0FgZwJDpac0+fCI6HTqR4XlSiDOZinMhS2FqwYglFUPspG6IhQ5vm8wobhFbPquJS/YIX/qkCHjL
zn3vDeiiSQ7CBoXcI4y5PdpjWzThYE+HNXj8NsLth0G9SBQqs8rp3gZvkOE34K/zSg7Yz/27ySXn
6WPV7oxKbN4DG1oUwbZ1Z+j24u9RwaL3kNWY4R3gw13mZwQo3ylGDqwImU1kKmhXEnAqsvsK1X92
8wehmjW2hr4TMsIe42kUz3LhCjqmr519EG5Q3rtCjDF0bSRg6RHVOlZaaRLXk4cA9uhuhL2+iw6l
tarQYh8Z8KIJPw+Xqs7Z8sdMcmftCaiwGeuKP0LLacdQuQ22YXknYUSdQgVfhbvQggEXyJxC9K3i
XeN9GpXpXSqY01YQ2ISj8g00gHIEHAnrAaE5w/cPvsyrCGTZy/81GM/xXZkOkuMqplgRBTAwS+DY
wP5kpVYOh9BlNFqDYDI0tvCBKuzRGYd6OhRgMSn/4rY8ysT754dTUg7NO+IK9SHgLJNakxJW6UDM
EiuSzFAzzebPHim9Sgap34d17TCJVp5YE5o1EBR0vG+HuZazvncPR1OyGCkp8KXE9MhKm7vpbfJz
mf2hyZZB9UAXduTzd7lJ7EVrHy8ddn7PnmQ2MSxwq2XoZdtGM2OW/bl0HDPRKyB89T2Ntjal9AEM
fftqK/QZNyoovq7CerWVb63GUpGbvZfxMP+jLcpk+yuUrjNfjtfsNefGbLH1baa0zm6Esc8U92qb
4ctYZLV01y0R1amHIR40C9nMfvDPRetNRVLpokgIYmGvNwD4Ef69inepx+PG7lPc7kiI2s7lioR+
5ocsnCHvFNRY56rCTyGckTyia0tLJJTnR+JIL/C08L14Ruob9odgThAO/yKOkvYSSIr8EzbJsQxi
wmycVNd4FbFVcFPSBNvO87+kVldChew12NsXPf7K3crG1W3m05Q2EJwOMkVK8Bv3m5aJ8ivalZpB
/9vPkZ8CT5NKKAB1xUoum9B0DJiSVYKtkNLjGHx11B14v8OOsujzugP75uHmQh42XwxR60Q1cHOz
iJFPK3NSX/h39WDjsrPLusUJaqH01Q16iJtfS7JaJtZH0cJ1wwtQhryBhaNAERjDNQOZlbUPLvJa
iG1td6H1Zzu7FFX3Ss3TzdsVJum110E1fTQdiaB0bYlQIj0lmEMJ58JK8Jb4smZCcLM2M5eClZSK
c8LsoSahzCyAGIC4qAQSQtjrezZreH5iPlz2mqDxkAC6hvTYab9tem8Shb3Ubh9fvraGs5RvGbN9
fh9+tG55cjEJIR2lR22CmtaI/oaRdkvSQUpHoYUXoyPu5mGSmmOMvpJm9NO/9jQQqBPVyW4GUyjX
bpoX8ZBatQbKbWBfxFmz/m/o5HMkE68BjsKDFe/wejKsEacG8kaVzhKjjVpdaXyyBN5+NmOLKjAw
H1IUTRPkhfvxRcn9dHZpYAMA+BspE2LzZUv1wyvx4EEcKQIksQhU8jSTrD9u20UmJPBZidOETvLK
vg+INx+YMDMhwC+86uNHWgpAOHkWr00ParG7PclWDeiUKbQvMAqQ+Afxi9GOtf76X94nJmNljq/T
qjeh57QZzy022+JoPULCMu3tlvFrcbn2EdO51uR5odBjHB0Qic8ZdIbZPTwky3YjXvSnq52tKNRr
LzHuxnG/gnsJRDcmTsKhYqkl93lxRUWK+dgzXimtXUf6dIJnePdlFejlE45TO5YmEnvl4+LX7qjf
3YDBiAMr1x7tVbMkBbOEkp6pF7H/ZIWNNQRcrMNpFfgZcNH5/kspak+rp+0FOP+xEhI02fZ9i6eW
/G6ohfBu8bg4ZizeX3MC/16gjDnQibsf/6163HfQuHxULvA+WHECAKG7FH6aNXe9tQx0NviDGSTW
lXrVBjzTstgfBRbvQupLSIXPQbH98QaeTRBrqgDAKV9f3Euqv7DUgjgNyXb2IaJu1vA/fmA1pIYK
XWoLnXbVw0cZA69PqiQD+O5BFIspGDOWOMmbFmZGw4LM3pJDLuUutRgRH+qPMqGeQKFpGhG41DfI
RFz9BloaMraiizraZmNKC76NXNlhzWsM1Qkvl+7eOrsovXvuZ1VOcC5p5TqDdw8/Gb6QWGgl/ZIJ
/DNpVeudCs34Jcem7KCSz6qSxeXyhQXMmxzAFaLxcOmFIi+ZHGaib4ze1UCbCucgO9+8HL+HI0/w
vgABUi6i8NiPsCVqVv/gYoCSjSGrywI5lUJmR8jTcE0gL3H54gvImWrJc4fL3sJ6L7G3mt6V4rGt
x61kvFAYiFi1MzHu7TCtzCD9cfcdfDCl+nXuFflZpK/HGhaZ9z0X/5GEs9ngXiw8/6bLSlo2v7B8
DR/RaLdJd5tAsZRhgc4mPEjxegjPdU86YPMwzMOkdgiZ2mKS+c5wCGKKKtiZCxDpHWATru6soKEM
uK65ZUzcT6fvjDToC7p34DIuwGsYdAsbA/kVVVLNKNpMIA29r5DaYgWmXxlWN0PoOediDopSNuJ2
QxbXjpGSl/2QjOFKG3wDYwJMU37mTA3x74TwwpvlMEVO0TDJkqtyYlpgxgY+X2eG0FTkdf/G1zyi
5tKZHBdfaTRr4hU8Ux09qAjGZlpIKNpN2HZJ5PcUYyz4I5wFtlkUfO2KTGaiv8/Ywc80ZaME17DK
i8vmcPRxAOV/b2/erU5LqQdIbBLXST6JIGhDo55MktLnBs9q/Zyc+GZv65qcNy6JbYzKaUDYzCjU
+WOmi3ISPQPC2xWdaJePjItaMrOeR9IWK/FTIsMKljWm14KaCs+vuvbUqhizEJRl91V7DjDrxR9Y
+haI6uaX4LlcR+6Lq1P1/2v3qctfxx0gVRGi7UCLb8TvMYblduhbf80mkE2rSXZmxF+6jvSSQvW7
/FtVjjyAVtHGAQVzc3IQjkeyPW1b2Rl5M1B2QfZso/GuXvq1mi0MdOM0Jb6m8DpumUlpO3LSda76
efkFAZCQEgg3dVaoiQ8NPF9jijCLR+0YO7Wy+n2n35o47VmzQFh14P3/HK4U3OnDQS9tpOe0wXnK
d4c+ZB7T4iqAzINOpT6bjTxLFJ/lc7u0T5MkxUmmG76UPLIa+EBwD0Nu15r5gjLNCYXrASbjSIW7
ZWtr1nHjAGNO6fgE45isZO7MnIRFDOpg090KWT+Bu3IeG7ygP32jzvtPVM+NmHyANBKdP6NQWAjE
SUEUxo5kYAtEx+6L0IMikbgbVd0prBbwY1yBr8+LK7C8z2UCaMG8WmcHdrK32qO9+gc1dEOrVTms
9EdDgaxgwg0T5a7/rWz/pNxmrIHKQpp4TuZv86S5rEg+EZncFJ/N/bd51Ubj0eKP+PI+nVKTUScc
CI3HIhFenQfAHay4xAOcRmdqnYgUtSgR3TiHfu1N3CwSQqJDSmB3y711Ri9GwU+CxSJTwH2MTtzE
NJawIdLZCbWoGeDLqFmDCAFKY0AZ/WUeKbYyoVO35bGfi63+GaMlWe/eExZJlvUKPARmDW34gmay
t+VptKzzQwZKsfC919OhfBMrWyVf08KyfKHDvw33aD0nQriWkkh4gm79EJx7orGAz9dLmpNqSR7I
hwsf6LiswQmCPlJ+Lsfn/oUW4HC+gNPViTD52xr2Yz7h3fr+YrU+QFG6A3LtWyDpCWwOvPy+zpS6
vTPY3rV1WfevkLOHHqJCoIL4FrcC05YAOZcA/4q6NjTwQC6PM06XUs00dpW9BUc+XIcubRufAXv8
r0nrzYy4+5Gxy+Qc+T9ghbheFiWOVI56kO+5ZpM045IvjiH9gwLOOs1OIPazN7l+K7gwTqZ5+G/y
nG2d9opJPDpdYtkdLySxpW08uIkNIgKBOkYYiwhPh1j2vzIyygo+XxwoYvoK4mhcszvRWL2X1UbI
sfX7Kg2cFkPoxau81oXOl5CBrnI+ZJvQD8DQnFaoQnyDj051taBYeLShAIzE2Maz1Q818ocJ3MHQ
Wylh6fSj6rNV4V9dNZ/smKDD2B74ckulw3/x9zNjzB0g7L2yEBHWGo0heKcui0XNTHKEfFM+gusj
uLd+nARPJOS/Nf5Bn2618RoFsebTb63ErNYPJxfgDUXb9q5TffCXLAt0i4ijYg+zHHqOrBNhtFZM
9pOgFq9F/rQrzojDv8SMyLphiO7viuBC+1u/vZnqF5b9HPwRm93mLA/z2PRvdsCiXVtTbQ03w2ay
1StuRF29Vt/7bjnKR7hetK5o419AsIDNWnqpaZHXbBIzdzXRye51PeqIKTunjr1fYdRjcpR7vzFn
1kUUgKj11tmiIDS0rWv8DW+uikxj/VGcewA0guJD6i347hZu2oj8DaXv87E3SKXF/vAWqJhDZnk/
pIK4ye0kePmsmLLa1xVTjGo6H1kshrQ5yWUDCEFaXsFCsNEFdIF9P1VQJ52YIEirAkEySeEgM5sq
0SnSxa/AwIn7tAj5Nj/7qdfdtSWhbG1t5nTDsgjJhNa2kW1EH7A4kZvOMpDDWt3AFeVzXvOjHhjE
af11myZCd2r5vu+4c7+MgIcwWaB4xUq98AhRmiHeWrz68bn+zdNmhR5t8sv5UTHDEhavvfGzw+oI
F5P99+NoVetrLPGPmZjjSj4+hypy2FRu7fOEWH1Ra0CsojzVes33o15H3wiPEWl9ZWytWkI1tVFv
kZ/pWyz3ghfOEuouKjud4A0Q2LUCxbYtiHx+sXg9ojhIw+KXyp/H0mGG9/o+bw8ovB+opUVPiSoD
+5PJYLTKURVGfJGgCKt+R5tmw9O3JWZi01D/gHv/u5l4zR7iYh06SUi28NDibXDXp6bxYpCfivAw
AQ2Rd4ktZ1bIv/VJYk1LjvGprI8NC4Kc95DnOTU1GvsBcfsn7LU7Gp1HP37Rf0Y8+nGy5OulYDLA
wFKh1S5GTwJergzN/xaOBK7WBG/n1Nwwswt71AO6WhBXdgD+t4oAd8cu+FCkL8rUzpkMMnJx9aZz
bNyKfkQTeYyqt0XkYB96h7OD2crIzz2U1vrReuD0yz7EEXbHdpkgCZjOGPMy/F4KZqBAtrZRDWfp
fe37AShhkucfFXIrzQEOWdaxQO98xj/TyRa3+Wx3rKeUGS8ULU4xfI2HeyzpZCcfw5ZT0s7lDfei
bTUNxWQbltRGUF4eFy/0q0xJt/vn0FH5h6gR1T9N0BezQbwe5Eed7ULqG1o3AfgSp3/RdCpGsXZX
UMvmPHQClQA2R1GzF3lxScZblelSpHCtda2ZqvaQArlo+Em4XSChXjeWsWhzuY8zUAFvmnpMq7Ce
8TCBUAwS3toIxuDfw2HkM1I9Mhf8ZBahAgKt/2nznQa42a4H9/RK+AFTYxjH6lJDP8MGZd3Z/ZFQ
Q94duFvk2rxYc+d36fFcDTIgyBSdnbz7U7yBd5B/nOCs35dNnLE3k3LaJEYU1uOscZCJQCPrs+vQ
yNrzdBd8Z+ih9wYeZtCjug5/QFO5K6xT7njwuDSVy4wG9o3QFsjQoOG4skvTLOlfvUpzDjfae33L
VTZ70LdEDv8qYjRyS1mDw7K0Ms8KutgnhJKdIMZaz8YnvVn6556jsbholirRRPXMCYwU1h1hnM5t
tMGwW5sNaFyObf+Ok4rtOUkOsO15zwYcsxWgLfdl3jiRC3nQ9DEwhnrqqh1cifbuxLW9ecotUXGT
nkVpHt8l1+qAvF+fdW9jnlURptcqf16e9HXWD8CKcT0kUBJzmvI4LT5KTltnHZ5UDKI1LOL2WAg0
kCZ7D2sj9RsGyFMhq9hLqXKYcKngbnAa618KivcFnsn/BjfmOJkKXd4EpinFGGalR/8O++IQu7oY
8LmHE7cnK28mOSNR5Le17D15tVoV6mFW1QjeQ9eVEMaBZPp7ZHvOrrYdsR6bJkZYD/JDV1sN7ro1
n1dzoSGaQudC4YMvUjiFoh82UDEKODNUSC1UCE0qGeuSCt0X5HM1qciAjVYngJ8pBwtPwJ09xQRC
oDQjpJLQ7PeEs5BAFVSpm/2nYQTXSoO9h975IlIditXhcj+ybKJ2eueMNWV/6b7JgIsY5Hh3DPuG
upE2FtlcE2Ae2grnHsxB8AXHlaXQAgmpG3t6YB8xUBT+DHjL4eyGm9aiLhLriPRkVXVQPxfmL7b9
JDBliEeqAsaQ6CWFvR6B6Edh43/TV5ZnxBMfeOBFsM87EV1L0R9Moq8y93QHarGp+Xc++W9PnPrG
WRTP+sttaG2atT6DxfGAdz3PxUv2gqVBHmz5BJo+g/82WbrGVcnGMF41tCci1VoCR3MX/bRMfPzH
bShZDTtpKsWx1SBbY+YAPBlow3k2zNqNmsbGJd9NBD4aeZXqB+j+AYSeHNAa/YGXlOrgkiUGCy34
suBQUg4qU4Tk+TPrXEtfDmzGdiwbLFnDvdB479ZAvrGJuLM/r6/JjOgWiXNQKplRQ3LzCWw4S5tj
K9Q5J1yCIyrTlclEWCNU4qvgBhlgbSX/5A+WxvP6psitxdDlCq9dUZPT3KtO2hJveuk9tkE35590
VIz6hZnSvuNR9+NcRPzY+NqSP6Zt5TZYdjeOdXWikFrbNI2n7C2SRmFF9SNRKSAvjT1gztu/nNoP
j+NRPTveje5oRiXmV0/LhRxqsNbo75bYDKxrrTlrw5kfz3SISKu/BMJK3ugPvO1I0R1j4fHukxca
pxkR4CB+vESzo6vj6SXTuiET1QS/UgSRaKiyKxKMJTxDcJUDyhp2dPWAcvlMiE8Qv0GBSy4ZEo8/
HVRMbQOw4mfqG8+GEqrGvf5pVGxCEqVLImSxib+atEv/zK6rzRhDt92ZKit614JDctkBoB81CsZz
rrtyFC/nfF0MgxSvgYPPiVz9PpyVyUVtWYSSB6L5jNI8bs7YwaWJsMFiyLvtF/Qn8wj8BP9+OCnc
0cY/cbqf3iDGxUvRKElJnuMVQOs2tG/ZpzBgHMfekmi0Gm+z/cSjwUE5KU2R9Jel3GIiAKa+D1bJ
kjhVeHlox0ce1Iq2oC6hnQzQNU6x+oHWALdGkxsP70Bp1b5HF/9fEmp28kC+7p677WyR8649joR1
I8N5HMqJ6LrjJO+oSna9o3kML0vKjqjQsI/5qsp8Fcu8E8/xAiuAt04Hsw9SXFwgxiZzemVU23ZD
PA6ef7mHYTdy6WouSi2PxIAYqjV8ugvUMkYb8y6xNkvn5AxMgqs+mEXzu18c+zWlnfG/bpkjXh+T
Wea+50O2EVhLfkhpPvELS28asv1FMLmgsTpHvgroA35vBervnWB2d6JxYT7y2CC0P/TNDWmEzlzv
JBu8tIytQGFTjeOaUFMZIb9SGSqIX7cXP5oQ+MKdBdl9PWIR5GaePmzr45F4l2SYNL+yC2jcWH3P
gc1Jpxw5U+94IVwWuQQAxtb1/ZNtPJH9LIQ1CY3yAAAch7u1mo9MEm+Ffk7QzrviOHh6zJe0zB/R
YjGYYLT4dDfM25yDd+2x4nxKGG91BKWppZFXb3MmscmLtTxlo1gdAjAa31koh8lq4Rmj0saYkYnT
SClOeFli0fonqv6nSuwOjr+c1i2E3mIge0J88IjTYPXWi4JnevX7Xht4PVE0Pbs9P1w1MdtWpSvY
2hZWmpC/SQHPkTq8K8y4zxMHhxU54dFTY1CLXWvBqmg/GL0lB78EoyAqCoYMSebtTEewvJWqdCKh
uMmaVeq+rL4ZPdkZDGobFTm0qYLWIj+42KgioCUO64tlMsdw4PeKNqlnAHi+D5y5/Lk/bkSeYruC
NyvO9Ewo4j0VHuMOeiLnMERbioPPvlcBf4CxRdDA2HPYZHEUTSLV0aRXqZNEBuqfwalYJQiXlSfE
5JOOm/yRqx+OYlnn70nHCBvnJtHpTHAx+tFGCNXmxlDTP81AfFyS+SC489ejIPbr3rtwtgsAdQpK
RParNZ8HHja33zcvDXRFsW2Tq8i99TupTkIa2awBV3xThEJSreRTU7TqjwlecEb0uUUlnFSH0IZH
ejtTzkdx/N4pD9QRGscA5g9oj36nlcPz9P7a8sQBcHMfLNt1cQijsggrq/r57fEHgx4unf/Ziltc
vIstfNFmCFf1k73z3OxxRGUB0+9cVp0kMZgVmhB63HMsPUss0zxslqkaM4rqUia+zBhi+Lq70yan
uTQhAUsyldLdbwviwcUG85wH47lc0Ctdp4bWiEmZoD9zS4EY2iDzgMRT4jcufpOZBca+BibuyuVI
11z/exffB6O41TrnaZhOfsanOroPDid6zJtBDn3I3iyVQ1h63CN+v8wYPWmuj4kzUiioZIuyAX1s
tE02H3sLPVHq+e5DaBSPwco5YBo0WcLuOPI8kZXLGYiUWbsXZAwHvDTpinxt8rG5gh+96NoRGlxw
dy1A0TBs7ssQFWVP1EjFTNJIdBrJb4RNBBtUGI5SDzLCp+jDodqels7WoW6g8QqdGJ0zQ5ITO5DP
6VMLxSMVOKoxtH7gKMs+WsRlCEf1rjgLJXkJAzbMkLJApzRNWJCBSagEDYvoKOc5nfaNmr1i5jlB
n+E5Afnituo0jpaEJk44mk4yXWVnhxLtRiYPO2Zy3wX+ExNIgSjj+dbSq1Mij1EQqa9ihLNZ0zGT
9YImbabqaKjB7d/P1DA6BB9JJR2VxWXF9S4FE4QUDBRuvX5vOKzdtb5A3aRO6C4iqr3dRbeFPS6p
sbaBmHK+DqyOoIb6wgS4TPpz48cikE1PBkmHMyDRQlU5u1G3+JZGv6bAOSE1Cu7abgNP5QwfVUm+
xRQLN772IoWHRHJj8Q46HNxtdMhyWewJFpchNbV+aadKX6EYijk1+MfrTsoA11FAcJp7t2MB5/qQ
Xz3ZOhC1/cC9xGk+zhpkkSo4RDEFP3MkY5mn2QzLTK1KRI7WR9p7wJGuqzGoEDeRiyxKvm0dRJBj
h0O4T6rw08t9H/olZY6IrcFWOwbzG+j5wb7tJX6YW6vH0yspstItzAjCarB5O8RBkTWWgRN+C4Ct
SSRQReIoruqisUThnCJD0rdJva5xr4sPLd7cSmGNq3XYerRJaeKGU//LAmFzgjGPabQvlJyxrOP0
E3+xSio4yZcDHbbzHMnau7SjsN3Kaa5Y5RAE2rBFUcyJNeEaQwtIWEGMlGZfzDwYpDt371xvgfav
kqB+gJN/+WvjWbWp/3y0PqD+Xgr9tD0CxV22HQ6UZPc+L3Bz1pq0R24U5lECtaRlXzhX2feRX+kj
4LW89ck4FYE7URc7FLFQcQeW0GVjVKXhQizTDCiKF5iXBnH5MR2LqdcMk0rNgjQhGH4NU4+Sf7kY
B7bQQpYua/Ut+LpDAlDma8kHW9Tmq4ruwniEC2RipoQfVhPVW9Q/vY1THYlPTk3rk/x+RoMBsVy+
OH2Drrqggj8tIroz/Hcpf3LAMrUjOYKOj5jufP2p0p/l0Epp4m/HLBkUr5bDRAe6xYHJo6T8K5bD
Ang7coEMywBbbzO6pNw8IFvA/7jxu0t0MG7h5gRXBbWWD9r1AOUe6m+BEG2dnOocgdYe8+blihLL
tnbnwTwHO/RKUCl3LPN50eZBthgUsmgvmI/23lV4or0Mb1GQqFBTmP6MdVIIgI6f0MCfQr+S4Vqv
kHXwtEMfbB1Mf9ut53230hQXv3u9Mnjs9hQV37WH2LP0PnNHV4VESOFv7Avypxp9zA25Vb3if2mj
f/ad9aYygi0210jbkM+5L9/cRw0uUYISf1WPBaVXgTljRTaxEdbJVAyNoIQHvt5/B95wYbAn/yq0
Bv0yt0iKr+NDDcLM1fBNuSGKj2Ebm07DkrEzaWR6XfnvFTX+kID/SgRG26s93Mf3Q8Avfef7KNXs
fQ76c6ns6ELlvkyQtoyVj+wvM2ongcRvpIx6YBIvMd5Z2vSqFBrbw1dc/WgZMKIzpdSeNRJN0sEf
5SI6SRs03uK+X6+I2ma/H1KTYpNpwPBCKmMtqQPx7MCfg8E8/bIU7ckRRKzPWkhcsElwZqDEoTEB
QBD0LcaIVqOv5zCoc2RtSszGg5ajQ+bML5wl2gxaZKjqHWIhSFOucW+8fip36XV6r635a7yn+WoW
YgCF3VIt3UIIBTOl1w0Q5psl5vrLpTpR582YtTWBDbZx8cnP3vXrzMc8Lx9oCOv4pyW18xT1AGKV
KJogQ6zfNA3nwPK+Lvk69QpU0DUAC7E3/XJ4cMrQ085Uyz7zO8GeDtcWNT1sgQNOQmaCUuwtao4V
Cg+TRIbn5izkudBimpdzTSCLeJgCGjKIPuYRIoEdx0WPbAxWGgxERYJwmWJpLHltYb4DmUkeC0gX
H7xtMZFl+dJjXl6Ya7gNeLau3jNUARkH32oHf+I2FNO0mtf576ERQYFAotxMdThp27HRDfh+GJC/
J07Mi/gQeqIPKxuHScnzr5NKPufaDFG8UnmwLE80K3XN976HKdrM55iXVVqUF6NGnmBavXcDrPtT
iO6Aipx6C7o/OBVIU/eE6DOeWpib/abU1iONbhwoZa2nZ1gQhEOU6Zw7STNeSlP7Xg/tpeySnCol
FdKSlC7ImbOpMLDWtY4Yi3BDHDfumCEkre7W95/derjIi20/j9Z46z9lozE8qRxM/jhcSlXGqxUn
tojvMKpZ0Rvukw/u4JajZwr6stNfScV2WXZtTeiLcaw+/fN+hn/X+ToRe5+/czxsHjlGmQO1xnrM
cGZlUroXX9lXz733veHMGJSFrw0RgzGQtRStqRw2HpxDKbko34ejALZnTK2X7HLtGwbN36RW6ygw
DR1k6vvJPBVGlT1ZmsH9BMf4n4daVwGsLy5IAvgaE9HpMJAw9Q6bjyLdITD+JdfBVtoQxt4qTwxP
IpfxeUi3RxzREKH77KQAnveMU8p3fSSDyiL/b/u8QLkVvP8WrLdi8DWIUfzbh8P2G5JDbIAArU3J
60xDItUG3t7Lm4EgYd1qVkZL7RR50Wy0Mv3VvzrL/SC+3/fFksWTU/ncS98DiUeAIw+2bu4X0yI0
zRiiSUzV4ezIIeHsuHLuVB8cqZhVKHfDqqZNoBQx7HQfDLMeLjPnE8sVNckq7VWz3loX4gsPgiGl
6bsC7i+JMy2UJrI+O3UddkZ4wh3SaKN7qvKzTXnm7qmcfTWRwE0lFYk12TY4PxNa6G+iyViZWVC0
jHbTuNksGS4IJ303KbKL245sJQLGpMmzEsapEirB62+rgj3K+m5o43Ex77pgsb+TM/w1ddNfx6Zc
gfWt8Rm0NdAo7/UhODWfNMC5bRTJQ6EUf04RxdnSRs2nt8/2aqffE5uarS4PBaw55DOK10kPgZEc
IC5kvoKvUOWtt3NUw92vBr12/E/s2gnty1nwHYS/VJjng/Ie86bYv/wglZR+ElKLTc1hFbRK8lLR
IcbeNVlYl7lui3hrfgQJvvgTEUUmtSFBynphF6/yUm/CH7b/WVWC89U8GZxN51p9wJ/ib0LuyJ6r
QhRavbxYC26eum0sTwWUrz7AFtJTXUtchk0TMT0GD4IzTmTL7yGnAEfaj8N1LEW8ein9JkaTm2Xi
Mw4twTcHszG1nBCxicaa3xAQLyobDfK5WS1e+iGBhM7yqwGFAzpa1EXf6204qtSerDlVtXNfdZmd
+29dRjm56NYZnXi2IkEVpr7awiRmTSQPXWcZzdpfQpaRofyiptuCD1PI8dCnn2cRuCWOte2l+9UZ
7KSqbDHpXw7YIunDtTKJGMy+e7ZZFN1gjnHyAcA6ejJV2R7dB6mknaMwJmkZCobj3XfVW8G5Qdkl
aq7bPS+Bl86pGQ25xstwazRSZZ+usYOa+LBAu1MIubq4IiWdq4BLTGEPD1jyugLXAWjRJ6XUKxPZ
yZs5iM3CLqkIG6yNlJwjBYfIVl3wh/SiXGaWLcEWA2q2WAAV5NpyG14jJjhmBaw6a8ncsHhWOnWp
hyimlcFMWoxLkPHkmAeJWACNpc5LctQ6+iHbOa3M9/bK/oUMOV4cUYua5HdsqK6KqFryXJpantnS
jywYKynRzNYmZoV/L3GHPzt0XZYKGXZPe3oxN4ANkv5bMjRLKURJlyTUQx1EJUNZahiW+D3CWp4a
tTt9LO8hGLz7KD2e/VFvyUx0YBcVMaUBGWcg5LdOMCYzzGJvBHOsCUwXLxnwgCCeWx7kAdo4nFUW
dN7cwmGTqsRPW6ZHA+7SVDdAbKRSgOZOmRDU6yyejtc5eizlpcqYCxsNK2zXXuKbionGvTw32ou3
c4WRkBvrbRXopDMAXx7/V6geSA+EFTRtrx0mwu5rXcxv5g92POUXps15WwdB8QTf6v9QB5L7lWIi
VXN+uYFR1FVABlVzq/YSgpmagmFXghHjhktM1mEsF63Rw8yY3bskJPFE83uJzut4ZjF0YLh0QkYD
k9DK1ZjSSOhKNlqE6tTQqmWxfXay+m86ObBslQ14UISCoR38ZPDSwzUW49Rj0L6FOFafnCAjKBxm
rSLybY14/f2ZxMOokptbmwC639xkZcIzo+Kf5UuqkgaBGQ5EHZcZzWGVeB/ZAkpswZN1zRART0Sv
GD4XXNaZFxywB0re6aWHH+xtVhgDY8rD9+30FrCVWZGFO8ng0LnXsv4Vk7r/irNET7prHnnTRU4z
J/ujJPgFAICtq/EyvcY9buP+5ZQGp+J+akllPFr05979GyBWco5EQOpy3TG5JzixhIm/8rShTC5I
Ie2yDfKrkQWxWk9ybxJ8wMbMID5vgEDJTi3mvibzKZsnxTpGXOIHDknGOMlpejaTunP1j+EZOomZ
DP86bAr75eY15bpr4y7AvvA+pBAJpt4g1xSCnqhQhBO5G30/abfdNBF0n1QtIPF+0HrmT1IegxHo
cT94yil97SYEQhnhjGGSoSyytc+qbTaRKkokXM5GYlrv9BPDNUt28Mj9HRjmPQrC3IYs2QcZkwQa
QWgQKj1Q0+PG3Tu+Ppc6SQoBlyGycKwyhAb1LIegkXcbvZ0lopeDGMOYVgtpIJZs82ihEAPGnz2V
6YCFxb9UurFmXWD9mxGXkQh5aExQNUgzxToNvf7JrFvQtxnZLW7egKwn+hxoBmJpMgGCCv5yZvnG
gapIAbCKAVjys/c2JRnSYdHL9aZ72x/BlFVu1LGC+WtSvUQOG4ogkTkGEp+MXor/7Cqogfj17SxI
2C5mUvGCzUwLbbaE+Uzbxu5tHwUqIuTJFo7mvkkM7Z5FcG1eIM6twcq4bG93pyJzrq4myP/4XFQk
Flrr+NszRPIsSjfRNXAKbFzsO1Q+13zwEc7clAyTSPgD9ZQV4bB0WYD1mBFWHevKGCwuiZ9LIGoS
NFR5cvjxfCO5GQdBBgWEtHoClExYWAHzHpgFG6kEWfIpYiTH+eQbQxe+K9CGsXHFbqKY5l7Mh1iL
2F5NxdLkkezLlNVGwg0cvKNiv5SLqRullYfKQxnUqor07/c85hZFKNisykoRLtCTSGi6weUj4ToQ
x+3ew6g1STfvBIApHET1mT1FnWDg/KW0PhI0zyiZSy847aod8SdMM5mxudmDwFfjxzs46ozTG5yt
AbOujmRFW1PaZ/w7LWQczWq60eOUsLfbFuYo0wr1wOIWvhItxboMZpVOMbYy3OqK+dwF4OLfuKSV
HKtHpoiXHdhXq/LnkJgXcIAA9uo6qclTRy296WHPHsRg/EHsVsLhuMoD71VkhnrTJ+6/gGkkTNP8
abZ1vLrd8n6Nkwhf6ooYrdbHP6hgXN35uBVFYAEPMjXwG9DCJx252AyER4Myaj/+1h2johRGIJ4f
VVSXCN7OUaxhly4xmJU/fYijSWfcwY/RJw6afSwVUwiSPFr+VUKvj4uJW4iMXlfHb9/eqQ80LLQB
K86ZoWOJEHIsIxLOZdgJm+OmoxfwON7sw45OoXn2jSMy3Wr3NeXS7XA+yCyXtbjtoDC2vAwnAu9+
lA9+TVxa/PJnuiF/4nk2IJevD8soNnt30R7iwk+HN6IpIvMQ+172QOvpoOJkYEzdXBukzVBc56VS
YdB8jJ8hky+UYA+i35YVBRZGboYMbYubd5WiqGN3f4ppwy8WpXOjj6dhORf9NBY/RkvtvX8950Ci
8laH9vXadzKIWJ1FvXP9gExMlb8+CjdncudUjcc7tIy12pDPAGVLLY0503pkxBiK6eEL8xqFDcxL
VkQL5txJpHUl+SsXYisQOdMDiNsB7jQBAQ0mWyhdEB9wqWlqgGEm74JPxVrgur7/Bx8QBHhQa88R
EQ5Oh30xB7McfWmXC+zTZuaPID/6x9wsnZ3OrRDJQ7hYNmCBYMzPrxE00eZvisJi9gXfpIRTC/vt
We4Vh813PPPixu6FFujAO1yTRGsJDZA7d7gmMUo/0OGnVQX8fOxqSKdx55LLgc3ublH7bhGFLVp2
2lTdkvnL2mvjqdDBiAlesoJW1Dy48j7jf6uJ8XOlfIL3UQ7b5dJFfbEmfoYI0NY51kGQGaY55o/S
nwR+mZe38CCpGPUhLcZho9V7Bqj+CcygoQmqAUjkTgmaPP/u4fLyDgWXcN5N0yZ2sxDSXSniAeX3
jYEqaf64KxeQsqsh7zYxy054yc5Yjj4aKvKjrfsaDS9OOp7HpeltzehDrRYeKMynxLvXThlS7MXj
rNonM6O5qZrkkA7NE00QxkYSg2qt/zVv8t7jcevzqgsLeuu2dyixxC9FJXbUS+z9uGM+XJuidbGV
CwcNZuC9AsfQZ1ow5ZeB4ZZANZk2njN//xzlnDVqhvFABAxqOC6n+ZUsbaVHe+K2k+OKM0oJYttj
M5RH05dysFIVkPVIq5PUtDiFrsrMeTBVXE+J31ES+kZBrqQohaGN6I03XZg/XwupDRrvN7LTYIuO
FQ7VodGemVebc/XycDTA8IBXXiUgmlXy9aPqKD9k8aMmrOnqgdu+f0eINCYGjuvNAFHpufHK0LJB
FH/6rLGDGN59XbWeskXuJW8hCkH/mnpMAdloLIc2XDZ+xhuA6iWInc02eh5DwM2s1c7PBfPaxiIP
r9uyskPq3YocpHz+jGSpKP4Ow1Wf2iewurVQs8NHhbBMAmunLny7MhdwGls6IWqEZK66gq/bZM+d
fYZmevxBsIOn0u2rnmKO5AlxKLIubcVW1BlV8yIAueDerWOdZ1WPmVBevUN+0GjS0BCn46ScJdAJ
B2WPglfCF0DMoYZVgfduqQPPOA0LdomhclxGOBWC/7u+GIodSNhy/wc9+poAOiLWRBzdjb0hpayl
XAAgRmnfRxeMKA7WsS+AJhJvpmAG3JO4Y32c5qjaMDLO2GNAjFBUmBLcAlA+LbZF6FzD/QkI1AVa
rjjxYiM8vqOVLZ6sQYPXaqjXKBtrNAYyRfmM3SrOGpFllx07pRhDrIz/xOOzRGRCAkphA5+ZPAx2
AWJED+FXfTExtZUA5Xev0050fDD1IMcr+3AD4JXJi46imC/JDUTtMeuERilH9WSSrfsCQkJ+wByy
oOVRaSXnpc0spoNFuyVhDBQEddGKyD3BKUQjCkvQxgFlNW2SCCkzTr1zhemVqKEBsqiEpKSVNAwh
AN7/zhun3HoAzdjLvZ7ajncoyv/JDrI1VMKBVgtFUFuvKg4Ds/ReQMERDqi2mJpxj6tAr73JIFjl
7PejDli/4Tm0bJQyjBkCkXJLaYfecrjxNXQ2jeduAZ2kTiRnb5WPScx0gBNzMnJh0YXyCZb7MLBF
xc7xeB+x+biHHcBx1Dw9ObCPc8GJVM310Om2zbd9xS2UP8cmxkc2QmZrWDpPQNkIb0IXZyS7oYuz
D/ANZLSfZnr278SBhguvLQyKYXadVttAKmy4Oll7uqorRCIMOv27UNl7hsp9ZYi8Hs7TZvf0jrnp
+FJjJuXDjK4jqWRd5xviVz7yoTwThohAzrIuNuHb9ro2igR85s7JqMfsZrg4BeI9DFyZHSqqRcXy
cw+iVdIm343guqzL9N+G6eeKQm2a+jh/aIRWeH6OwxRWj16bOT4JezzZxFcO/+eTundURO1oCclj
GZpNc80csEikigKAo46BRW0dw4kbYPpipUInt2JdA00Bdi/6fFMJtWICXTGolN+SMyT+nxW7Dnfu
RP/Qrof/u0R8hxk80jYBZgEyiU9rQw3448dRyK2FjFgDA+HtuUTfYccDtUD0/OLZ2pSj+2MgIyIX
OIy0YaQB0QyoB+wsV0I/rn9kmxEYhCpJdviLH9I56vUlIf7+4x3eOIMXSf7VMD8dHbZjLrt4miwu
d4bBqX0A9b6sC8puF7bdD/KpAZAGsVIfpGvYJjVrvMWAUugxKSVMXpbVKPv0nseUZpo58FJ0y50V
yTYrQeLpOZuA79oGJ+2WZtK2E/KkSgGsMAeBB0SajCQjtieyW3JIY2k2o9Y7pTfnlo2f6xoQ+BdV
Tc6O9jdwTtave4KCZ0fvYmaMGeKGzj4N59qFXU8GFP+svObmA80+Jn65IMC6kPjt9hApm3LCoPpD
ot1iBQnrzixkNEMBFuyOM81As08MqAbPo+Ha1ClfWgkCJSJ3PIlXZIiUICb/T8sHXyORO6B/iflB
MF8DtJOOXZ8NJuG57h1MzDL817nTCu/mCpcLEhwkcC7Q71paQFtFAdsv/pnqDTDHpPIROCCDYIlr
n9WvoNidVFyuvJ30nHB17FiKFENcNiS2f8nBb3m7jFxssYZIWpq9+gSRCwWJk8ApgWLSVHOrT0GU
Qr4d1ZIeH1PERXr4s2s55eGLBCwyCgjh8hRUzue+XClMiUJAFqez5Skr41k/+bWOTGD2468r9X3I
v/q8BFWkpp6KHrivk45k1TvU/x5VABF/kKdGDCPfvdmtjxcbUfFjcLXhIRntGBOq+zo5ejjFpkKa
7PBfm1fT0hzXx/Mdz0hUiMs2QTE6U+U2zdWqFuZ33+qXesgaw1ndpFLTNDyRjVLDwVMEJD94Q2AW
WzIV6XCPhSXFw0/orHglqVMJuGjheVMWN3TJzUDF7HFgyrmWWlqvGS8X62RYWX5kiWFm0v+SjS3T
LGuO7PPDNtBn5tnYNImRgZPgBIDeX92gRYmK7U0ozyD7SPnPkHO//UjlFi+CwcbkeqUkO4bIKHou
NTOdXZeaWg2QzBgxFwAVndHsn3VRFl7NclYSmwFbZhyd/9W99f2pu2i9GuDkqhCzOLAxydYSpfi1
vhei/Lx31BtP7LKMKPHTnM9i0apvUeZ1UmszKWg7xZttolsFRlWaLsS5LKCm3SHkH7/xhUWwJYKf
YQJcVJL9c6VyOrs9B9dGGZONJzOOurxDqcdknUoL95GV/yLfyx8GSAEjZSA5BY7pZIjMF7LrcTyR
kNEvpLm3jdBVgikgcTvuzgw9u1fLt5WRUZRs3nlJzWDvT+7nQbh5BSHRUh4px/c8QMzF6vXBJJ7a
jH85c+gHxrtwBtywl87/mRX6+dCMYU4kkTWwwbn/J/EDIwExcM6UitRk0ch2290mf4wFAyLr+FeF
RU6wrYTRbnlvQtDcKJsPv5RmOdijAMzglfmqA683UGPqgeIwgEHvjJV2pQmXmimswkVX3ag7lGji
V3Ch7gACydwRnET+VkKZSPf7XrVUvD/5CR3fj3VB5uLyfp1hRUOlnC+B4Ip2dJelq1JNcSu1ipG0
XmpDV6rrHmH5/1X/8W3aKbTkOukqipAnJRntJsn24vV6O26y3lFuCMnB7BGbG86sUIgoBjkYw2cL
bOQavepha0d2oWjN4DIlOhyp2lA8HC7fRWfwZkZFpxdhVFatJwGz1ilB+XFWKHo+NuUpNeZx0D6D
X3rQj9m/dRXoVC7mm/YGayCp7z7KLhQl3K+TzvruMlwu02gT5glW+MOWt3BXWM0EW5QyaFdKoyZK
RkqqJCPVC9draoL+5oWid7z+jjJC3xeN/I9qrFAXj8FhwajJo/uwhBXLbbQvC8eFUSqXCOS9LF8v
B3EeExF8GEGt2wUwmtiDf28ycuyJYgv/JflIv4hec+zwHrINh6tmV4OONQzNgBOLcjc1fEb22X8o
G7zOwkUZsZ4f9wppBTxmCpocP3QIQ14f53lb/REsfrgd/hLirZC5XADYLTyn30SMEbwoE3w2dfIy
7Ew3TcwA4eC9vouQvkR9lrBXv4M4fWSaQ9y2LYH4kZpKPUbj6GNjFeterZirnajEf/Iq4uurSscC
2RLLEm87k5Rqgw2BPMR2YSMAISJSNbVD+j4isUCUrgcLRyPm2h3KY60Q9eEmdAYfQdol5xO9O3dY
zm5lrN3tk/J2jnkDXY21O/NPWdvATMsyqZx+kD0c8akGSHT8ZOFmpNZXonztXv25wa671KS98dSK
2qOinBd/qCKPwWDpdcUYeYG3uamxvGD/t3hzPXfW+RNX3mRqoJzpBjvQ5od7O4HQJ8TyF3NW6PP3
MhoDJ1i/c1N5YDEf1Hz1YsvJ8MvR+iN1gMRBaVxnCGOAZuvXWFuLEh9kl95DQu3V7evyJH/xMsY7
dEckTYbnd9m5YeCNlzmoZYKZQqMvTcW+2zpeeSNvqe/3N4YYhcTe2m7JE5J6w7Mk1rDfwvDCHfjf
r/2L1GUFERlk0Xhn5RBOUh3khgLfjdf7/ViHP8Grld9BTPYtG36976vJEHNORtDtG8CrK24kCgeM
L4Iam4IDTUPFwraU9MsQGaPHYNRuyj/f+2tBblS6kOe77l5BzpxomTziXttMgH8kKCPiQs/IfkSN
abDIuvx9CbeIMiFDYQIOR9bF+NeE6rNjxX2F/eAvyevDgWShmDZZhRCnabUBsvrpCGJJLxnShatD
sgReededmdigrrrkKBbx+H2PQQzGBf9ptT292qWNi0YZcub9kIhbaD91Sjzxe14Kk5eiya/06blJ
1tC/nY020i2Fj1vaGUdnlyS+QI4agFuMPsWpkifJ9NvF1u7qPHYeR1bn1sMz4IUgkrJUd50j3P8o
fxfY/F+fl2hfdmkoVZlQ+dmwOQp5GobnD5DqIPc5q66Hdpk8Te6/UCFyW+CVroAQoj5WC1LjftAT
1ytvsVFFjun+K1US7/7ZCeh0H6jKKLMAwZBRmt5JgcMX05ilAsB95fIIPzRYevKS5mvLZ1Q/Rr+q
gtvS1Wcp1VtKmnj7Q3pdYlVoz2lrWcFX/JpnovKXCqhClqklTWe3j+Tt3yLxPZq7NTRHa3yjwhWI
B+DB3j4IZIZOAlAeD+L9af2aYTJ5QcAAyDYUfvcn/RKBeMBCr5HEtNmIRIK/XLUZDRio8Dd+IBDX
n4fxpoYB2Z+f8QPf0CSH7hbxIBvXAixk9JwhEh1zRWeDPRolgQdht+ur8ARp5dGiodg3Pfn678DA
GYgptMBgfD5OKnm0d+XeffPNBBvbkr2eotAPWmEpJ386vuxV0u9lX4FlNzFYmR5I8PfM3REGrXQC
ASERMmdKNZJ9C1/Kghc0r4KUxcrVUQdsTk+ZNs8vytXWaZCE8juwi9Kt0PX1qaSR06HEZrpsWYyF
YP74GXIpoBrhpecD7x8BDskxDaQ83zkwhVgy0mt0UTX1G2dip1B8JWOjunstbPXGaI6xPe/vgLqq
z4hcRvKMVYNOVkNVP4FWH5qwI8TC7e83bqcnPfvGfGl843LwU4OZRHgwWffzagJFnu9ANalOKWoN
acbfaSYdutPrYF4giAoI3X4Lwt/tvmxSzlJDXIyNf3oActv/BTHQ1Hg3LB+wxItAnmjUyYL/9xk+
JNpHcwNctd1jcpBWwvcacSSlJZsFT7W7K0No1rN7CpTdyjKj3+Odwr918o5ZvjB+lbQPaZmejYoo
Ba+mxxEu1+TqFtUOh1ddigTb6uhFe+OKxy8/36yfeQg7kgIqz+iXVSxkqfDsk3NY7Z0DWUnM9qwE
gvlYioE06QDyapBycnWX1JbaJJwCPfOHDWiw7J9eRsE5ze052b4SktWQjAqyqUGRKJI/Dp617KAD
WpsKT6U6AdWX6YodmkqbhehP7qTQ+ckhVwZh2j4CK+WDVlBcvyN4Hpm0DVYWDSFDA1ChrjfJgYng
UR//QmT4mKWFu7r98woFW/ZnCMrrjquBxMqUdmH6CZJbsOL5roTe+oriBc3ipd2KRBQQ6WDi5Xho
UMekhy5e2aZiWrgWLLqswJ8p3z40+UGMsOldSk/j+lKdVqDfFBRpKIxsnadRUK5Vvgpayn03QVO+
LqriVcdLnvPGRJHcSNzDFW5J0iqUhwVqWaor8fa+uRSZFYp6OAQlQnmn93waoXz2CBHp2pXDwv4K
yRzjDPuvGBWBl5zISseHjkjbnNw0abwwsjxHCWBhEXZ4uyY3a4KEolwfiage6ETBuPr7miFFp+tg
G+R2IPOaaMOH/UD3U4G0zEJpxWP2Tbzcbw6CxI/WICMr8xA2pDxiNKZ8ib68eosTj3qhldE+WOyt
RO9fVEWoym7+VqJO72PbEDOsfc9Y+130d/5BWO31XwKTOTCVQHXcIFswodbMN3vplbm6Lzlj7W6P
eQ1WqL16ZcFmV5qwdHtVkm0s9vwNkMbbif0DFu/GoArCCXOuqpborpCFUIxObFthscO1MgUP8nOy
2tTKBhR6F+ThmofxKuTF95H3DdbQUtlMIGfJ48IAL7D9HqzA/UWPaVXvu2tE3uIW8rrERWh2rDoa
lcXnEicj0myv4qoisqBeFleThUfUic7KsilFeNgfMiPC48U+abTLO/k7pVziMpy1VAm153p4iu0Z
sClrWh+Arp+uGQURAXCq920DEUQ2g+eEABEhIbZ1BRWbVC8gDorohaPfQsKVNNQMZgqqBIx/Ez59
l/Z43/8h8GbgSPloOhyrkdMnw/qpfdC0QbOjiyzhrvGd5uXZt5S8sZz0FvbSPk+VpazbRdwiA4oS
iMzh481s2kAy/2A0r1CygsFKMpQ9CJlZl6r07snw9+5s3k5P0qC5uq/R9OEZHrZGKtxd8IJ4X6sP
yXgFd+Mnl7Xc7zjwXrxWjKweCMShPGqHEXNflpYqLOhlPYNEOD97/wKypMMRDt75n7xsE61yTtV4
zwY+/Rc6TpTvHrtuonR6PYLcFPRr1fyKYdyD/RMECt9PJoaCsTsryAAM1U0ZH9vlimrdw/j1xDGA
dTLRCyM2Sg2ijsPvEm7mWbqtHJumA6Uw3mxMmq9B6VRB2nIYRc7U7vj5vTZtiP2qPDRDZ6sHxrkO
9m8l/kcU7uE7gSyeuS2gz3JAbLlHjpxR/mKMsDUsTa1DQXbxIaNESVoCF9U8AWzmaX1NW6fpGgJH
jQK7gr+uFSFthOzNKeVtR7rKemZ4+ltbkd+lI99KWIimx4ztQqalC4KsEKfDEqGGRHV5ALmxzlR7
tOpRrBM5ZFQQkICPxsbyAdbSyB3XOUetkz46Zu4O3Lg3z8pRGy28RuxK8mS6EIv8/+pSmvZMjgEf
I+fLSc3kIFCqll/g3AF1oE7L6gWWD7ZUUCEMa7l3KumNSEf5VjsXR5A2uYnjcyYuVKWbqatDWoft
Mea9wVaKKOVHzTGa6WZVNhPp/cwYh3m0J1BMe9TSFup6la4o2AlSyx/dkQtFXnsmVNycH91NFYHe
WyWqPlIZrMZm7/JS+WfXSZe8+ph72iB+3q/MJMBij8ZL2Ifg3POQL9Vy6YPkNxHWyR/TUNb4xM0W
VOy3GO6bossuAo244R5D/0htNSCEpNd/vIJZ7ciEqbZiXVbP9RSfCAKtmvcRjKZHCGTvD+DwLoJV
D6DLODagXNeF2e22lnU1q8DXTwBPQRh+43ViLJJTQ/3gutjj1thyTEke+618hglKSIsflnacT0us
hVIlz74ncRNDlddt8ynSXWiAaNx4VHfVdesevxIbhIb8yGLBZ1aKCge71aThdcSsdqJ5LS6q5r7n
jsP5C9KWDQmiAB3gzrcCL5WMh9sMbhyxNTpHwsqx8/GFd/AQHBsI5HatQv6Ig/fiWWpBNoM4Ntq8
5AvRduWPCK8LMnFVUecbAg/Jwvu9jaXq+IJQjLNtCT1ZF+KqKJXc6afV6vxuTMybrFAPWR9ueGB9
Dm6HVD6bWGN80U5et+rU9vJwc+Vnur2zKA/UtK60gj27oQg0U9ji0+rt+gv09IwGdFLoPaQBtrhN
ndPLCGV5VJCB1+ECWxYXDmgReAmrZBdNSSeIsmQ2hnBczd5vY37LCj0Z0ptncPIPmxkUHIZf2OhG
xbeP4b4XdRM+67VDJrWEGy0MMzLQteHBf5MQ7CKu6LQFvwyY4xu5H8hRPDoKvXGUeb3jvxOUZfWr
Iy38hdJ/P3ns2oPiXt3IIr86XaECzm+LID8o+RpwzH5fKTQV52/jNrp7/KTbh5my/FE7ea3YlIpS
0nzLepEYXbCuelZlbEYnEJiEuSPYYP+QEPwSJCirwI9oeIt2NozV2+Vhnky3jw/mJFS3jWlwFy9b
06ijJDanPDWcnfPAbmUH9YexMFgjUaJUvEdECPEoWFZMp27HpUS5XDmmriPWhuPnXFDmBfZz6xnz
lPyuPPf+3V5NSkHtlhcRmcTX+lh1cSj2IDOGsG33S7faC2UeKmwiyGNJyi+GcoAPoOvA8OSfomVf
RH6N557+7jzlZf+mKiNJyfARAXO1ExMPjb74oNAMI6tvkq1cBJffwVvDsqJwGzarRhZs+9m1VZLl
bmdwD2MiUAzKG9lDKjOZ4JUl0wvxeACwP/z3bG3c6Z7KXTyP/7XLXtPcO3W05qKEXGm2f/8PlD02
sNpffxvDDVH9NajxQ116CS2tfm0EhginYkbj8rSQdNycG3MpuYIWp5GOPlqbeDgC9uV7x+iOG6Eb
bz+ZZjQ9ffSAJAZ/BNjwcO5rUG1mtyeUmx8IMebEUTXzdCFbtuZl7BINAp54E1ut6ekendvTVEYb
gnMt9iGXUJTaZFnmF4IVWE0Bxs9QnfCvOPXFrq/1TCSIhSpv83lSBidLynGwLsoiU5uOOev/lIhT
lDGph1PUjZOpsMOnTd+jcT1A0dP3pZyYViTv7DWusI6CvtOcU9akqCawgixkfW1JL/xROuN4ZXT4
Uy3/G2AU1ScthZ3tHhOtcKLuRX4EWyeP88GzHQzAq9QCtqRb0k1JR2NMO8ZVzAocBqyqXaORivqA
yenwdmxwl3744gbM2K0xbsa3bqnTXqe85tcKcRSwsIISLKSqrx5RIENMdonyybXlxnfE0sfvIoAL
K6IkqJwHnxOtH5L00GgL1gPL0YsjCrhnDxrN1SOHNwyMU/CNXzfPqziaSbRwrDrQOqOxYqtXsIl+
ElKdGC4mDRYZTWGHlIeQqfgebF5hJYe4decz/eHfJN1Q1klPhqGTks835zNG71wrOXitKVcZTFVu
bnK/4SUlDSo9LncCE0O3aOH/atMQ4pLkrA7yCCRmO87YGX+2w7O7T3JLH7mPL7+SoZZUDK0KILn4
Dxg+VWI9K/VYbZ3AGPe2uLJmxCQxJMnTcUTQ/A8ZPUPHKfTi5dcPQFd/wHumNW38/ryUmhhK9iyZ
wirK5TpqpXDu1UW7EHQp8aAYJmhHe88t2hoIe3cWiMNfdVfLEheS/EQJ4MBoVT6zNmU5Ojx93/vl
7aIXl0KDDKhoBN7Tk6we7lkSGzd9iSNBmVzd0POUtiQqMMgMjF6Pc3vVp/t1cE6CsKdsoZ/MrSiX
lYp8CakZMzvCZkHnMFRvp39e0K/kRtXjbxYIoS22HOVK5ycwtyF7ahrgYC9ivXq8hb+VcYLItxgi
W6Y6KzeKxQQ8QlhfF/Q7iczzX3yVEYhP8kv9kH+sgza0l9mu8g+w1l7a3Lpm8fdLug+WGgLcj0Vd
vWmzznDA9/pcKH05UAPnVA9INuLrDJ62BXla68l4+t414ByY8430T0bsyueqznk0Yv1F30SkVpOD
pRVLf7t8HobtB+uRk5Mv4qKMOkfISOrKXd8QVN78VlHQgU8eGZ2FOCDV7F2gAMSyaK5hiLgtK4cW
kCx0FsYoucPKUIK/FBi+10PZA6AA9s68XFw3hvLh6Wc48HhsGSK5M4d0bprNM4ARrsym8XQone9I
SVYcDDk11gdHRKPvnUFwQ8WpZGihM8aNWhJqhLwE3QKin5HlP6oCHvlGK41wjhL6ft7qsOJ1tiZF
NLIuhuhD0tTw7DTxnH/fRjpNEMKFg+JQbiPEbPZv4ZxaOP8NB97AP/yZZm3HKPYFEYN5fRY5DZx8
e/crzdNYQIJOnedI6/KJDwSA+Zh1iZDeJ4eob7YDpr2s44jOnvr5Mv4iJsmalG4AIPLBAcprtg/8
Pq73b81fHfHG6vJbWPyYtRCp0ZqUnBG5VShcXk29g1cWT4u8pYrB0lNyAGEjVWFRwuR4N0Q6kVMB
evZ4BE/Hf2sjCG+Lj4ybe7tHsuElGeqCeOYX2eThmeBTz2POa7clY+kN8SXQWqYDBnAUle+T42Bd
X+Wf/DBR7Dzsf/srdpcGRPpoa3REefKGBR8r1Em1SSQHXrfj9R4FcAc1H5l5ak4dxQeHsN3audxB
E+cFi1rZnhpWfna5dHhY7z/195Cn/uyZl17VN7f6LCGyPA04M7IsLWifR7BEa4n6VStB0Uq3JtaW
Xlwba807MqPtyLUrxYErscURfwjx2sBUKDyiyN3715VuwH1C+F/ALAaqMtkPqo/pZOPSoZP51/xv
Vlsj3f5teqbuWufFLLGD24VGR+p+Kr8sN2apVYk1mfaEWUZkqbBeEAM+uMuQ/RrwBAQ+SH11LMVb
4HTs/Bg/HVXwpu1esru8Ytv/cXKaIFXp+lRgvCJ0QwoP1OSMGT5IolgCHtLgE8dZ++5gD8B2eUbQ
HtIoC2hJXH83ZiT54CXof19KJPbzBMAYa9rwCnNxM7ccgk2A/d6MvDe82CX8fitCh3o2+J+bGmcD
KKm7vJ84faF/yT6AHSGKEyvBDMSH/t/VaWGfu+xJ9uTvgtExD5oJA6QG6bpywuCyiT1+S6l8EjJN
SeXgLVx9OxIwWv5pO1VS+HEr+UCuaEm1EfaCCjO3qNjlqtDzJcxQGhFhQCYkji7IVpU7Q6xSyBZx
srLf/o9fUM+y5TbDQChrbMP+4EAkUo0K/C0XhHRes/1TZc/r5pjGyYCLGXocZt0GLCJL9nu73w5r
i8uNZnJi3nGEiDwBzIegN8oM3f8oCYaqSvEMcb+0rFObQYb4hlYByZWYpYBUN6+oDP84oB8Lo6PY
HUdYu3gczNYu7kscS1ALoOKMyXdyR1fiMlXPltBcChpftIQ8eMHBQddFGa1XSXM+qQiSjLw7eVG8
S8jCjmJO03DrdG1Z3SHHUmzPbwBaCobkG6KeR6N8bOQ5mpuQM6LLXb48Vgrcw/7cuxdmnxwqtluH
SOr7GhzeRvNUJY8TwBkGzEfo82nelbr2JE+OuvV722IgAkF65NYnRsG5bUDAkcoy8B6dy8qcDs0Q
zdFXPor3i65U5oAYUnPYj+21YyV0YzLbnIYIg91TdAS5Sdwtrcw+ivFdqQX+LZx4GE+efcvP0lMI
erccJsAzPkMTpLzoFu2KjntBneQ9LhZEvTRPiVK/yag+xTtZlZHjldn/cSQjgFVue4DNN+wS0WuM
ix9wdqEiAmZrniURnHZPPjHioLcUS7nb6VQtGm4efFRO8pi6TSTq7xIvt20RbQotStsNruytnswm
eW9B1anZQWJj4c8Osio+BYnDPd4jxshBFJ6omxu3rf+jErKoibp57+KeeCuDEvMRlNimabrdUvnR
J0vJJqVx1rv2IOZ4vdIzEay3W4nGHJyVJEF52cyIeHhg2QXNxBxZeGZdsoui3FjUtTyBjxPGZ0Qm
0WSG/qpa3W51997eIMSdhJ42Jq3LfUbucjCqQ8S/xYfMfTp6niMEvlRKQx4mSQSCn2LbYjfCU88o
t+qv/bwMPkxjneK0QhMYAVv57NrqRMrLF10KL0e/HS0jFYhfBMv6Z5zhnFkzreXYIq+0vyKxs/TN
Tvc1uUNk2hO5mTKhzC18l4K36jkLq579Pto59sHxxCceE4mftSXqYdFUIPc6yCxyqG2aDPTMet6/
uV9rZPn2wW9cHCuLoyXrJJ5pZJczbI265qibRR2qtEr5VpapLTyWEyKe0wkY3jyEk3w/jiV9Z4Bl
Y09dkIAnA1q6IfxlUcfqmRB8d5vls4CfTWYJtKNY6FCuU3/d5iJpseguLFVWFYs/dtj9EfPmPDq5
eXctCpa+mBNmtwwtlredBUZ2zSYQlDdmosN52NDPLAtiSGkDoDivPO+kDK4Y+G003yInWkV0shlT
RjNmB383XnObv5fneD7dgMx0IourtHsVTf0PxEda1k1mBVMTSukRW9VJI17+FLVER+nHW6ZmKFiR
dpvFlJjoqBS548ZvkTEmM/GI/N0DzsXWpUvQ5jCej897rLLubL1F7QpcpjwBAMX2L9Qi2AkTV0Et
l/SE0ci6Tj0gtPdo9vUDSX3zjj0Ie0BdehVWXI3Xt7lxGNA0UPA9r8uQjjzRYvQyJAjuSpUR477S
ta9hbZBDOU7rDwmz0deTKPuxElJzAYvF0VshTUapmMXbYUepitZXpVXTpXMn0KNnV28S7G0JSQZq
LMD8QXuh1kWfgkkY2f7DVmuYOWLlmA0DFP76dMi9651OEBmmFqw5Hy0P8T1fWyApYha8Y8qUDv0p
KwyT0iDbfa503eAYBI5CO6YviVdBtwJrHH9X+eCsyMZ4jTvWxVyUQ95gkF16tMd3vrlzVfDoEUYc
E3W/K/4oACOXPOpU2ERTFZIfQwVbJ4Kp5IywYkYlK4jxpujSyX97QbCCgdQZwkXhWNAlNLFoETQ2
TFx0FVlEp7+RX5S2ixN3z9KwTM3YZAtCAvOjNBh0qFfFFhkmWpMMK0fYVF6R283iG1O8bUwGP1un
q/mKTopFy2bXWuHaemwUMPbwO3vYNN+gfqdw9RqE0ZNd+SjeNlbf/R6aRVOApoHyoFropteGRFQX
Vlu7kIFB0FfpNvLxFszJzhza0DNFmAVO9GfZbKsZTgcqVBCkGJIdHtLPcIWBCp9l+s13PhFN+/Rl
WhwCjfgHT7suBV3/BSBLzKTPKW3FVZAEalcIqcmut92UyiLEhgk8IniwZdXbXa7i+RCbdaZ6Aa1X
/LQvW619l5B6wlggd8HRMweXHvgnmS21HZQsaSv+gOC9OPgMkDAUVmQiPSPKGpTfJyr/7Ix642XH
Fr/TNM+7cojg+rS/MMVUsQ8CovwAa7FGjjVS58V73N+3WcCCm+Vx6TKKCG51APMIRewxNnyVPvPt
vmyTKoxbtHw+kNf1EBfNrigQCfbesThzGhs2EN9tH/G77XpN0YLoRZbU4g2df359ffmtjgGPd8wi
Con69OmLpifn/KdSqnUIFjFyH9Jm8OOjnorh4yhFWPWnCyjd1Fh/Q8c6qQz0wAb6rmBxq9oRIqUX
4RYb1M8lNoGFP88WftB+DW6YGPMgS1fxi2zuFP/I8fG4okLzZJX2QzwvJik8Kuii0Iwi8v+fjFHh
jLYmW7f0v/y/IhPnZ7Wh0uZyDAlyWuFfSEgv5T1ewLxAVYD/9jxTrpPaoCgOwgDuaHvlcQ0OGD8+
7ADgdVPTtcPg2YGHsWy9Mv+3cT/yTRZVWSCCLUV8MaAAth5i/rkOLMjw7qFl01qJKOKbKiLhSPZ/
omf0UKjskZcOZr+VKROKKRN+PXiWIOHsCQE2WVHW2EIGE1+in79/bLYfwHBbf2tBLGT6IWB4EeNb
AslVHvdI5U/M95PLoGEXFaZoecjYq8Yy/5qfRccSVmOBMdhGnar/MqeR5j8lfH1pAmlKA1jocTD5
rcNX/Wer7rhcY717Ep438RKU5nZdvJjskG9lCc9j6ubKSfAWY93lXfZaI1GDEK9dR0ZZRU588Kgx
cdH2tINfMBstln/pGmDBh3iAvbnZtTAlZO5zNkzZceQjUjrC7WgIEmMuUM5J/K0aX5Ygqs8Pzgqo
mxwPxl+X3tHUekyV2nuvD+Hgm68Jcz+4sJtOLhYvJVuAe83tS6/e2hcfy1MggRYj+/KUa7WsD9Js
g43MjbOTjYmXsbz4igJDIvoBTw8B0LII77MrruhFk97YXPJz0681TiOqYHnF9DVYoNg65RoJ9jJ9
DsK9GPF0dUnmvWRMj5MaSFGA4o1jIyIfKGP/MElbMRoFa4NAnHyse5hB2qDytzoitTnNHOEzmZMe
VGDMY3ng+zEtldsYVgoWcJb/u3jf/lpylt40x0pZZyG2VznxLOwJtFsK1jByWlc5X/pPUKCJgOZj
NIiwQDcBDFZwAH0WbV3bAmqlnG2TPMe2LfIQwsw1RdYLa8v8EdG4zKjrb+DIVD3nWyV6s4v+w8gE
IuAs+iC0mhV0gEBirKqnHqXtIfqmSWWADjcxejOXM7/l8GJ5ZL/ECY9zVvwmh4yjz/02YvOktzAL
DE6DnagEisUdFEvacJx/Akl00iKGqap9FF8FcSp81qwmjUy90lHM5yvcK/SmrO8h4olxCCJuHc4/
4fKv/Ik973XJKfeQcfyRmwu+iKdZKbZcjHYE1QhB6/aZdMUGco8rEtmA6dU6sE17SxHHiAl6uNol
qQfAjrjoR8sLiJ/H2q5OKtva300J5lSCO8BJ9ihqHUqnlKNuBjzlU8+2xoBeF/8eGj/qYnY/Kpeo
sVpKVQKS9mZQwDmkqaMos3VV4qdmx3C/9zXz/HoJlrEsSD5VvzlIGaCvRU9cTp2CiSIpGOyR/h0/
CEa4LQhnBifBk4Vpp6xuRHKJPKFntAempJCQQ/bG7s04C3XcmvRKmYAU2Th3DMgvJeTisMxIQOfa
+b8EDeaTxmDHGLlqqYiomcLTkLjkVcDaeK37OafyAi897OVnlxbDFJfXG3qaR2Y7iljj4R8pOE3g
/yN01zdvqXRslhu42sdKN5Ge5leqf+c+Tt7UY4Z+jerDQh12hYkBu3vfe9R6zSWSsS+6KRkYOMnK
Pfb43yMLtuL5nWollZiw7XafVqOEWAGOKx1t2UkGP685jhCyqOykfs4VP6ua38EtjqdYdoNKyMoO
vY7vXeGFZR3aiZloUowmiIaZg9rlonCVG5sOXhcQvjo6rB7lDvj9Krc9xBOZ/cCwIrMRur3aRJr9
FsOSuGMuohvZ8+HLcTuenjVWRuG/ZdcidgX0echrnuFfuDk/svMonVH5AHLETctExFtj6lHsuAsU
hGTAJYSZYfPfD60VC55c9OGtiV/zZN7j0AAksq/wwEWTffr+3+uiS3tqsBPvwIxTLVJeVusjHDQ8
3PBoAkO/kiNO9Souvps0VP2uiAqNZI3RCJmDxPuHimZcqj4UvQCEt8efycHjdz9C1PsNh3pO6Gzx
BMfaHVrojubTVtTYI3YE2i7AZts6ObtElzs4ZMQAdlbIFQHW3gOlwQB1ciHrxQJYs6/u2wLz1XQY
oX/M4B+HFX7T2ChpdRAw/24WU/lIZ1rx+KtcL70YM4LQDoJspIbBLiNX5dpNLsh7J0YgZ/MWb7eg
TtWoDhGUws/nQ+vJe7h46P3bxIBiWx9S7d1oz+qeWl+GaLcMWIukV6BUPXKWR0slVZjW8p+sPUL2
aNRktZstmW/Ypo03RwLTLvgMUTmvrO+x/YF60803kj46aaTIdfjvkzqFAi8Cc4fVVvDlv3p5v4TO
7gxgg+QfcOjJRsLENQ8yhLHvY6dt+Rq4n8JlExb6rN0wvK0QRjoa0ecGE/nxHe+dXCfSW+7nY1MN
XMFkuuEbgTYt7QuXuvIkOIysKzsdQpbfRloTLJFY6KaT3MGS2jdZgX678NtRHN0B/Ai8w3ruxcWL
hLimV07S89w9Widu9UQRpm+LzlRxxmK7F0LI6NROM4aJMm1U05SvmNtFKgw5G4p3O4IiR5yCbEuV
vlMaEdT81CHjD6KUGyiqV1vaTytiWViKJapcCgmBBoEqk+WhWzj8CO6fBII6e4BwarMv3sa8vHEu
9B1nq6zJikBL0OztkCr+TKGI6zCUkA3bzLFn2rrYXy0+KxYotNFQhuc/HRggkCQAsEG/1oxkBxzS
FNB1n3yS8JVEa6qdPDgPDAZ+4XcIMqmYJOZDgvHdiHULO1XVq2+2Kc/isdy8EE4iA/1scsxkiW8a
h5llOTYMFWxc5m6P4aO/jhzYUIL5g4T+tCrWgpqU4saalDuz5b5bS1ld7m6TMUgkvOUxEfXtCDWt
HOw3XqJjR4iqC3cWkeh0zkq0EvcME34Kz/NbkRb4fk1TDu5D3pG/ypf0yogNsSiF87Ai60IRok/g
TB7ZH7Ah3hFTPuUswVd+7/k3dxq++pv/8z3Y4xDMSSJQAONcsKNL/OH1rPfYpOgZ1VwtJBDUVkks
R45wLWKFNBjetISQ1O4sXOdMU49z4YGplDtEBbhllzwo9fVymszP9xURoZWszVmWgrHxJtWKgVi5
kNVAQk1TumONWSDPBB8QIhZqZdRRPRjgWb+mn30SDqlgimQp0YwQAOlxRpGtFfkhE1aY4FCC9uTg
kpAipvvu62GY0df/cfAi7N78o/5Y5t5AMhU1JTlCdh8/JKnLAtsbzZv3pJzuamVMOIBiE61ZBQOD
DtrkRjdBL6u/3v1SgM/t520oUSAmgakp2vBpX1GPxrvI0eZc9QOs0fuhIZZvsrkXwfg3vykxL2V/
XZa4WgEFMD9+BUkwN8i6cgXRV8ebRQPZ0npfqTtY9iVYC5yLD/WB5bq3t8vWNr7mkQtdbCUiLXpt
jehPNjGpxf+M3HAr66leHNXYvfDUdQJMWFenBYYii9Im2jp+XG5ddwpEPnggBSl7nQBpaiULnT37
jTb7JESYWJTXtDWmJQfpn7lEr4hEJSIILZTWps/jQ/pfqWKbF/NMzWzWursgP8pOw4wlrN827IG4
G9HpiXynLUgSe6j7Zx+5Bx5O7pdoM5d8iWtxBpQio2gDgZlstqnBJL7JzEJsGj9C/yfFBpaJ0nAG
z8mw2L5Bh5G2kjZGNXjsZ+nL0jJlbUk+evs1zYfbNI0WwgSiskxRk1CNlsa4CRzlGoRnVNnvfhVB
bMxiyl23RsOdlOPYjFbuVUYKSwjbpL9YO7NKw6kAYVx6DTg6bueWYlph9hodif5azjEHMq6Hdrpo
Nf04DmvdmgSmlluyu3Aq64BVO/OZm4LKTuWBsr2WEPp8GCzqNAS9nUJ92xM38ctFKsUd8Fp0CskX
TvDX/P6lRGSZL1XwcCx9U2rZyWvW/3PkqMoQ/zj1zZ3pt55IpcPhq/HA78s2Tt+I88Qy4m1IgdI6
FX+zOuiL40PihuqE8czXYyVmECzpcefcgEEs670Fu0uFBDggMqVEzz2RjT+dc6e6JYsRlQBYI34Z
9mp5E/rMfZDFMrbhsgjdDxAlD9WTT9cb6dYyNlLW/Ioum60e9YngxzQO7rLbgg37MLO6LWGEFJEI
CROuTZEc90+1lpYRwNLF/nKZJFX3AgW5S4Kz8KDMnuyAiW23blkujNtkGXOfe78ayLuctKzcBgl1
mh3Eo+duJs2Fu/BsoCjUBJxn/Rp9AxoWJ/fpQPCA8tJMHhfXsMuFxtvZ5JhQVjfvLiGrZ5fQkhCx
m40abrKtCvOT0JaHNeDTtO9qQM+/RZYtfOGJONFdx5+4+YeLK6/WhXIcEohsnT4Yy+79kwY1iinF
2V1cWKDsPrDACnwdWjrRlYtYocKiKw+7erJBHVa8vMWmBysdg04djr/5K1E8vEBZJ0fL7NXdpxgD
TIn/cCdmNZtN2lfAelwlip6Xwu5LCjFRb+yxN+/Sv5QDefFec+Gom1kfLOzExntD+1Kneu7+KfZZ
fL5RsUcwbnmUXTUNJQLTm5tQ6UPXj41+VE1OLQ2CMhJY7rYjiapqlDqrybcIWqKmu6AGT3yTzlKM
St8pUyxb8fqLoY8xh8tYJvzgR3MYOZSu0pqZNMwdd6y+OxzsiA8pg/V5tHghf6cIrf2a6esE425O
T6qz0W6fdienKHGZWS9+j6O6PfhKkyqhv/ATf1c+GfVpGMR2iN+OpJrEznDtLqAd5T71gHnOeby1
LwJaBRxozH9FcY/zqzlufmbDtuxHBjaLBfehtS6vEL9xnkKqV7fIrER4hRu1Dzu2++Q9XWfcCN1G
yXGPnPUIoKrqO9Lx/9EVimuEf4PfqXMV/OnDEFpWbydO+2d5HoU+X6jn0+SZwhKCIaOtiznGdMRv
gM8yqybSnCCzpyCLZkEKGy+cWEpKPtskPCzL5fxh/ot9ha03UWL2hf+ShY8QeFpReySTISJ00SMR
vMWgM9um55ecBtrt59xyfLFvOUdK2Ms2t1UQ00AgwENdw3Ke17jxfaYEDsTQop3ow3T421MZxtqX
D5tAflrMMUQ+nLE8ae+gbAJJvPobzvHyA4QjzCYkjLrt5PA58+MotFOODgVG4Zr7EO2NrO+SZnL7
xFB+nMPhcFW87AaKgAyaBE93ZpOWK6E9B8xzXUtiPzmXPGi/KGAYGrgvl0e1yY24JGUYWAdrjFIx
t4w/OsZE5sqLabnMZ7wNSZ4Sn3Szz4hmvHrbvCmxwWyMiks14mMqQXcNUbcSDJdy8WJ9c5QfBFN6
KxOttL51l9H9lZP7pTbp+vrF9F14VJobkAfcRUgyiymmOlyDjT6dOOoiSwuRykSzZ9A2Uhr4f038
1rZc4N9XQaVyjVk/3ENVwizx/484ktwInWwIFD0CoBJ3o6PjIGUpljYhQdT6DGt0uoIwjPt933bq
wC0wRdFAbDdcduFziihKeneKlj8p1LiLbjT6Z9r3hR+Jo3B1UVx4W3WUA3p/RzfrE5Q8Afv8PPAi
DiYCQbMrt6PbToTP294kdZlwTku8dEDcaQXi3HR6FkDwWlD/dSVZDActLUXIkbGx/8fCYb6jc0S1
f9vA8yFMvVBVDW5RRz/ucw9pSfYmxuOdRPteSXbZdR5emnJQJVOjgV07ulAuy8ZrSeO2jBKBoJFC
qjnTDdRZDufY29op+zYVqarL1loceDrzpHoBgFazhDLiR7x5CciRtnxQ02TUIUtkH7GYUIMi8m+x
JtDeShw5hSKlKreIA5CvceezUNO9ld3Fg4sGyY6tpaoBTWOG1GsYSu8RkdL8uygoJihxtlTDsHbr
JV4ufvoAvVn/bh0WUFpkcFmTRibY1xxv0lmVIPg2w7nDaxCZnFgJyCGO05HMWdODgDB9pNQ6LAgy
g4/ue2/q6NHrb1p+g3Foknbd8NSSDS7m8OSpDPwejtc/rD55RlrKR7YbOBXYUJCeMKv9kCdqsPK3
bXlDCJ1SMETTBykIYQ6Mr01vujqBmhRXSgfQWM/yiufMZjogk8RDpYhmCaWBA4dbIBueRyyEQAl6
pjiiWxJ+UzLPallaGu9Fifi1Dg9jSxbwuT4/jGG9q84m+d1MuCT1dojzMcqleEJRpJwXuUBlCDJv
x+RPl1lp37w1mpbIGcC6T+bM5r/b6Ydg6ktM9VsLDp9O4juaiOufHRlHMTOAP1v1CtlXV4dOID4m
6o5fB4xFm+q6uTfzRUO/LoyQLMLc+lQej0jimxOdEVo+tLkYcL15f+HK5NGYiIlPFu7vzzizM7Dq
GSPS4RqHp99ZgUdoMCDbtrD9mWU6UUl4iyduNQoX8IBCfrzvIFXC3CK4V/iSwjfH2Bf85h7EIIF6
26rQ/89zEp20tc/syh+gxR8ccj60gHCh/06Zl50juktwYYScLROHGYwxCdf0kN22/Ygjj6eFOasE
VTHk9d4fw0zxlynaUeDRFWEMrbczrdE68jSe+25UvABTkOtFL6SELVe1F35vjT6IQJUdY/KSPtRI
qs30uVDlnMKc7/5q6d9JyN7AbnQf+GYp53P4/pnjjDcOZ6KvbdZz4cYRJnkBoNWX0nWQ3V1Asg1p
cNzrZdJtJZvvFSOAP0/AT5uh+GONTO/8GK9XAtauCU0DkctbVbzNPT9dl/rh354tkW+FDXNwy56u
Jobt2RBXHWo/n4dRWiVSVVdMhPS5SYhGMz/UkDO4/wq00JLjBtLrWSYACl+6d0izVuYE0SMw58c/
+dTl8VFnlUi5XND3JuPPF8Or0Of2Nml0hwAfYpphnf9v1CoVOAs2y1uXQ5uYM9n1P0MDHaGuFpII
7N8EiqTeMBo8XZa9hLw7fpxyY9tbEL7HicVapwnR9hRD0r7/DtoVLHgN+xenfuxR3D7GkE9VH7+B
FV2qjI5RJ0O6G/tDSHT2YbKzbd9WRhAPELqEOj3Eio1d9mQKi5Epzf6BiAvtsKFvyEvhUwwgmSe9
sG+6TenMjWX75cs1NcHt8vn0tnkYcASEWhHGX/rtvhJSP8XS+uWxJhvUN6wpX5Gq2+0hO1Kbaalt
ppb7XCnPcP/G0RXvb1dqzcUeCSXj503EHtvyXa9VQVjWY/5n2a0lntwauzhSqbf/uP5CljPnkH+j
VXF/GfLpVNyhlyLXh6BFAP0j2vDaRo6AFK7rfV472ZborHP+JSjWJXNmE0OGIhiFjyPijb6oMIyK
ZQNf5JrkuNP9AByFCqDQZW+cAwPSAIE7q5fWAVHfk1tg4kIRmS2QRR98r8FRjBdDR8YuPzQ6O45e
z1lRVr9L5fatKchiM6FV2JWqn/tvfMamiTbQwn8W6PsKQUZwvfGg6vPHfDi+BBJDWXSICb3Cdit4
rhdK8Mq3LglKDDk2ZG+JAZG7IA0ziX4DIUGKDCURMWa0NFuQJmiQeLhuTgX1cndKY/KzXkuoUWOR
h3oO2kbyShiVV4cd0zHFXBD9rSwtsJM5K7vgVuMtBn6vnXlD757Jm8/QegqF9FKe7yFC1rjytDwI
ifCDZqyZAmfsXGx8QOfEZgvjA/Hwjpv3DldAW+D07DwyhWxcOjWUkwO0seN8EGR0UjbVymxua4Sg
kN0AHa6aByL/zhvqmjNY+UdIDldVf01PNBW/1t8yRj7CaYspzGC+jW+DzObqQGviEtOXxTNaoLMZ
QiwNu+Whf8gdAUxzME8MNSmxWw/xng0BQCxIDMWSGYjgl/qiX850mcNKjb4tVJeDG3fUHSb2VpBa
zORP1boq55rMbQJfbr6G7mCdpMUUXl7MQtDdbeSrQkkPUSXDl2MdPU7NRRC3E/ANz4dhzFVX0AYA
Siq6YaDxTBE50P43GSUp2tXIjlXm9Bh11UEU9p+vqDUUtk4rEWTZ8H8V0VQ6+NXCeaN2Nhfnmlq9
oHzVtIjAbq/QcewKHhHsk1XlRTrI3NKLD8mzpMGMKKYLy6gHTmqQA8aYJ5QtI9w8fTezL/QuEJee
0I4lmVHtTpc4ciTxpD6l2jpGKZdSGHy9VI/WQ5tm3biJOBvM8pGF93QuOlIuXDGcGgTWMTIywPsy
M9ckjd1M5q+UC72RGPpYmAJA8guqMu0wE8jcU8DZ3Mdg7+lzjA61s0F52xYIiGLZkT0XWbaEAwd5
NptpFkC3ei0O8279GzOu8TY26KJ8mrctkuU8fgqcv6xxdXAydIgI4gomGrel1OJ+9WUtouII9EhG
CBNnONtNWRSHLaeUM5pgS6b8qsKzXKGoh2YsOG8lZe2ESiRfN7PML/oLsTZ4YTFib3tvODSpAEHb
fr3Qr0Mhib8rkM3dIb/uiCIMzRTwbiW4X2rJr0Mf18qBnSV25j2+PXMV7jYSM2dqHh5oB8K7UOOg
MiwAoET54rNI3TcHY7mGvtbxLwmorsB0CAvLH53TShLM+FrA2Flv8ne11gDpyPAAi0JRq/wsaR7M
oazZnWVfHQ9gzWffPcm90q49NELIJtEBX9g3m03E5Yn9nFCvKCxXEk0xoTHxqDz902R63CULeWIb
NCCj+GJr8EfN/P2qaOTm4U762G/0/Qjo0tKuHlZlLl6JEs3Sv1dddrr8OyaNR+ZV8M+gdLmoyjNy
D6H6RTO3tZrIaJkgWjVpjUjaDENmfxmPlC85iGdRmCsgs6bTWBNMg6d1PSb9b0qblgEuaQ601lDa
1ldRUN7hA0+8WTYtLrRjLbYmsTWXrEc9DFSp7ohjEUaBGK3cT99rUc3NEShLng5IgOJwxNU4J1d6
Wshki9gru9CNxis8r4e+li88oBdJVFA9HSevKBfthIW4laOONPhMEodmbwY/kNjzxUbWwySX6N0p
ZpMcCSmYcKPuiSb/ceYQd2Wr/3ftfNuJE/wUwVan6KLmVaoj1d9rfpnq5Nn0+MWbYEvn5F5fwj6A
vEprrV4DaST+QQqi5qNHFJQ2lu8kcz3oafh2V42OPtG6x+u/dI/TDKCJiYmcQSLD8knEfhTO6S0a
JE9Ms81QsR7xTZzdjBfns+SU2d76ioDALbaKU9DzalYxMCa7qO0mqzPB1+UOA0rAsnvJ/dUalIIA
Ia2+H74wzovY7H6wqzifqjrHCi/VrLE6Gmq/EQCD5phxYzrOtZlYPSjttU7ZwF+iWplWXdii1DpU
EnbT63KHzZCbHAJnQVl8y9ik2MyVPHndSsj5VwKKpvflPYBeYSM8D/jtROprGrDPK0oVjKHzbNBV
oaBkslBCpUorHLpUS7JVNbC3tRIArzAgo5pC0R5k4ihnS7hboH/uWmYvCtgp/E44iEoRLuwMNZ8+
gRVCJG8J9AueW55KmHMK/rJNuzwE2xmBN4CbXexa50Y3hdMAxsma6hryqmAiXDVb3QQAz2pAVQjn
rMNuEAyl5tjRb1FLIlqq8y3DcWar9s6DEn16z3QY6Oo6b2MPBBz3spxNQNkFMCd/7arwuJXfj+wX
O4KdjbN7zef6PJX5dal4Fgk64hswVsK3NAA6iLGAI64X3E9JpJZkc/YHRM5sEJZotVlcb9qK12Ph
KT3dUDJVnDGl2kMgEWWL0S7JQ7P1ZQ6yFNFZ3JcuDQG9lHLbDOdl+L/LxM3AC4r1r3niMdfuweDS
jZZkv2xG3NsuzhNL3+KC+yXZkVpupnUkHeHJyXSQpuUZsqNbrrF7+FQdveKWqPaOJY8uRNyLmqNY
ZqDrr4TLn//KWuu+sX7/flymIDSLHNjjF+UDjEIuef5GbqAL+YghIFepUzbsEf1Cecv9v9gneVlp
Dc7x7tSIU0tvNBq74z3dvLgPLG0mb7Lo5VIdulLuHWjTZxgMYkya7Ex8OLMM0fLMV0AOnfFWt6vt
34VlgASoepMDOhMy5QHbjSnUbxRVQcPSzlGQ49gW00zlIPHM7yBgqxhcvKIhH9hSirZuf0wRAKIx
h3Nt3K6MZDwIaPZljid3vgsQJZDacBhK05nBWvrHEpjEXw+QDulctAI1a+f6nPq6gZC5sMvUVtn4
VhNMEozlp23qBgkcgoQpS2OIQSi+PulMVlABft7tKZaHIxot828B3WqzJVn6VeQFaLGIg/IkoLe0
R3X1eYLO+4bTsvIb5vELu9XJYd9ZmRl/pZkAopyxocO7CD/bRzSiP7fgp5RTb861DxtYvh/11L4O
pOwM+ntjVTQgtm1WGcELmmnu3uJMmuQIDdglLJYbCTUk2lAWPV6utGAMuLb6xZz+iEilhKQEAFCT
bbtQyhHaOMInjK26D06wbpwSn1Gm4A5CDoAlF5F8VtuJ6HzYcljDgIViUxigiP8mSAZG4MKso3hb
9x+xy+wQ/MDE3HZkcZ/40kifQuk9N1Zo8c8FIUOXJO7o/so3S+95bk015ZGiEk8z8xkilSsxG1kO
ItRcL1nh7W0tCVTtszFJvmi4azQSN8YZo2K/QlOb8odikDHlEJmvVN4yznBxYmK/wOmmDkDuOja8
phEmSHO+zHDugweD7snDTEfi1mhZbUrdb7/E9Zt3my5tveKT4aXnjfBWBCgPxuWhou1UmD10wEXx
BizKzqUlEtqiEzNSV+NRlzUIX+l3WjqXCQF6zF6LCPTm28AjkFVGoOpJDA0iFqT0nhSOjlNVfQ92
EtpuwEecaDLGBuWIl14tJxMD50BMtAgg2fqrnXEdrPeojhvtHZJI6FWF4FQD3LJ0S68/PEBrzZ13
4LHKFMb0WmmXdXBA7Sj6oxUo6eQsnH54iR0h5Ea4gY9lIhKk3flwScTnOVMsRgEquswXMs85OBtb
1FahVteTVwOR9Dyc9CBkHAqAp4EBRQrVtZanIwNB+AYYq7tRTyPCBMdHy2QLGWkGTGWTQkr6KaAr
y5a9jfGNtW05iU/6pSbRkvqgMHZOSWWpkmAe0P27pHR/YS/RsD8gf/eLtwdmxetb2oSXEIt1xEMo
cuFfTvWbqJe44FFoXmVzGbWG5vSU8lpL8CslZaMkizGFUuEDGSGX+9IaUzfCPnyX9QzYRKySRdeO
7mOd1sX9ZC/ZHTq9+IeD+tBFjs3GqTNMSD7t6iEqipZskQAtMVMeafv83su/go8qxXoSuCwpDAsA
gPDArbA1mM9CnJI+34DdZmx4WvpZS0/ACgnmC0CfPLfDhLmmCCmwthinTKQvU/BvjJOHX88kIwGF
+rGdAps4XbVEkWNJgmpOHfPdJ+HENPDuhSh3iENdWuP8fii3yk9h08aC17snzFDNVGW/BlxIhcT2
QZu4YXN13A0Iu5+vqPzC85YUnxVZTEyO8BsouK2Vc3hvc2UbP105tZ4pGV+798YUbqox9qkt1b/L
9qhMrxuIB8yryHEtXN6NYXN1L6EEbHxV1rU/9LOmSMTLTcLrIaQloKcLpRUnGPUKh/ijDwURmj+C
USO5yufJ3/ygXc+T6r2oJGQvlfhExogYyrce0GDJedKDxYL3ENdi53pQGarMu6xgHE2qc38gXwn3
rsp5PFEdQxN0tMhxFJbXsQpe+SFboC6BfxpBql9AO2gT2aAltNdrllkN4KyQ4g5ug5rOfTnSfWxu
CIt41fSeQa21S2L9UQy/qzdum2PY1lQhP+XcWvhzFLYZXEizsWpahDnxIDcHqiL7nAMSVTjJiYnx
Mk+lA59FajORF+OSdFd/hKI6UnPH0j1bezHLsFqzcQpojjP5surv/b9PdvIlM/wAPujS5duGrNbO
srkJejk/F1ZHpU7HtTawlGjHOGt4yy4zNBbIuFGWdPobyGeap4nFWiDeyOenEMh83jsQnKXwp8rd
WsrLyzL2BcDNLST62+s3gj8GhM26vpxIB7H7FFP7oP8sdOZkAsTc/FQCFww+UIaIKSjtRCoVsIFj
e4lFwocXz/VUpEbpGg/WHAUQJVtJxueFIyZQhSLA9cH/Fg0vwUzx/tnXOpMBCLVmsOUBIT+LoydA
d5pWVqIT8BsKEJADVrMa+3YEO3inJnFmZ7ItWnsVlBostf8/uT0zA4iVMAFj9GYWJWvnc7GMu8VK
KsCMlCcgg4BZyZlIEXPOc1w0sNDimhE6fo951jNxTrUal3o9XEYjzKCGHDhxk/MNvyIlHtAHQVzj
Xr96NKwQQKnaRtpAfr8hr+Dgfrz/JyXBxGzs0W2Jmem+jHD5ICcooSowdmBsUowjRxgQojXuQGRI
qDcumgpe42Nk3L44nYoAkf2pBabbKMIqIMZbBkqxAfS0ezbNZJAnFuUUjbA8XUbUfC5dV2SoOT7b
KTccY5236BB2L0gfoNvQqxRPCs+mBL8Gx6SadZDpSkxWi0Ie5rpZEwzcjzvefZ9g+GTudJXaF1aQ
+zNuyZIBt16IE7BbRDpDdOE9jWKjjbARtN2/qboGd0w12tWC284jCBQj7gyANPzrnwFCj4EEVwPm
4tE68SivfxL4hpAh7J8RnsKQcg/Y70edD0NXUZEdh9cl1pKQ2OiE0teDfHcDEpvLGoHfuW8kUQ9V
r/CPIXyhXl7TVJw0mm4tEgtkfQrz2UTudqd48MKfELOhcAP6zV3kPeM/3Iaub8uGKavJqF6Ji+5a
riovqujmsMGHjXVPEaoTCS/GfIQo0nr0vzEL+E6ZhT6LC/Efh5WAHfric7V2Lkt0mkcaJhboGCo8
XVnXWZOUHzYCjcIQNxme7OfI0JLANqiSimSnWpd7LXMZ7wn/glMS+9ADpfKYvATFnFh6RvEcdWG6
OHn9WoQBsCBRtkw4VPzPXOa+TtyFsWqYgldR4hlgrfFVf+XCTThYdWsg07RqNJODdnx2aRCkqQKz
MiLi4rKs2HHUkRFZMIEf6bWncyAs5G17ip0TkZ9zpJHlK4WAGH6a9y8vB4BwAZBqfs6VBE5CDQzL
TAsJSgAYDVeW6ig1bFsMPts0jruN/BoAz8g++30KxaFzo7WqaR/I041MFCMtmR8CCrvktLzbowkT
X6Lj1MM1+DfSHr70PKivi/EDh/9bc/GguNJsJ6/LclYrzcr0XGkUhyYF6ye8QsNjgzQZGbWja0n7
lKpGM8uygHV1AHCz0gt52o6sml3KSjeAXcXhBOTWEqF8L48Rf2o6sW7bR92w2RN0a/M4yTQttKgf
7ci5Wp5lkjFf6Q2L11kmE1okpHmG6AncpOys0IGpC50Cde9YCrsRW71roMVR3MrA26bYLSwDv8Fr
+5jpN5n33xpy2pxuhsnvmpCv9hbqLVV29YZoAWsEgKpgwbp2d1dZw/XaGfgPrQ0etXVG9lpCkR3i
ahxnAMnbinAwf/ZaGfyaz0yO31hf5Mof8nMv6d51wDNihvN5JUkMwiTMncygx5QGKY3/r4oGGCOn
6oh/N9YyCaroRCF/3Lff7W9nBgktHhrOd6o67La+505v2l69wv9e6SGFaCZdxDlj1lTVMCDPu5RZ
5K28UhSZ2dEmPDGdbEpLij6wYaEmwV1mlWwbZHVaCol+YT3NSZaK+Y1IvA9xQQJCnHgZERGtpCIY
MMREkTHfmECyWjCDat6RDr24CeTsaPfwZ1GvPUcWuRvgreaHUI7wus548KyzCSlleGB1wypwNhkN
0VVW2KZgXsVgTOk9WVrTvCYGkU87O8lYLdRKT1egD9Hs62jF9ksu7rfNfjmUPjWDkhmyntc0evom
2P8l/plYgkhwwHmam9Mf2QdONZppIlZOzqP8RHR3NbCCx4csbDydWipT7B8HTcJZ0OVY/35bucBd
2nw7IZy5jHg1bqM2/CTRHwcAvAKweHICQZZ7OrV/CEArVEK0dZmUPPIgBOcvZxi0DdFy7Ug13WMB
UacaAKrCHch++zdHe3liQuBnTJUnS9Wi2gj2dHmnCr3yL5GqflVo+HhlUX9PrUUxy3vpNWBiStBO
X5WM3WppMLh5ZCzWR4meOm0rF1MmVwKlXabQtoGrz4+3zLK73fN/tM284RGFqv/eYsfqOY0J/8ND
T58KdLLVp/mPAq4Mcke7RsBAfZ87KRJqbEeybgklcgnj5WLfyebvKkX3SEy/A2rYhvLi6TkVsTZT
VY36i86bTMtfcPp/31XnbRf2suqCsuELyZ7/MR/tYfsiuWnLlnCbD90RGeUtpsf5TlzUxtxDC+tR
Lps4a0fjEpNk01NhoQ+ddXa2U5/oT/LvYJSMgyMbFbB8W/5Cq+Ozl95jhbtGCx/yGq/gT8CsWsYS
TFsWN+OPT4aeSMofYxFsaHaupmrVCciqsTwMGAUF/FKWVJyjLasUAe42Mg/2unxBck9uFJKM6vaD
zNi7kkrcuW1B4wNf79nYHJx10nLj6GOAWoRCy6IFdOUzfpi/T7OZ1DjGoVk2nQYbqgvc8uelezim
NeOt4PmGll9XXJjq4w7IRol9eOj3IYhPpnvXaZrOcQv68/p+mFAzMGhT8ukbp/W/UViWbRgDb+U3
V5vgpEBcm14rgrOHTs7XSb5bNn2TO1xblqxgM4BngVelh9v6HnxI0siHGu6w3z74doN1fK2mZKHC
JSh4jn2bIz+8f1jp3pO3f7ls5rGa8616w3eBaI/sA0WkdqE2fWcGUrQ8lJQ4pLaeC4apNHwCNGT1
lhb18pW6KQN4UuWlRIuRlS/DraD5SOT1D56aKLYT61fMxvFHyvdF28GnX2PWTh7L+WnA5n0d1nfv
Pnp7yhc/52qMODYzWdEwVKEcBT2/GWPk4mVtYMdYTRXH/jD5Q73SPLeIGsYrdDh00PnF9QvojRjp
CsPnXldaYafPvs7c/ADpNwBMNGIt/P5ceUrA+WAE71BnPbksFzYDxinnv+j0tP5NfQMeUGX4xl6P
OHrO8Gx4/gHIbzONBYp2dzFNuZhDzUfbzj3Z76QhzMk6O703RM6bbAtewGTninGYFF9isuc2yeAk
vU9yxNiMr8PfBL3iEcxWfBqrQ/LCmPch3l2HsZ5n3eIbDv/kH39cV6a9sY+6IoJD3iIt99kXb+e1
I9Bp/tXkHnxyNZbFogOJGQ/mMpT/jFnYDxSOSRqK2p0P6vz2AnU6g5+AwbfiQyiplCZeeIN9upZB
fGswXWTbQCLiFcyKL+SCcfh0ZzW7H3RnQqK7djEQEwa2iWy3U94BfUL/cq36BsD8c0MO+Ufd0jMm
mMlkYfGR5AiInzHE2MPCcv9/BTLH4aFHF4JPnhCvxUxwnPZvA5BpyUBVchAs0+XO+USHHsfHVGpW
5FciiCqEBf91SA14OIQdUYAYqyl6UeKwHtHQXm37bjUQCaS8lyB3SfpS81WHKi4axzgoxMVhCNBX
DUjyWVUPMZ2ZQeKS75v4GSKZGyedlBtWwNPHuQefekQx/o95fvgpHmUG0Gpp4/gkAOnbPtFNVsG+
zNn+vNpI5Ccr0ynym2Poz1y47Fq8mf7fbbcI/qRxu6i7/GNnABEEE5l1e6KCEVBnPnK9GXRAjznL
ODt7GZD7AcYiLh0NQlujgqua7zbEB63XMs93pfHmGudv/V8muTtdD/qsbzy4xNGS0y53mKHbsrAA
oSe7jYMaZpURSpXiTbjgM263zSpsOgp+KHC28JWWVO3uFyI8V/FdEHeXG6P9DzT9W/JEEs9jj+Nt
/eu7w9wzTvCFBpMOHVMphyaPLjR2TFYLZVgEe/arVmtsuVBHic1yVkFkbpjvqUpmIzF4XpFN6yrW
RkxYDeMT7Nlpfy5cxrJ8iUV8RUsD1nAQ2pjbgDE8mfYrFbQUhH/BxLxlyKb9fECBTeRa8w3sjm/n
ePTSmiIzLGgaKu8wGojy6nSHXznSNSfGDeR87HkFO9DMSp/5zMt1Btk/40BQH2nw809KWDVbnUn7
f1GddLGLeYI3M5Jdoc8/73pqUy7rtKIs7ZgyQ1bXT1fPahik6KdDC6RjuxRApiuHAIXQSYOkb80o
BlKNKwCZHt5gRDtmsoTHvVHQCsokct4EuiOzzDitCaP8aedje/nl3QrBfPnQkZ2Qce9PjxQUQ209
7MwHFFtWx8l70SZW4Q890Hxi1D4FT1DWAHeZCwD8iFxJnG+sUuB2mtK+askig3eZGkM4ZZGMBcW9
LyS471+KXYfrjDZMETPdhhC6p8yURQ2LO0mPqbMc1Sx05r7lE6VqJDOiD7+l9E/XT2h0rJKdUlo8
G/VsnuIQ63oJ8uP4qoO4aPRDrbXt8uC69u9WmurC/yDKlsEUVJxjYs7osDaHys9Lt6yJwvLWQUXc
6gjiR8Bu8wbG9Y8DzVrknpSHZaQriHrhTfPYGnI/04qepD/45gZoqQ9fW1NORSm0yzdNUOQUuLrt
+YkXEbrWDtbdnwU7TLX+k++v8HgdD/mQYaKXuKmxVSlHVE0Nrb+jJlC62fF/HAWTd3jHntcDjJMQ
gUvv+u2xCwcAC+lp0FdEnZh1zWxj10nr5OPhOdRh31XEZfszThvj4XGrHsUAT9qgphZ4viVRSqT3
V8EvFX0d1m++QyaZM+D8ci15d8qSCTNsBEFY2hJKR5lo2IAQTDv8ISSVSmh9cO8JCy41yjNW9g2F
kYWAYrNrCGcRzRSusQV75J1ueRWroCS1oHeaSBAb63w9q3s4H0XBCRhnpNoEpvblS+5jE1T/gcAy
EFDfC7wun/0+NjNjXpDdq3M687L50i4xpQzrpCzAyUL89Dza8kMEwxSzwbgujq22e7KVXlZZdkfe
+OsGjPpZYxe2C3pCHZJaJr5pRQq5a9kE+UNh75PiW4ELRUYU4t6Y9Zt4NMxfwiKQA3bPyLibA2Mw
5uJKRjspSwf21V+gQwyGl7UnPlbmoq3b8ZRcs5j/z23xxX4ssfwUw/25BPK1G3M22W+ShnrwhnYk
B8CTk83AUZ7Z5P82czJo98BytWqeUM+qvAm9F7xFsuaGBcn1n++S7mkQbi2x3sS8ayTkE6oNhjCi
WVxiPF/qLisWcmpHbufkPNL7Kk9hi3NF7Jo+30CzGqy0XawslpEr383jp5TefSiVGoK9NTtwDbmr
Ayj66iPyeTsH3M/ciDStMk9kijT92GUiHEDoj/6TtQGXB+L72JGmJbQhkchLi6qrA36ykQy+uT4E
nxfiziFerIkOzTJIghJu9EMFXd7GErH35trKnkfygnvUG7gcXFux6fu1Wr8BAE5364SCKJ+DlGO4
J71sLk10hw00nfIJOcbXJx2Ae2GbwE8NXlfzcCRpVw3h04JlFiuxYEnxqd61dBJ0DcK72kOLypx0
vTTfmVXUyJmU7msr31ESEXuAVZxy5LkvhRq85JQSHeK1leWWmvV1dJI7k4+VHr2K2GZG//Yvp9Np
fxxxLi70x+OGzMwiZhpBi3dBpSf/pAxBwtAFpvGUiQcOuwfO/IWgk7iLLZIjmpobi8HkHdKaiOJw
H5GS+MVW1zTC4rwlgf2T5oJ5YAJ52Zpe4FBLUCeuqniHdimMxEfyHFNltJPA/nqITU2g6KRfK3ep
4M824R53lLln9yIOhhH/dhfLPRyrvylOwysmZqKXZHPS1SQQDjJMcfQiniZeUxVrjjBgEet4FimL
qpuStZoGr4VQtLYcqWhQpACYxlnRuqXrZUPeG/uijQjQbnw3GF+LMj30A2DPOuX/mZdVtAYfmk85
jZ21df7yEn/5l40TW6ZWFwzl/IcvkL4F25bJ2QW98Zfu8qI6KagSj0UKdQvY5qb6F+G8D+TXInMN
sGHvaN2g0UplmI8ReHXDeA+GSPco/lpWYQcnoowkwA2lO5Lk1rBzMdv15LmR1EAtZMxvl7op+CLn
CO2g9t67wOzuXP/T0TBYh9db3uHI340rOZz2sDYFOb2RZPAlYJpOPYTz8knFT2QD1jiee4mW7jIr
tpfPAA51xxeLnPB1of1179xBLZlvd2oBbL/Mz056fRKeo6Fhb/NARjIFMhQHWswKOAMXRRvi7T0l
KRYchmZUE77ytgkJeGU/PkeEkCGJW6IRxQt/kiaXV2iouxIgE1T6gbg9IeazbAsozNvz4KvSdTDM
a2IFRb2yAa4o8PAPuKFFvgvmmEZdMNqxDivqFa+E5uEg+COYugXYccCD6PhbDllZSqko5BnaRkxH
AvfwkUC5ZzaPTuCG4rFLI/BpcFqhEPXb85wG31+MuSXdfis8z3BD5u1ZE2TsolG2dlkXTCj56Q1s
zt4kgJKernu3GQcwgYbQwdBauB8TnPkAbXe7UdPLrKkgolE0UfVbaj87uwB7+2q8SG2h8xXzFPUu
lJmZQ0b1KIa9T0hw5rqJEgrpipzjX/uWrI+XWRnqFpWRpuJOCdq3oc2Nqd2CtQ5hSdj54ybWjIyJ
6O27wOOKOmjkak5mdWy8J/rUpH+QT0LiZJHEHwIexITtaMPTIaD8zeXnyLC1qcAtVQjVAvfMAIZZ
4iKivo7xb25cLvvOAO6Vw2eQL18KNOyg6cANUmiU8TsxI//nUahlP8+tIAVlc1nlLKXqQxQkc6Ag
+XjqjzTnxB+qIBC6P4E52Dw99KwR2AP8M5lp8AseJcapE1d8z/kGaB6Dsqs2eL6GWha9G0izO4CG
TPUj77u2mKhYnqJkGIhOnxFISSCKdWOpBC2/U/YE0lUXs7WXFR9DuXsOasRLC3Q8QAZ+EvpLX7CS
yCBJVkGU1cUIeX0ZD4QRwC5z5Dvm0NUkBF5rC+FIRw7jCC9XiDq0BYLrmzik/FyfGZVkzgQTgiqV
CQV3YMnm6sk9ZHJWorsBeRoEMu7yjqYn1KzZUUj3iyMyJXAJDs73XOy5bGU0dt5+uZhemiYpvacP
bBYgaQ5vaODONbpcpfr9KGQQAIqDDplax1vT0kyl/raMX7k3xyWGTApajLzXxe0wqxJp7vP6rz/+
o9mzgtBYUGavAkRvaNcBk/E9qCR3WhIPrlaa8OyJxU+DRCuj0DN/62nhlAZ8T/6Xr3hvmxtxAWvp
2p5H4F/ZyGTN/GoW9KxyUOtd4NS9BmqHsLfJ4qElWPZJzvAg0WWCquL9doSgLpfD4hydVIoH28kk
Vcwl5mdR4iTLuYwax9vPr29VRDhkF/sKkvF+TRXpycyg/aLz3V+p89qI4+AYBsUfW7w/e1KM+7pa
kiQFTBc6ANrAwwInwKV+9zons7WmaTVYGz8y+FWf7oGWL0xdOSA0Dq688ETcfF8CbaQzabMPDfdN
EBOla4F3uKX68FIuj2fSGqSf3gk/ErOQyzVhyJulDzS+RueDzre9fiFT3NZMYt9x0awArAHth5QK
8LENs5XgJVxaYuClOauKGhn52xpEddFaD6pTs1PrWpz04GcNCdZslvkpSgS8UEbBBKwlEsjFoMN+
9SC6rV7zQig2yMRH4MzPdVE8l9OFOy8xSS6LcXysc+Twav6QH1uzAUYy1s6K4rq2KoISR0kl5slx
ASKOqa5n6pM8cUcinCdGS5p7XtOpaY9R+UpeIgH1jaIiZ3vMy7XYJehpvo+8so/6ImJXRSb9H4Q6
yi+yqFrDZCSxpHKb718PgwqMdrOb2EP4ukqdf97nJsdeyRWoAols5bH9s8VN8PtOZHirRAETyH2h
upSiK8ZCRCU5IXzdO32WbT0BHQlqYk7qPr16nbc2mK9phEPW34cf43ErwVgmHinjhENv/K4d8+0O
mu4P3j1JVGkijJG7ixIWgF03dbbFTwziIqakGaRqlpDvKtOxiBagXfpWd6sDw5KQDvmVp6hvFpJP
RW3Tc7f8yeDRFbiYyjamIA7+JMVYLTOGThWJ72cq/e/a3sGjcYwFkewjQs9dQCxwnNI5xgCwxWK6
20UuJL2lYIWfoTWQbIETgBbVWofZGh4SQ1pV+sNPWj39OlqIqGBQ8nE2hvP0mXAVN+NSbJ/V+kJs
nNWPuvP/rc95AMAH53iYCxD3iXUQY8nSTrXTWn23SVXr0V562f6QHBEMsYWlWfn+bI0c1DHrnOzJ
Muu9a2JSYI6ov6NygRHLl47NrLsfBxEl6wm9bmk2AiVn+alYVHqy+ZJk56jUle7fxmNzqflYJJAu
pfqNfs3AEc6h+rANlCqFZ4UjsUBr+27e8Ee3sIAwg4+0ZJfjIO/zh0hK//DKjKwjngQTclJUEnpd
dHRbYaJ2UHBFWydfFKw920a7tFeMfO3vFJIghTOsEfbN8wJY/87MRCr0rKgzvxAA5IDvQ3nDQME0
wYiGk78abrkDSSlXCJCmTrT4FWa8YOmImEsqHLrq+LgI+Z4QcYXCj67cqEKbmSy6u6c1+3QAHzd3
p8M51jx5Q2qfUvIHClVS/00UY74GIbSU3/HLg6i2v7VyibW4/hck4oIoyykkzpikyv2EXVha7+hP
KaP0POBogLgySU512GAQUdH3xKglvyWLyWIJ0rtRWEVVoKYpW0BewmFCLVQylccYEbYnl1v3oAqU
U81pkoV1t/h4Sfie81LQ9b+rzthbzQWwQ1OH2qdCU6BVcuu7QN6ejTKhvSomp9QmNDeFPIaoTdGd
m73JrLc1mAAxYdQUD9LaTm+dmgwAEwp3lNhyd2sW13325TTuonp2eHTV9dcBAUkNUNlKFmE6SWeO
C0GdiKAOH4VgUFYoyhQpoDo4dQxYLX7WdhCqMOCj+oSif0zXwoE0qxtly6h6BqrPxE3e1kNqATgp
R9iPnKUw7trGhVkje5zBVYp+gDlMI4FQfkNw+sa7uJfLT6R25L2kytzqh98CHYeuel2R/HyMMwhP
A45TD2jRXSwTpl/Z3mvDxuI1yMvN2S6yvJzJkI9tBur3kHhVWmOwtkF3REOxyfkFnQDVFCGFsHRh
eJ7IwVPEnkVY7zZpZ/fnnOCbvGERrV0E3JLFAmW8pLRuKMmVIRGfi/567WbEjLkAFejLy8Cwpk3t
ZbOawLobjtzYUSW/1/AZpKwc6tmipcvy3LlLTG23aKz9IP8HJeQF4RVazk6T2gvaxSvvWBAdmsoV
6oBNJB+/L4F7JN85Y21OTBIBb8qYCF7Gpa0ZUwcFG4N9FlAxmOfNUTPEzFl5ALhMqoyw5AQ9rjmr
CyJG3+b9wx0P/lZd961DP9v8PO3Egvm7J/vlSEZ9OknQQq7KMMdD4O+Ck5ik3Rmlr+dhwRrxs8f5
NIN2VywiOczNPcgUDA8ucTQoqIoaJ3dsNx3T45ojRUtUTVzya39dTIycxbX0eydJfnLlVMMZ7mSw
TiIRUsHtJJ6uMoeR8wKUVAoJTEJM8oY9dYr1bp8OvkdsDUOsvXJ6IvngeKSy3ARAwvf+sniaUSa4
d/MeGF/saArs2eBBbMRkujlCtY1z+waobduI8b1N+ByQFqft6KoO6Y/PGKoD+d2wqRV+oAvGv4MF
wTA3QQf/e8LCjKMxT2RpSE5vNpCD1RRmIiTT0bsChGMFoCNhJyj/35bD4+3ausfN6ysuVZExGPGa
1Y3vKn77A3aycDiwioYiptQpZVID4nKEPn5sqW27Enad2ohWMZdVnF3gejv9NlUS3rJTLQnJA/3l
neTnvjnkGKGYfTsNdEHSWIQn/tdVy9KlHODMvK7vAH4CuEGwSuibRuGIp4UwD1cri5qxvMhF9PWi
Rk0eTOxTIv1u7NA1olVndKrEiK4BLcKPWswNPVGeBFeoWPI9p66RhVHhwMlenDNOjdmKdBJuNmtT
bPIF5I64kn5hPmlwzA2dxU68UGnH3fULuXnmfROmS05gXiHd4hm2pXJtLlev9EW8EIDshDjLnAV3
NddyXgK34oVfYwq5hArRrfKEoBVFQtrd1SmLp27s3z2B3z/6Z4fDMBZtz9ufZxAQA7K+nJzXDWr6
nyRl8yNCQkDD2YgG5qx+0jee5sfbbumlzYvw8wPlre/W/cPnBdZ08q7PWpJDovpQsKvNJBs7Sm6z
ei4roJE7uwKTn+ZWkzT68RiLUwb/FQSou41IyCGijLKrsM9V1HZmaocDxTLROyKYkS9fAae7z7Cy
bpg/wGKSZVBZfj096C9OumuFtwzw0xQn43/cLNl2IPysW03U93zQbMQ26vHunzc36njOW5udB31N
1G5OAeimehXJmsY2eSbw8GckVIEgVULzq2LLZbstVcME6bliP4+yPOUsawurqtuYRTnuyrOHLT5x
rFbUJ62xCMlgMIYZnEpUmmtKuRWx3ahT2QvmY065l4ySxz1zFv+M0X0Sbfy5HlrYIe8spzvdtMpe
dhdY3eAVnSExuPYXeX6qMViXbkKy1XbWQiFp8Z3psl5wBwQq4F7Azi2aVngRaC8ObL2+77cpCubc
N/jLpDumdfvopwFPhh4iyPZAdkMQcbhuFuUIutY2WDVS9Mv//aIvqgl1PuhX6BQqoY18qkBNHw40
98emiUQgfLT41836hSJc/x8TXGhrOlblkmeOdX6oXhREFM9IVw9wQ54ciZOkBij0CPZuRNVurFHc
H63zrCguDqdxY8Fp+krzUmvME7XAkUIEnExB5G720Wdd/LQrP9dUg6vN31nEueWwNPsj7v4qvkdc
/nCeBEbyeL5JyrM8oSIfzaHR2rlbFOrRd5W88+zkr8XXoWt3gozqujJK5JrGk2rI95vrNbQ9ZiMA
VnNj2QYC6rF9hlgJHwfdnkGvNaPw1lGp/Jx4Ng2DEK2Z+DVGgsUfbeJKLehdzQrPAPJVFHWj3Vsx
kb7OndY8SxQcc1Oas3oHyHftlBqtj+kRRGZfhwI9Sa/vmDSpGG8Qq5Rcw1tOBb9JO25elvQ1hfC6
bkGqIrXX6rWhDoSJiqMh2wcfsxI1+p//e9DysBRAGkA38RmBS7dv0yLjpNaafU8PBjw68+wI/nVp
woXGYyE370yFO7oIyJqFhUC/VUEQU5uCwZMRGvSnN0QVH+BKPpJoii4YsxE+bPKrNUg8RRjlQav0
bRW3R9HaOqJIuQS3Ogrso3pyLgcVN90XpmQoFVEhMvWIEttL+FJzVrE3Ux2FhMzrVQrZe5D3Jtmd
rkKlZ7d4GskEtB6jvDwyIqiThxAtlSWDihufD5XTxcMc5U3RYa5N9BChfBz+wTJItinvSdOr65e/
E9KwMCfkoXJcfzVgA08lREpr+d/61sSEQXC9tBL0+o72e/f2KvZk7veBJQLaIs1Q5iZip/s2MeB8
Q2Y6o1N+V1jtqCPLzwM823mkLNw/Zen7dNSe4C8rwB43k6Arw+P1C9ui5K5PaIS+rz0V0ZRdDqtt
+dFa0X9C4Re2YXBv+GG2p97fDGHBTLEoN+jcCwnz63ONdJVTxMwWyDP69jWo2V41oix4wCgPg/Nk
3GG8n4VakiyPLNsdb11VivwZGx7oqOOCGSVRhBSo5Pme82fildKl6XByKp2CigF9Ezt3AmDNcTvx
K3gG76RkwZE4Wu2gn8wNvs4xiCtuVzK3XejqvY4+wBtPYmn/5QMhTznSoF8NtKYlKZdqsuG3u+5S
SIAl5pGSgwfPtEgr3ih/vfxzgJU7wHzTlU65jToN2bHq5oG5MgR3FaJuSqKqEbNP3Usma18aIZQ+
Ux7zu+bsJEfBfxIR8waFZWAHlyaSJNKh6IUxIV83QzdG5zrM/0AxXiVNiypAn4BTnbbtmTOicw3H
/uLkp4dRX1Uw9XIZqhxDGK4wnL5tXzF3EpX1xkLtYcsIn8b8M6HAoioYgh52cj8Y5xF4mKKAHphi
9QsuNRhvKmX63QSTyWOvcEep18YEGLq3wgh9Y70AKVODe1UcHjtXLefFuiYLvGwQmncCFRmC48K1
+qq0GG7sicFs8LUF98AIcK36xqNfff6gAnXWq2AmwinHdnSNbWLMw6HnT8ERKIjsZ3NwcSbXWgKY
9NADcgvqdpoLpKt0+J31wogQ62QUZDk/o4RFfHdEc4oEC2Cm/83E0eVRldpwDiS9dVh/C1lqrs2P
JG0Zps1acxYJHyLnqhgZ/ClKRVje+mOWT3JPpYqOBX5ouAGXyu0v0TTL6uo7UGIneg6ikqBIeVvd
FhPHs+k5GgPzxtI5WTPnBq+iCjbdL9C4d2iVwCMW7HX9kmncxnGIuaXY4VQ7xR0DTUcLbJNG5JcL
aIpQo3HFeg5u4x/CI0PMqtHH4zQaOoFgryY5gHU1x8mnAgrMtFAuomir09LzvMNxe4r3tP3PzROs
MCoxTOIDL2lZuR79RU5THJnyLwwqBiNXN5kFig7n5ya4NrBL63SwsqsnehES4q5Nzx+lM7xpRiK8
heSlJ+ksKR5tspUvuWvo/XynIx86h4GTcbGkwFL/G8e8RiQtEvFXPzTkcHoszllUv3PwvRtjbGYL
G95z1jGT2OGzsMFkrkCQEpQXUpDQSSAkQ1BXSp/tjgfsIKyTZ6zO/AJyAEXAscHxXWfgkzXsl3Pm
t9eD7jT2dMH4JC1hvFkd/RlMvhnuQD+KisftbnIHLd/779S+VMdOrJFdQdmOsT5cb+Dp8pA2pnHT
lQcy/6zSEnby2Yafn6ml8VjGYFMyrirPNAQsJs2Xx+VlvXyTsjP2QHeludLL/W5wMwGxA9C3ADkW
GcVuymS9gbu7Z5xPonwzmx7CqAgjZCq2gZRQjkM/sTEFsAS9FkADFXKiq2hhvczGLvdwtdWaz/u+
fJZ4dcU4Pi4CG+Zjc2tJBTOW+Ls5XYAf9/0IaAogCn/dhnfDBDD12BH6hHgHJc2+OvG14xTmmLE/
gEmwz0DDdVdiwJafQW2O/mhyHaL7i7NIv/BArGAoA8jQ/EV8UgnwqyAHRlfRaBxWRzgJ9l8ghMUp
3rkx/H9VzR/9yIc5Oxys4Ca7hJYIM2xgl8NVFeK1tUDt3pXewAuFLZD6JJhvkMdTdywqrHuw6ZLx
0RUfd0GSpGAEwPeCmlZbdqY4Uy6cCIGDFECg+obLfEI2urvAFC5ciBM59taxl8RcaU1n6SfRlYCT
hVQ4fuNrHlsS7e2IOL5+XNbcMXQoqdX794HuIzjglfFJu1AvYJFS+HiKrQrwR0TzHpZYqkfoTn9s
X7Hiz8oPvBcAatfFnAzLbLRWt4YaOr2fwhLDXApbfSHYQNAsA/Np2/fAtnpBMz/13Hl/O7JVwQwI
vGvkZn4W6pkJTHbO98Nri5hF8uR6iNbEza5n09d8p7DqkhsSEKXe0vhoyxUnTTpmDm48Ezx5Nn0o
U+Ws/Z6wymtzk4Armg5bNDT4MLJeDsExpRaupWanmctEWmbNZ407XN44l6bofVAP4Xt+t6gt14c0
wRPIPBGHs5bLGWpBa+AlJ2FG87vJeArFXsTJ6uCcBuYh8aYgYgdpnBdGQrJ9qLSD3wlQvEmdk2lm
kmIfZHfWd4kW10Ucf3aU+TBB/2pVrfrmDALrHpXWZ03iXmQ02tovDgKYFmCsW6VGmwWg27B3mmap
wZMyUe+X5aEMCabkrAIzDm4ZIWVRASBPU2U29jHmzYBJBhK5STbwrDwKUcxTnb2dQx6G9VACP862
sVBnqN9p1dXMe5fgZhDMIZL7JkNsqwf5Ss3S75d67R4sRc02WjxuzCm9znnfv8GHX3K+QFhSxVC1
tPTbwonRYxu/mHEq+UXAA/v1kWPs/UfLRRp4MWTwFBzOeAUkUuyKKUWli+W8fjv3FvCH/u7uxGP6
1nF2fNrONqN0Mwg4O631BJ8dnAo3pejPU1gl13ISxiaZAQJ6pMM1w6FvMCEftpBK6grHnzqs/YEQ
cyd4rOKCwKTw+kRDLkwiI4ZYeCZbxmoAlCUFHPA2Q5CduqisGZPU5Sa3joe+XjdKCjApcOfzkBMq
ciOF7WrX9SuG/m1XIdDGR8GKK2CcbME7Ind4KYzJ/BJFwZ5Pqsgb5Hxe+mmZicMh3eHbbdJVWudo
3IuaMc/xBpl0+OIEj25cw+NkRdsgrVuvaNACCZ3+lHcGvYfjh2V9ZnjvwrAwBMqinr5oXUpG1FNt
DnzyMDelYvhL3tNWRm38HpiEqegJv0oR+GTrdktNKqVAIztjT5wHQRbNIlJpoRqOZ7nQMVnRwNBH
roM+fZ3jslC6/dZCrWa5m7evK7kUqsajYqnNOt27Wm333o23hpvWf+Skerfdk1VMEzfLz7MrwQUX
Wch5l7gZxSJUFQDb19Z1UoMm2UwQp/BHQEMO4isMfArJPMrFKGvpYnyQ292UClW9SHWJWD+k25Eq
PuVaFeQ9uDTTu1GmstymGtJb3DZe5zc4kF8TqX+mxVYt8p03Uw3d3qZ67lGr6jK3ue2/JOeCg5iv
b9msB9FqgrMO6+R2iLHcfkCPjbnuj3DlECaEbktpEcmr1OueIiDnsMy/hwOAsdGbC2h0D14xzwO2
+fD6i9GD9QEDostAl5PtAB8BsUMj8+CiqQB2SYQBu1bc5rclYU359ASVlMa8eRtUUg6En3zbJj1X
UDMQFJ78dFkqHQNwzvrnSJf5/tpb0k7l9BIzR+0oZGF0I5JqWQggzAnoDfJg2SG92x+/Ow/BZ9M2
JG9pjah1GxY4ZEcO1DLdqyCTQCRj4XHzbCiotEFq7HvsbewVdLOEebnn6HkYJvNTUPDDhpjglmYk
DqLJC4Mu9rP0lahLstIX1mbxWgfvzhJ3tzFJMSpBBu9dnFTYFufHhCBYo2IWDeDyfaFHUmORbh/D
ryK3VwhNy1SWahfKAuR1IZaogrIA3q+F/Kl0CR+p0CxqFLKWZxbfpzVYZVumPMCvZT1OkezyjEs8
tOd+cFPJAFczejkL251Wnk9CxmkQYmiVBhAkf45DulSvDTJKEmJp2spIsL+Tiy/rumeX6Y6AE0tk
rvgs7WQ99DV4dzeBJNriHcaztYkD3xMAhteH1PIm4n+cwYZQlksLWZmKwoHECudVxJbLRlSJZh+U
Ng7O95qcWsvkYYlGRU1nxAnuV9FmZoEYIiHiCfvC506ER68Znn3pNJqc8dcuVq/jfdSPBWs9Jgcv
V49MeYzFHyQausW/8HAB6V2jDMgPhbZ9r7xjsIs+T79UaYca6eTLPfsD325Js+XXK/U45rlb5pEK
HbkKnEwd9SSJukfB7feVO8EX16sIpgRw8mxHpZ6/bJuYwyUeRygxuLZOnn6B9fdKa5omhXyyhG4X
WGnVHRQi+7oUTR1tq/isxFccC8Iasrza+HQibEvDzSbjYDq9CxvCP0x+v3SaevQI/l/x4ccnUr74
WCYmzQkXi0wosjI0+P0jzk9kRtD5D3g1qZ3q1BFA8NcnZC28cHuYmSvNmCIzPVldYJ1dk4sEFCqA
vxgJYOvco9mLAOXgYCmmLuvYX+bNe/oyMhwbA50pbOKZ6k5o55jSLu66kb12LuectoN8e6Lu/vqc
Qm4AA9WMB9tNaTLkkYYIoBJ1h88thYsAOcX6EE4ZL6wmsBtK+Mtc9EeBY84J5MHPP8tO6OVD2v3N
8x7+HVM5B39B1nzw4FwvmFW3a7wqcBblegJ84+1D1qqmgLWlwTUYbxYJfOptRVEKAcsZFS5g4x7M
Vjwoc0f4NAWhw1NEW2p8wheG8bkRbNCF9uRxBKFhFAR2aJ40vX3tau8+S/xKeCcHxg2F638ZvDMN
cIpqdnB1Iy2DYsfhcEICqjsfPQF6nF37GjbY/R0e40GJKZLXgscqYw6WI0S2zi3jqK17gXZFm/2c
20BC/DcEEIKrAoQPvT5qujCM8rpcJ1H9sdJ1YWOBWb9N+kEznVpyvKx1lunzQrlKaWsYsXZZnl59
wpu/w1Yp0n7hfWGYh6ndnCM9K9XV3V3BrwESsc1tUMzGMWPiBB5eGE1HIv9ATkV7hNshOFxxdC3o
R5P1GDzDtuwzUWGfeRvt0N9I+0WgB+gaKEMZDSsIp3enr3u3r9TLJ31jgPkJwa9Z2J5Z44WmSwGr
Y47pkFYFj9vt9DHfCpb3cPNjcKSerXUXeEECes7Dh6B8EJafNXnfQLt4Lm8wtYq+wEoWEdeUwrc0
rVoz6J1W9e4Yve59tjwuravjtCnJx33QXFh2R6vo5MkkQCfDsBsEDfLPy4p3IYtZCL5gMvFLzZhF
cOUc/XQqm6ez+8jVzuu28lW7IHYiuPl6NKG7hQ5SySSu5iayBbTi/muUn9IH9e0LnP5elbAT67dq
2qmHMVtvWxrdzicQXz6T0qgB6p9Dd1u1BcbWzjpnI0NuB/KzmyciZIcz9d5Ekkp4TDXFa0GzUiML
1UW2mMftLeeB9vBOub3TqsixU9FHQA4tMeB4eWMnXswRSKk65HRbUJfwCUbLPgQHITesdRIA7v8q
c+p39Bvqx0mMqH6Whefx3KOJtBB1zi2dKE9GEJ3Vna5nvNRJRE3UZYDyxk7HvJEu73YpWMI4p6wy
PMbw1bR00bz6vXDWPENifol8MD327dKOZ6txi/weG7SOWTtSbM/1DGgUCQYLhwrzRvrV3OzmWjTv
Nwv3YqF0IHSG9T9uE4/EjVtz1mEWF0BYz2LXPklMHCPhhCYhA/Iow/1NG0mGG5ZEDhV2Ktuk+DaG
J5UCFmvSoBUGTthaZiBLnQLXz69X5Z5QpunLsBoleoCmEqM3oHXqRZKrWquMO3P4j8VSP4W1SYMR
cJpepUzdmNfP6jVq100hI7r6S3zS8v3Yv0o/l3fi0mlaHefFtu/EEPznY6EhdcsdwRBrnwEQEiOC
mM0WmeT4mXlW6Z2nHgKpvpc2hG4nIsecCIc/+cXVhLif1sjHZOPLdjOfhkI1uzaKHPEkXXTuvg8C
BSPOi4akwZQttGz3Tjwmih+NaaL3TqWMY2f2/W2wQEiWBEO19JG7KZeMJ319JtRR6LfE5x2M3dRY
tRM3Mi9buqYmggo7fk4sEYNfK6FgNDOIR0Q5gTmKctUr6Q4Br18Uu9s30LAxDo+VuAO1eLHTefj7
x3dejQjZDa0cYlWCjPH8cbAJ/0n+6zigNoka9ZvrCo8LSOcjAY//Jr7dTh54M95/TCH0xYQvY+v/
OUTqU5T2uyrdyWHcpBJhhM+tIB19dMQjFXK87TKj+wAZUhM28uGu2gIDs/UhVARxhAjU6q3pY8Od
n3Pd4LySMCGsCI9u6Ym/Rg/JERrc8nHB9U5ojex6E+9pWr+0CpeOUT0u/vbtD7RsX/MpRSuZgEeq
KrGQ1QshWgVnlSDNx82cXggoZ8BrWTTtBXbrvvddo5NcJZfag35BGG0gOKy/YtvALnZCQq7oCuhT
Q7Q6ibil96DAk2z32bQ7uuVLfVnP3W8O8VdPlSZ7/4NrHVRW4HLMfGokJtzsM34Golgp/VHio99p
kb309U3tX2+DUOXQ2n3/KHJ802H29HL21gQ4/ZqhD6EAc7nT9v8NLVpDnwcba/8LbYrOD8AT1QcF
UE9UIBjqNXbmOTsIpFBUgsAo/v5p7PopjPf6Ja94U0h1vJL93leECAv7AHTZKxIUsd5MCt9DthbI
2tYcGAnE4C+7ZxNoWiSprZ9mRyQNOP9Hz3NZlWCgXamBauj1XWml2Rv45jCF973h5zT/cagk7+Fg
6KNFIpLps+JEtEwSz2SR1SDyY+91u3KL5/cIbht60p7Bb4MchDUWOdl/Av7W5s67t6+PnPLb9lgF
CNHntkaIW3ZrEl0850+eFYHbPhFb/UMW2fE5OKOqgp3hxi6Cjb9yP5cJESPcA3BVn/JkYjDPW+1z
VxegB4ShgvmCPBWEsGjA4dF3oTU9MHE/Tk+0zpBr0yV7cCdKFg6agGIdXUCJ7pTwlnKH7sf+wJkv
B3BuFArNo5gVRb9e8ZnNnGRvVWXqNADAIqPYAJSKAmEg83sTDuV8RQcRXHt5T3IpzjQQ9h7MjDth
QfIKeXQ5IpyvP3NqwEaYmtJRNRP9h7xEA9DDczOiyXei9sxCH7ZYYkTXuHR68vhZJvk+FNY0WCk7
+kww1KInajexIsVG/j1CE/j2JR5aAczuiznZidfM2SNgEIM4HX8UHKLcw+BzfE8sCk5TiARNeIyw
ejnaf5wag0TSc/hge4lDOYdf7+bSmY7WilZnsJFNpqajaZ5Y5MnjzoYk2FMcMpCkdog+mVBuJSSR
Bwe6JiuyrPJBCVxRMM1+Foxso980yYMUD7Bi3FDpte0YA8kPe9pdxctSabTpJyQvSjdvhSpYrmhQ
ANYdA+CdJQjBANQtQn0Kqt/wlmfnP4A3sqVDGMJmv5K4S1oFix0F0V9QAlOE+eU6ew6NwW+HMIwq
DyEh3GM9ysLHC5mhoHCZtV+7izF4Gm/tLainW1p9kOI+Es11jU67IbghmUj9XOe3AjnB5gdxsskQ
asvdx/P6Sb0MI4pFZCuveUx6luwqDcCIimtioLvZSejD4+Hmxc/Zls0FXLZdzgG49Ev4DL+gWKDX
ak80Im8jhUl+3cNhAbBX/35Bxl5ygW4xPYIhkgS+FJ2XKTJl7S9IfmHQyaVgfq+7Netv8kc/ICfO
2ar2Wxk5znA3nl+S0tSDDvtCG95OBBrJrbKID7Bgo+QWDirqYyDE3TmSdhRa2MZW+GwnehNIJb5o
HH1METc+Jx7mUp+FW5iViCnB5ZoYKSlJbsXj5rVOge9Tg8LI8RlESxTZIi6JMKUgju8KTI6GH0cd
R+YMrp5SpaqssnpzlE3dZOjmw4vt0kIL77CLgLX5llHz8SlGe3XoM2pjXjLITRID/dnkiBVPn5M8
KMjT4pHCrIYvIiiqogxrojgPsyF04Feu3ZWsBNdwQ/zDkMKF5Lq2dLRn6RTx+qOvCG9wMPeK5nsR
XC32TCZ+VzRY7STbmWcxSphdqfyhNUBqzoJ0erMQW013L35QrhIMe2+Fdpl4srwaIEFFV8Q+Ulns
Vu3J0tf2g8TERA3Vhv8oe7Gccxu+XGvbOWy7IHUOXFErAvjDUpT+sViM0K3Dk3RayZamtivdjRxS
ZCeg/e37lr7Yf7PEIS1efFIEBhXKEdnihwv8krrSnVnsp6flTJLNc/SSQkyq+2WoBkJy8UFN54PW
+aYz5Iloy0/afH7tubplxsj18JN5AR6cGGiYgFqv9qyMimHki8eRoznHtLXTjn7KCR9Sw/ac4Nkp
PqEVDbs0tlxHuLhoHYXz5AsK/Ptk+pFWgMHHIKsvyeYEXdZDhVKKACPRcuKReyCl5xrTfnYewvvv
1qTieDE1M3Q5lqgVI7EDirP+Mc9UFeMQJtRPBCgLRGLOTlmaicpQwnfE6QMK1F1Xj1EFLwv8rY15
OHE+cB8qFXpPvPlhOHXehZy9cE+LTIjKPE/THTuB9h1WIvuwvOr1LyWrPBNo9hv09e0CYG0b5vI/
DsD/6HtT9JKFBeGDjcss6jHhguo1GfzibSxY8Q0oM2LjYDudWcAxIDt3C4ZV0rl8QIzL07y9g80V
AKpa8pjTwXMSv3AsGO5H6p3PHo0SB0a19cKdBLKtc4KP8a9uAhEepjimJi/SFAkDAAlr/LMWVqJx
msDvvRgR4uQvFAcCFcneKwRoOQe0AWWp99j4IuhnY/+7zz7YIzr/xgnOtdlEvW0aXpQYkmFqp7WJ
uvbDrMuYKT33cXpxBUDGIzt3sX3lBweSKJBeKi38DVjStaHft+hLQj59VOhuPbDjUNWtqBhRPz+h
EtQHjitDO4YPZLkntfhL5s+4RUrxrFtA9C2sNxOZRwgow4YzKAlC8GRHpW7B2hYQYO5Kt0ECVsD1
k3G/LOJhcQbivlwWwRAcmBF1DhOVpv+BhMmfIYUFIPMFLR9Rvx4tUMZM3Hw8jTnXOl73vDMQwric
V3kU6gnOpuXC4ec33LLnhcw/YIK2aJ0oxBYDVoeW9er5obCcZYWwYLNDjCajAgL8r88U4CFo0kE1
uWkZahL1w8q8H+Llye/geeuk68DSfxGeXMA2leLghqZ3udKb9xledDLcyL00IpeW9Nui3/dt4Jus
lN+SBnGxYYXbzWiZzlbac+2k27B69Mf61p/xXXhI3vbn48135EvoUrEKRgTgMyxhVOLcg8HXguc4
rWPnmKAa7XSjpI8XhMN7+zFpKcWdN90rbeI69/FplStBJE85Hg+jCTPSsIKk2TLu1YBD7wdv/8PB
0YuHM+HaEMbbOj2oxsky5y3YWb1GrlHc6hw+WacSruJQC7VZGSljvbPheWAN3FL79na7au7IV/c3
oDe86I2BJtlY27PbAD70x7rJ0UqIgY3mit+Vez0B+OTt/bPRo48bWayJFbWE1P0SsBuXms0N4guu
gPgMP3HD3ge5z3XJtCibnCUCfaAnf4xbQMq7qyjVemPWNI13YBfARcjDNXw28AH4MDU+EmubQ9Sq
s6Kq6eUR/e/UvaqL1auKuzs1vnqLT3ggOV3NlGeEG+VAxlp/06gdTlWFuPaY27bbtkXOTzOldQoh
yR0TGlgV3Eg+arC1A6vj0xlVRwkXwagvPQ7IVDdSbrTrpBKKsWcG+tzQu8i6i/D/vlo0bNlLbL/+
jH46oApmRqotGzlBR38opa8XDJ1EfoBF+nOV9oSUeiBJU7RRnNwfzXuIPhvKQVdS13LRmfZSnZwf
m/U6sZYLAneP2+2yStBqNJEu8HtGI0AsGSoMwM3tIgVBgDFZSMEeXQKg1X/bDksT+AIwsyjBuyKU
Qo8VciYbrXzJyflD0BSLJJl95U5Pc3m66rdAGmWDfblgxw1W9Ge1w4B5PT3du0B2icUdSmhLWqug
1/gD56Tdtl639A9lfJx3UYBZynLv5XW9RSLoww4USoCu0if9I2aqIDWrTOcCSJAiW/XXtkAMNPAY
PERjcsSmRZju1PRIB8R7y0fnt2gx4DmmP3sUiBaXS0oBl784+Zgwd0eIEvOxoAY1Jo+jgmJvPxAf
R6PnKS2yof0UDeU//mjCwGhQ8inYuzwlk30tm9ltSvJCXTXakDQHgr6xt7TI3Mjrc/zmtn8Cc/XZ
/lhhx3IM1GLNHDWFhD5V3zpkah+P92TbBQeDlXZXmWXkoY2F7+wQJPuxAyGLvEitezaHdQCocbnD
QgKfPiDnR5n8DzasmUMvxpRXR4YlB0cEP3WuoI29iF3uKtFrRbpwOh+aT2H+EDTdBncjKmar6ZTm
RVuPMXt6aGAHFxOv3nwPgEeqeXsJup003cdGFq0WNcJtSeYwe7fj/1921nR3mZge3JdRhPHw3DmZ
A+g2Z4Qss/LP61i8LkU53ngJ++DCz2eqpgwwtmUTHtcUiGS0Bu+kC7tXDzxCq4oB3HmNqibFqTew
YuCsSYa9Hgvh2ABfHs1N/V0yT+zr9lEG0r+qXfdgo6tbYZSSyDfidZUj5yZZySWI9vmoLzazLaYg
ZGGxwbFS/gRswxIjTAAGaxskMjA4gEkpTDaBFl8OKZrYwJ3ZNueHLOzHg/SV0FbSQuyyVWGXv77a
fwneLW4gdWYTqPqarN3wRLo2515WSk5WVv1NxpKaM+YBkhRD2aqf6e0fQZg9McrTFrPqsPWjDwU1
r/wFtM4RiOQPW7BGWM0oWXZAUEBcRyaaz6hT2JkO0fghwpwjTgRL4O1IYB0/Rx5qXFxuQJ9FIATk
6EPOaLiwfFXToZl7ua1uA0ZIQN9dpo9lX5ju2+pUqB/UcYng2jA5VMuot7L0/FLpA8nzmuk6KPsB
HvF0y/7/rK0dR3xwlDTRODHuoYzIJeFxDN95fG3MVpW+X6di3ffUq0Bdshni9697ILaz2XKsfMsr
JqLq0vbwZx5Wr+k/EHgYRwqehCrK2rrc1uWTuuJIOt7wGtGxdLzZ57gzcqxuyoTRTVwl1f0xcy6U
ong2QU4n+UGu37g/7JmPMHmP7/Vsp+6EYuN2qOnhbbgkDGwzqe/1LueXHb0SVeyNd0LZ0pPnPitR
2O9uA8VybNhpC7lvEdvaScauE2/3NWOdmyi2D5AENA27k4jlhKPF+9+8lWICXqKI+RUVqYMT3LlY
dMi1FhGDTCw9zQAh6jB9JO/GME22vGKDPUzGpJbOizH1uBBghv6/+i2iBL1aNGsKgG7bxd0DrvdZ
Fn5Ym9/pNr4s1yyw0zZevEPjbNXNpT9lxG/tbF0yIS78X5QG41A/cSHo98um6nJ0TUkLJ1a6m5VJ
vEXhnMNC2lAOgEB24SPHyYnRLz7QhlMVc1SvN1vxVqW/c8qrV1iH80zUVFyB3LeLo0iwLNnfU6xQ
6zCDwEdN3LQwcEId9NESg3WUPjBG3590CiATP9avvWqkcahZVrFnseDubWCUZFfGys7Myyf1yMYA
7T98VfEPzhwmcRa3r5RfYU5RMG6LeACDdZJQ4OH5WlC4FhzaH6Z1z1t9msoyYxPwJlRhDxQdbxyP
zSz+LjURDgG2DecqgIuos9Q+zEjRgw8dc5Mkts1fQsIYDJjnDiODcGUd4ulDHZEb6CZE10RNKp6K
2wsmEflhUIWyQJnBc2n2dRY+uLLGOt5JXDqmMmlHZNN9uED3aRwsUVDp8GFDOdAgXpgCQ7bUKgWE
BOACKTvAQoOWgkOiZGclDOzrdR+SDzTvG/EvdzYeHiQ/A8uMpS6ExpL142UdLM1SjSxPFbylKmDE
vRwO1o5QWcoYkYlKjdQmPJPXtLjkns0nNcqzgrzaXg4GyDpxjsT1hBvw74HBuMo1qPvgWLuiKSxg
YRYeOP7fxupGwR/rhnqYfOEcVfspk1pgo04+Jy94Lxjs7mtUOQagofo2FJotQyBrjQjcC6/anL0g
K85A6nJIHHiD1rOliJZ+tGIv6Wdmuoa+zVH4CiQ1BlOWh0FXKMuqFIOx8A0NgVwGJgDWY7SHRFG+
XT9g0Kq1Bs8IkL+fIYAVUnnbGn5eouwE/7rXn/vJx1xjjBqqHZRO2jGAGoQjowD5xt9a6FhimYQn
1XHDaClH6jkc3ztEztzvkc7ZaGEeCzOOrIqfmiVUEio9CgjJmLnYJPb8WQvA+xuDwzJGoSn2Fj8O
5U5TBRcvJKTFtWGdod0hLilt4TOlL5F5Iy5fO3SVDV10oOUCEeo+N8WL/7QbbjyDPKyFe/cfTLsu
Nv982vcGCHNUmXda+cScKTB5+N8I45zjryz/UoVA7YFL3nMDrh6aE/Ubi6uBxMpI50wAiTln/2Og
GXCXu/plL+MCoWN8u2Gb+2CAJBeE1SjlF+QB3a4ZmEUvdgfE9/2w62mXHi/pSJ4wm+QCKvmdq2Jg
hAeWC9042aXqUO3ycsYabknKBNV91LAnJbtHkf7S2tPSag89xK81PgYLe7IJsXBnZKHWEJXXtimq
o6rG5ZwspE+MMt4XxLBqTIJmHtm+smACam9S38J/4W04N9biHQw9baA++eZiuqq1H+nqqGYMjAk0
d2zRWehnB9IHPvfdQwSxA/KPumEsaGB6ANy+Dn3/EqFla/OHs4NtZHQ/ArXRIsUJIvhn/RqxuRD/
pt+LYn4zE5xe4STtI89y5Y/lBtLvn52dqr/5JRsKbySHva8kHumsR20uK1+ndTm8TPu9+mY+W2hu
dphfQovqmN0Rt/d7xLsuTt8vyuiCyz4xaMjetuwDjjlpMllwy/8OFS6x+ttNaPwPzsYfEVSNzf1N
krq02b+dv+uPcmIKCbkUZDhGfZi/8fn6R8gjDyb8ddJGGQMowv/vukn0OsKGphNpZhC+kidVAaVv
3iSBYuMdfl0SaYEELU7S72pXGVUYGpsdA7b8ZMM3/2QRQiSizmUF/KzLc8jd1YkiV7G/QBT5wnOF
11TC86j+6NQ3BolQAA3OROMNkN1S6wyDfk7E+Ap/Fu9SUQGHLq6+631Ltl9RisnNOIQDETdOfiWm
S2g4smFA2p1fGPrrWH+RZpYdRhfdw4FEs7V2IivSG58gPX/lft/vM+m4P1SbVJyWh67xRQcv0140
grMqe6Vkz22jqfe4KlQrhJkkcwHt7XHA5KrgzGYGzmJDMdOaPGgGV1ZbLMbP6CIH5AHircPietSN
k9es2BTrSJfw0iaIi0nFiRyI4U/QQBjY+vRuFpJk/tBRH5F5KLpMLxowjvW/151sOxdsS1widDsH
B2o+kbDViSQNXl15XbslkmULPANkuqQ2s3nLA3PIxl307Vry/0Yt+m0Njs/HV9RqrW3H1S8BDcU1
0RM88DeDjxxkk2rEz/zKNf1GQ7nJ4R5OjXwqt0ktDJZzupkuqTT+sFcwAgtVGrGF5CDWqeiIssWg
wxzRx/NMLifQ8N0d3LE+kYO3pwi2Zjc6RTJFofA1sf1ndjDzKPAT1J4mcL4Tgipp1Du1gYFB/y0B
rCuR3IkGhZ6CF4XgDXAam5YHKO2GO3QdXPVVZoGhQC/3eAqk2f2dLW/sLEql9itE0lj5VfGEugif
HQjxsQ4EiIv2V6MzJEBr/h7kw2ANO6kIBEEX1YMBCmhtp1xiMCbixoD1ijN4IKICKXWROAVNWUG6
iunItHOT7kNNLfrh0/BJETMeimTFhrLVpaugfMgU6LfX1PKbIYk4knRLn/hsbazStzeSC8jR0S+N
2WxjVjjZCJ6xlg6NgGmyDSWARWu+hf3v/7g8DeVZkiVWw3cM5X1Hen5YVEzIl2EEi1GoZuXCTZiG
BPA9VJ18Os1r1Ya7Y2gVmAxh2X5313mrrAPQMZLcTyDEj9ZEx5T5X/Pq3CeK8ic3omHJgEIcgFCC
GtGlEaHky1y2nLtz8ZK6tZm7KX8bT6ms31EKHzYvhZ7eiI30ajeWfuosNxWjcyGPS6TbLOvtl8J/
4WMsYU8ipUMhmGXIOsSmmpicw34YUZ8+K7VpUr3y85EGf3ITyFVyAOSUmZwnWhwvSRn8aKAFEYOr
wBIHDKVbZ/rLcSyQ7CkQh78NvduF+kirIrgiEvAdrwt6Ma+FebNoauHT4gdEyki974I53c3Zw1v+
Jz0BfGL+oJYAxYYplRM2OwreTNk8JY5fNxHOZ16CdyO7PeZfeS0ZfBcbT4hi4jTyawVn+DhAP8fG
j0IrWZ6+dIy5u5BEQzt1SQHEZXOAUhxy3tKNNODBKNdqpLkae9Rgg93W9sqW27tQhNiz+Tp+UyjT
PO8PARJ8S+I+xgKq9Fbs/wAbm4VnBu6fquWBDeD3HANkg/g+h8Xjx5RJtfE8wnijBn4chOAp9t6D
nZKSxEE8pX4Ew1dnUX/Fc6JjeC/2Rv8qv4UwEe2QjgD7K5SUYznYQ9eOZGl3yEejTro2wwSdv5l2
GelLRfl7LXoZGIxv2gS610bkFrMeWNYwnYWQTow2dGdeoS5B0l/8VIIpRa73IXYRTrUblNnU6/ye
/FXU6oBF4ek/lmjZuZhqxgmdoeMq/UqkDEOOAnJbyodRnqc69/BpZBmBP9SkHsaHQV2ddA9gVcLv
DjX99R+9jWNWWBb6p8fU4V16PAi6lRBbBvcFUHOx1nguJV4cA8A8dxBL9cSzvj3TykqFIQbEmjUQ
t2vhk3YFzcYdl5LPqaZXbg/7iGP4qJpZS0gGlqIC5K7DB1qGDXbzr4YW1b++/u3210vtZ+FzPsH7
mLLoHAH982YoSZ6nKJvN6LGRETqdYUSNZ73azWJp4YaLFkdJjHQulJRPLaZaqlut2kq6wEXqLyo1
6OY701vSy1TKgoltI0Id8oDOtVXlE+ixf5Uxvi2r5PHmIBx6LIz34wt2dBhedW+6655OqyXwZ4QS
k/tZR+GqL0OOEOJsVdtxGgOXzD5crG5oa0K+xX72QmBxKIs9DtKM+xbkbQo7tIkZHuLEBoX4x8g6
qv0qPQQxbR6fd55T4iqmBZkynVEsS5ws4XFDtoNNCZOjE1Rv3+dBetwt5XaA0NTPy6GZcw4QHKP6
JID7oB/hpEsdd3SgTxCe/Eio3uIf83rp2JFh0hHW1RooUuOaoAS12JMfZCMzF789NFXoD7MG2M6J
9SQTEF/Q5WkdV1Bz1G9IKVsc8VJxnSUMG4xMSowCOq6yAc2Qo89wULY3aXTzmtoRJDk5aOwi/zQx
EbrcNhbKiWKNgOk041tXuj3lQKgA1jWTe7i6L81bcPbVZMz7N4QVPZOHqT7lOslTHd6P9DtYjmRS
3UwqlvRcLFE2p3zK5DIPgvQ7H160x8l05fdoWtWlx9FIcW3f9EHzu5sERBJ6q0zCfQTQUxZOhY4B
t7vgDHc62snZejfKdqxSwYKfjUjQ5PfB1YnTvLQOb08IfN9qTRqbUmqK6kgq7gxL+2A7RbMUSDxQ
CwPK2oyP19q0AIUywved09QMFltfg5eRR2p+DanJfhsYNJoJu75t8cNP3xmiMY/6bwQZIM0UzREp
QlJ5nLO0e80YUl9ZqeRyhKoEtQ9MfKsJotF7KIgydgJkfB9u3202cFwbeQFtkWwsAF1CYjr9aL8G
VZLGRBJpElGiAgHoHJViO1Ex6WNdBkui24txeRATZDgAlg4Z5EORAlD5sjeJY6VIwKGSklAmwCCA
qf+qaMO+R3Ng035tAVbdt0nMJ3eN5spPa6YftPaewW4mpNN9My2rbz7eI90bvijVkDoGdYbBoL9Q
o/jxGDCIwVuVeHUyYU7hBL5t7D1gGFEpc89WP61R8gUObwjlrI8458q8T3IRxJxp1gHsYpgvo+Iq
asa8KR50FpzMIjRXNzxulEPViUcdHRRqpNyybvvpKyW6c2vMTfyB04spaGgF3KupHHBlWUDHUCMl
fc7nvjht6DObcORRGNh7/rDB9aJDmTFEt/06ghlbveS2PK2Njy/tBqaWt3m9Ur3y/WBtUjTvnq2W
uOKrUzqVehCQNTHxOHTsiPjNWaop0tlM0bev18VzZMBrd83ak2XiJYwBabJw7zzn2jwvtRFvsuTx
t5XXJHcqgKlJaxC4+trDR0Id84RLcmfLBp8WCGXlacPRQOpLkrWeiqJvNrfs9vTRosjfpe6JEeG7
i6js6yYAq+ovjMY7IohJZYU0DoWwRiilCtlRRjvS3xxga5KoIEsRaEJqpWzin7va9hN8XKydjP7m
zaapq/f4zTXn2tWr2soK4e8xRalUI3as8BKdqGxUV8Qs2xTNGDi4HUuV5nv95wycRLStN1htzPUq
tEmCUaPTEErE4bFiEXKnD8IG0VmE086NIOmJ4Ty7O8P1S0uyEvJ13NRuFsm7ackRlru5DhAOa5Yr
yomnfkf191txZDjUD/PosU0l0q/5U0Fy6/DNfvwtzuHB7+PbpQt6lKxTKLHo+Fi2vOaghMN5wpcO
aPduflr8A443OoNNJJfNfjKGOqayVP+h4j4Z0UuxSRhF3/qskpNT5vvV5W2/u3SZaKz4IMT1xFev
5Rj3XZbjXZVBiLhJKjQrVCrG326zNhTvUnsPwlFx3T/674M02JDs4/jWPEo/3I2lxgZiad5YPG8R
HZbMPzpu7ydCF2oEfvdGa4HuIjsvx5Q3aGAPJyPqBsCM8SXqGrBbVTGf9lsmfjWBlppTD83SHZcY
6DXtU6/U0KXHnfB/hOyWZZSu5ZmtFiPQIjhhvPKJUbA/quE6ETsN9N7rHq0gzmGy/aZcO3KE/qn0
pZ1cDo65fxvPg8hxuETXRxd+TzFVxJkt+Ar7CxS+0yrCGQXQ0cR2bqPFRrnCqrG00lpDDkHtetfA
2JiDLh5pWJ9jUcNLaZDWv3uN31UXnamGRXrkRZ16I80d7b+V+tge8fXQSkSMdkSGyAG0irFrK901
Yua/hPVHip29tey+o0klGntDh66QxQ3Bp27Ovor00nyjtPp6MwCUDJtUKTWxRN4LkwRPyUk54pu4
CvstU8OfR8raB63F/RMc8cPDdaXootueKg+BjceXACuxP3k3R+xecUCMpvKkJXsdYKV+rq8FHwps
KUePNizd5sK+QuD7HBDM4yW0ooaViOFyFMQ6L5m3/l6WV1mZtny0ADxOnvDSctkp6Fli+quh7Wwg
MCkx/ZwEI/zIMFO/VRUb90kvLlQgvTYoKAFbedNFyH6wWQVVf9FBPanixMaGztMNGmSEK3DlISfl
9y6M7gTpVp//hZ/NzkquZ8OyDlUpzHyO82QAmo3wpXek0GZmkbR9qjrLFNhpILlF3vwDiBrkjW3b
FzBqwNuATu1jZMtEFFreY7gPPEnjPkVxv8iJrR6j6FIbLAWE39AtudPxY0c0oaWVd/9wRVbo9cVh
XKajoVA11Wo1hUtR28HzC+ZWHnySaWG9zFGIu8vWnhOF1SvYEH7wBBDME6MKumVpSIlIWGiiUY9I
vZGCVawuWSQUKKzmuU2iEMGSqpQPdhn/x3buoIJ7YcmK0794Adq8ZJHUAhWRhB6gsGsHwRPmxR9I
JT4RQtKUmxQsEgHEC/5+gOOKng0+atUVmRMTrdNGzyW64UKOUKfLhlU6qolnsqSfw2TC9n0W5qlS
o8FvgJbqwgfFdrR4Wg6dhYUQ5EQtSrd50xARFz813QKb+8N4w0qEaoC+dgagt3keICcJ70doOO/S
m7osMPJ7EPfJXcu2bExvRSj0vuDJLuGxWKTIBKVgCpuq5VQAGhbQO0ePm89PAIjwmTLDwZOPJKGq
0RpQLu41Xu6a7gBj8T9H7F8qHC4KM023qZ5cuDKilOGYC1/VRh5DadTRvuPQ0heNSl992SwN1hAh
d/RQJtVOhGTQfeWNoJu7X8L1cwSRgM+QbiroEB+hyPwN+JDqAqkF/CZYBeyOOCE65F27HwUYOCFE
zEB8+iQ8Yrchy7MhuiPvkCouuyz2Mqs+r7ddvqsa5WpVgeMarEsWt1GDmWEspfVPbaOljhfQIyMM
VrWVd6PNSPhzZt0/C16ihlZRXkEyI/Ahhy6rEQhcG1QKW3ocvTInG4ArJ6HO4+7Tgbd1lFgySdRz
ULdmCVYCoPoUWWtTXHW0cuU4rwPh+aWCHB4m2Wsac1WT+Gr2uxwDmLoaW5q7mQ6NiM3mwc4z0UZM
rrOFnhxWZof3r+KPLqL8Q2/ibZ/mj3Y46HptVE2Wybb6nti/sCsRFyrbBFZ//CdHZYwyoxR4+WKr
46wLIXfU/IBHgbju08Jf7yQlrFzhp4Nsk3f8l1v8MZwe1NKLU8FDOLwgOpwMbjc3xMaKKZAwHh3M
ZMtOvkPWrOXbsO25j8lUZn3zkeCydVNyjQr8dX9paZa/uXmJhhEMwYV75dG5j6pffYPgTCbQcY4K
FReHVm30VAgRwwWv1xrXZqAkQ1MQgFBAzv3UphNzCg0kUH5XsTt9ULnt0cKuOrTwdGjxT4mjQzar
QVld2B2S1IHHZnV45h5AG92BY+Cy9N7BpfniG3L7Zt7WsspjC+MJqn3WdLRko1xGfqg/dSrhllAO
ZBEWd3/d/Inc7i2JnK8Gkfc8I0KNn0QEqgDNtPlpyJpFYGx7y6smytT0tkwsglWhUlM3hpKpb8sH
qA45am0aWPL1G8r7DZjdAimDV0wweq2BekKmNcwdqGwkkPgt30P3uWLnqlJtJXuJNXa0b+RrNWHO
xBLO1yofVtuu9ykixm1gQeLbMmTvKdSVpLAgZWwT8SZPE7mLZZRppONtLZZCBqusE9NkzC2x99HN
MNpSFkWXeMfYZv4eDem7ZFanktg4gVZe4MCCiDpWcjv3hPUMyoumNYJMgIz2NFOXMUSZI/KJwYXH
zqFj5mTorcSpGW555pYHxDMmgVaiv9FszjtMWgx/aSSYHO42HUX0QYhQ3GYYPz615i/09Im/i6r8
25Wr/4zT2AFqd9D51JodOEV5MymBXBWL/lzGCAAsSkDovXfRfrVTEawoGyb61NaKQwzt/xGa9CYB
+PZnRadofM02ZP0HDK/ej4tseWpgyDpQb5ogRA4kwvbjy8DJGyP5AeV6K+IZW9j1HKVxPoq9Pg+J
zWJqNH+2IKWX4WEcRbUqfaPJU/BxCdYu438DZGGd/n1imzQazenbk65MFzgSnw/v7L3CSIGRrpjS
Br3qwWXkB4MKt3cSp+9hhQ52DbwueDvBk7gP636D/8BIIbmWlYvxIgqphgRdMWOOsKmnU3aIrf0C
ZMM9/cBdJV0WSzoYeptNfsSom3SLFsgANJO4MoYw8pMZ8CGYhYZvIYPG9fww6SaYy9NgLmfhGu9W
YFZsy8toIXP8mbR8HiKRnUUORQN7XTusUTH292hfjhX19YkCQ2UZFEfYflqE9SqyVvuMmR+tvAmp
NWR9kM0yqd1NDmwgpJVD3TtkhpOAirFmQudF03G/5aeCRmozh+n6NXfWcpuP51UDxwt7kg/Q0YXX
rUWfsJCQbfY8ADdDOLv16aUwsl9yrdEMSQ1oBKEW7pxKdk+7xtuk9kJRwD8weMGDIrTtU3eZTOki
fWXPI6173vluVD7oVady8+lWoc3Fs7CembsH8zSOtvRDyWKz5M06/H/Js9IbWM37lnLthlnwuA55
+WjagUPlUy8tewC9sCuBtR9m9m3rSCx6KIfnjBOt7PO/VPg6FEH7booMAClPdHlZ9vozUIOeRj47
qtOWrtSbCPjsPi5OQwnHbA6iVR2wh7PlF0qEGL3F8azC/Snf5GdJgFm3hUQigaXUkzsIy96SH9dw
Yc61fJwpfnWlMCddDnm2P1pcAiL/wd3xYuZ/wEW/F0eDZu7SCPQDrRz9GZ0EZ9369rm9A1AroZzU
P8XMgGMpycs1cPvSChjvM1nScO5gnQgLtR0Ac/3o/2pa1BeR79JdhcpJJ4sMn0plmbdhMj0G9oBV
bS6uFXNkkRDJqJvKObqVMxM+UZSFzAMG9V+cSlovYfT05FsAqiomh3v75dprw293InWqO3+jCIi/
EXVnpink1XhxqdXdKOJky5U+TJsBEV1gHqtviaEosdLkgq/0nYMqYXP2ofj05MwOL2NA+fMagxp2
tz2LPO0bRG/fZ0CE/YvSv4C9EJMjQH6dkX6ccdzL7jfcsz3XisPTDHq1Jh5r0MzcyvPHSbPBZpuJ
u9zgpbaSOuehZpF2GApd1aFet4eE2afzbRLLgavBGjyZkGaGAuQLV80CUltX6qlM8KwjPwTs076L
lY4oGKxjxVDeOhBRmcQ5TAXsz/bJ+P0xUiC9cxnAfQmfSWHMWQkWTBXLmRZ0w5pDczA3Ddri3Hy1
Rp7pfgbiQosqqmXdwIqXF4oLlBfweJcUBE6NTc5CT1gwVpnq24y1xDFdLvoMjWvHax+LGPZovHUd
ROFWaNm4bspFQOZcKv4bmfOHG3jlz+JgRTVvRWJn6w3YUmRPDcwkEnR3uVbPBPbswVMHoAMM7yWF
p42D22LlTI9tIEJhhB0b0qmpNvJO1ko+tBF3P31z6QGCadkFRaomiX9TtH/nAe+J+uRfCzpTKGKn
8lzizJMYFHb6EqFQzEMc7JjFN9i2+otooxijryScxQLV0jk103bH7vvtxcgJrKZBfhuCGJpTi14C
VDtmIBAdejLn4RM6MLS/zGIp7ZwdS46wrAgDEPjHifeqT1fj5Vq+Yd9YIbnV/HKsyle69Vj8IfP4
O8vFqeuQgaR4Zt79vS7at2T8qa8spryl/IZ++m2Nfd6OP+Ly0QK3R2FPIN/aLX8tVEax6tnJUAgF
m10wcVb5zlosEiw/3KCB6W+751mZjgY+gEPMPwOrU/DSDhuYEDyk/P+8mMKU65e4GJUhykrH2C90
RU09bqZWCRbnUZuSouhRTMbN8AGH6bv6lkmuYrnWUBae1gglRgwFrfH461mQS9zh7I0jB49AwbCo
4elA2ucAnct0RPvhUCwz1EFEPWT3h3Wm0bM1siDtZIjRAroNgsXyrfCbvwSooPnV+CV6j/u+p3FQ
SWe3N/vpVElZf6P3v2FLyRazlxOOoBUpLeg7PEWYYbwOHkeZfdxnwKcv7fR85cNCd6qgrXHiDUmK
TZk2AluurD2UbZJFZA36G7V7S1mfvudKVHrTOTu4Kjom1z8OtGhb/Cemc9LyySvCX4ns723B5cG7
PXO/w8FDjuwu5K29ijNd5ln4T+tD8HLlXb6LRdQisr/UAlwgBhWJ8e0ArNXSWDQ/2y+WrVb4U2W9
qq7kMspyBO02Pul143IOv3JfrCHtCF5K0KRsFxtiKG2JsFnaZs1HjRHtxmSX301QF+FLwaWOssY/
MNNzC3tN/dTjXnsLiaYrAeqAAI/7WUFUDhs2XQQuifke/VAGgJRYTRS96t8Ew9G0kwJm3Ke/CBuZ
O28B0ecGAZ+WbUJTL7yKVRl2tPRteGZ6htiXAEEI+2jPVxqJJOCt0pXN0c/SKN6au1cq7wXbB3y/
CxH4S7WKdjaf9BOmqGPUJ/6yzgJX9cI7R8m8Jm/VjMyXZTMkBjFx4j1C+bsysjvK8sZkAihZMHNc
7sisuTiNfUHrIg8qqCiRq4zt8M+ak01NWcPjVrlihY3ZGkPDUYGnqbPgdM4ZranJRwsq0v4CW+zD
5ySJSbPFOgbAYJtMLDULpk1BhfoG3/u5lZY8w0JBIUUaQ01EwwZTgdLo2BMcSsYelUXr8IkaqEj0
/PeJV+Cdb2yZA9NNJ/amWLqKP3W0pK80l3mVbR6wW1jv812ku9UNqAmQkhcfqanSJUzFvovxi5Um
si5P0m2m9f/+cQ1oDnhnWdGOauerPus3k4zx68bsTEDsvl+TY0Be6wYT1SlmkGDXMaSEDsSkTz0y
ypClk8uluxcBPyptWzJ8LNHQW8XpOYft+olDOvlmRjJcrFUt5PFdeLXyVuwKyvW7V/KPUbBZ5tYH
9X5kApY3QgaODKdP3kijC0tumsGNBwJ/kHm3n2K31WIYJmnX2CK+VOb7E3zxL3SVPFqI7LKDV4Na
A1G3tNWUbF2HmEYKeYs9jp+Yhn8KK/ZHrRD8ikSUP8oBExknGBEn5eEiwwa74h5eM4GHKcFstkMS
2sl2xlDXCq25YBMclovdTw334v782BOuwwOB2ywMaP6Ls6Tqt0KAhJe5dkRdRlpGnp/GGEjb2ehW
Qx8KcwHO/Zr8qxBaR5BSG4LzVcmeHWeF93G9xJ/m1Y7AllaoAvPOEny5knqns1I9GtyXDBHDnHch
a4CcFPezGm4DuP5iJL/UpVNhPyJkCL+CuEZg8MUwDZ3twrak0oNTmgD8CcytSNy7wZQbuwx1KZJJ
E4H0Z5PVifPYvHv/s64IDe7I8qY8oyKgbTOzWLl0u0MJ31ZkIy9ocp0TO3IsOMPZ7/eerH1gRagk
8jkFE2PUMaoS9qsRmXVQY2N/EMfb+6NepZ9gOc/p7ULrmyvSGsUAIsDpocdUimN+orYjc8bkYx2H
slR27guYhRpaa4oDsM7YK2o6gmcwU+0HNiKS01nHurqxiW6frvP5DyYPza85u1mmnAG2hSDEifEB
7qQ62PCK6MDx6uzsSlEpMkpbxXk3mni+ZA55c98BXnsjWoymLmneRCV7ROOoiXGJX9y3xQWpbt4z
Zf+JInIP9Q7K2d7SjXi3LaTnP0JqmoRlpbb9wZVybMqJvc/XXWkf5TQyk1TP3hfKFNH7F2tC1uIg
qrC5lBIN6Zy6K1VgfoDpCRiOaC7oLkRhSp3FiYqmlSMyzPTp6U/YrdPXIDcJinzFwLUTHoZ+h3tJ
1qj7tT/ZBtmptbP/SKMKY4+cGWJha8j3sA7qQ95qya9P5cX+uuK4XWMWef7nnqoTqmo6stmK2xgJ
WLEN6iXQ0/eYN8MWcKrGa58/Ej+cOWmO8UGnSECXYDAFGZORs19jzqjQrEO3F6gNNT0smHTC+Bbo
gAXic2cDu2A1Km1q3w+g1i0Y+vZhW1sULlThRYKpfQ5/8rg0zS2jybR5pvu6i5SJkwPOESm4ZFff
11DvJMjEme7VkpBjhuopcdYJkrbTpsAVLvgn0CVeBad1hWbHEnV4y2Va7SQyHUPmxLVEklYaaAxd
lYnn+EXYZz43dnujJ0+uGKchoNrFbDWKNKCsYJ3NZpp9ouOMcSyqtzu7NRpepcIinfE5qraHh3Ho
nzq3gnLxrzflMqBZIoKZG959/7qmmrR8y7zk2LqESYUE55zOZaQYS1bFCC4bsMn/jDqI7F3msTdj
/aA0fzHX5p0OfHR9CSWki6CKNRmF1RmcCdn7p3nC3aL29FefgFVa3Y4q71+RSsnFaDWglvobTXZW
dSc0fsMU7+oA9n7ma6sSEdibkR0E7ylb1M9Ui+TsS5BxW2ZzckgZgpqLn/L/1fY0hyHsJjr3lMPN
zx+u4kqBfSoKUkIeRjTCi5//zmFfvDr4k6o8dJ7ATHo0IlvyF/ldtyFekeFxAF8k9iPBx988pJJr
3ggX5/XBQ58LnY714Fppp3SWS4oGnBXCERMu7m++sFGkfJFDD4n0DK9muzWPXcfeU9pbVJOGrMvU
7NEuBQVdUdboRjLeGMb0vmOe2ePhMgwMa9xaeYCtAVaCPeCS0Cn+JBZA/a39oRWTtPwkEthACw+r
l1g7WT7sbFrMt05nXHGdEph0uQEnRriBjXkdjmfL1Bg5W9FTnoJGTawUuhAayXtWBI6QiTEY+b+Q
IIEeuWAPem2Yb3h8Z0Gr4PnOZBc2wcSveTfM77qPF7IOQqxy6AtD1l87vmMCXIbAQg2Vaihtcf9W
+NzOJlQnXA5d+Nw2Bbq+DpI73iv1+J9RX9h/K1o1IR8MBHxvLB/gGo0gNvo5lKHzaxvJZfA8fqCH
gXn25vBT0jc7PDJEtnTfS9wHcBV/XB71QkAGlox31xuZ/Sj/mDzdMqZ/3384/bHSou0xto5L57VI
EWCaIlFzE82on9lXTP0UPi3UanUjYS97K2lkslOsoOUivd+GFwNxCevn8EBnedejIvdC0n9Kz1Zt
Pr2Eu0kPy2biqecoitYcrRZMuiT6dQ+AFH++KsOrLaBJkJeytho1BCgH7kZ0rfLa7Ay28qvrHP9w
yZQvpf+10Ude3E7WweIdhDYC0QGp/Fa2wol48nEgbxa3Gx/k2+IqrSEhQXDm/av5Cl0T25N/EhWx
Fj3vh8F4lJCT1VNCoSWYNBfgcSQRuQtC5gqO1duiy17RWI/g7oSonkgStk8sU0AXRwU6MOEKZTtA
DeKcoYyDAK9R5huLYChpAt42h+kBfJnKdRbgEk7jy/awUZxllpFnZFHiDJ2nPd0BXO6EJJ84JYpO
J8ykkSsxFlLhfUKHJN2VwN1rX7dSL5hUTtj0Hw9wDOdfxszNDiBJS7Bl7XZKwFQHYdgF5jo1pJ9q
8v4nVbdQyLPEys3M7ftJfRtaZXqz37MVXzgz1FxmRpj+MZ3tOgVVtJZ2me4ftACG+KGddu2Sf/pV
cxoEiPO1MsBVQlSb1qyGuicao+tgQE6G4kJC7SEEJOi3OSKIZIzbWyNQ+UfunN1351jp4nLYxokI
z4gZ1JWv6MYPdCbPUqUxJJv5bMLJTolomnsO+S236MkaLvvhYH8VsnTQGDXaWBjIXDPh+gvJ8Hv+
Gqxr2cjec1Vvi+cqK2e2P29gqCC9g7EGnDBP1kLPQkS/4OQL56pCVRup4voZDGWaHLNzDlWFPtqb
a704VWWoFWbVvMndTeG//lTD5Xnqv3guOJsVhrrY2FViTQUFPtf61EypItWs0az3Ue5NcaSYUMcU
sAAp7O5XphaAhq8SJDzbSEKTuTd32HgT1JrJ+MQVaaDxK0EskSyH0gfydoqWKMtwtRhAE+QkGXO5
QOh34FpeWuzB6MaQiW1tGqvM5W4U1nMPERwqSH7ouWtA69C8zTR+CRyrxeZdM0+PUzF0AKqD/qTo
v3nZMJ7/n+KLShCM8FVKKfWeqbp5wdx8YgBw67v0/XKHTqHYs8OabWW0jX30+CPA2PTx7yYdTSge
M12gWRERRoR0xo+1g5aoBfRqVTEt8RISYpj7/D4srtN1lof6xlfd7bnIrqPJvtMmFhdkN4n33k21
J2CjSrzk5syhnwqSs7KUjaV11vzWjO4p5nxf5+s+niR4fNZF7CZ9RfxsMhvDYraKlFRTv/vCo42A
eGHh/x/igbQh69H7sHwlUp6THZgAGpfHKizur3yInzz1V+qQI+94hGcVlwqSuK7+ZJgoM5qzWJS8
/GOtxzbBgA4FIjxIYe+bL/u/xC/sa3K4ZDN6KwlrdF9JjXIHC6GPxdFa4eqDQs5VkEUQ4VKfTJ3X
NklQYlyukvcZ9VdQ0tVO0Cb0qfS2BM3dWGlmUvZrgm0yvwmgWIQOlRuaQwGQZOfAQAErqbt0z309
oGWFeFA4LNve47G/mS6XLp2iB3Vf3l++bNjy7PQ046SY6lyaAkM/XSOHKn+Lm+x3srdTFutGfqSM
6d5eRZ5wTytu7yPoX5Aaw6mY7dm/WPYIkxRyLFOJaHfj1gw6/ejO2EFQZXLs+SmfZZRujshFQ+tV
Hv2lO45lXZmrgXn+Zpcq3VziRq0UYw6PaW+oIKu/vKdKihlaDINQj8IEB3NfRdjO0N6ddPmaQFR8
NHs63laaxkH4gIs3iVVNpJLe3OkiP1ao7Tx44NpXmtvFTJc/HGyWairMhjEYZsn164flXm3UY+EI
4FxYA15IVBHqt77t0rE/5ql/ocDv1Ee9U+1GLgNGW/F3xxCmd15CL+73spZeML3LBQIPKB61TiQr
at0TYh0ZHYF6ctnSIR7esQW+h2z2quuNYY0DDyF5IVzmHqvYOC/Rj7BJ1ckIXzhSjaDM3AW17qxx
ox86ygkyQCjrPKRFh/RbgO1sx6M7g+hPXCzjKDYHR5M/7O17cZwE9ffb6E61wxgDhY5fTh7XA5yK
kcotlhtBVQmOav4OAKJWF9ewn/DWbzeHab2DC+s90yCCObdNyC1aADnevJIHASLmES9MMZTA03+z
0pVKzfDUlQLdPgoCB8LlkHDKq7gLTusf0BI2TWxLfEdgKZRUCb5mP91eItccYpgcUgjzUhz1U1G6
aTegjEXl1/0W8dqSoOmHx9G50Cep/pZtgBoMZwCj78VU2PGqjZmX9m8LhIIYd2kTkTVE/O/zuoa3
brlKuO7e7F/PyB9OXK4tinHROcYEFxdQ+YWdtZ5Tvw8Bwg8qPxpmphFs5wFouKyBSzUmwi7v3gSR
hUz+Y20t74eBL9nxToKbi6VIhgnGCAdrsbW6QQ2jpkTnd5a+S6INONER1Ws7SbwJ9Z5dtjcyhSWw
3+eTDyH0Es2ROUK5IUSnevJYxJSt/CYZ4UfN1WRf8g96y1KjxA2x+Xbm/Zwigx7r2QRrG2fqhon1
cVjlQnuvllAjIZ0MREYEsWyAIgGQSl4FZDKvLgn40WvX8BPgMHHX3Xb/6S449g6Vmu/pqSLhRT/T
ejn+wt+sRE0xaNvOS897ovn1SR1uUxiomZERCEoZry1t53jZ0uVj2lfCQvsK7CXo9QQk0mhGjAbR
VbPTjfhQ04IJPYqWa+XSpMo5JIW1QapjObXj3aAQghVkO4hDhNfcDxb1qyHDCDK7r4rrmqhv4eq5
cvF3/bq71Y6/dejU9AtBFKDjq8EX0dKZBsCfoOTG25Eglxqquun4hGFCxOuGCnFTtefY3es0+R7C
q0AbdyOnOq/azDGe744SJqL7oC2pO66nkqwBUrUS721+ezCLfGy0a8mDf1ii6teQSXU35as1WOQ/
7hucz89xLfRkpxS4EkmB26+3x13W4vw/3xmN7J2d8SjgtoduR4hV12bRGQqKxzCoqclpnHD+dMu9
GdXEna7lPz+T3Y3kpxD4AlmZsbEHvNv1mscA0cZxHZ4HEDzX3zvRBcNsmYTtpf94PeGE1CD3SD6v
b8ppRAD1XeTvx3JfE6n2XinrCgjdjuzFPgJwqgcamIffYqUroQjeyOhaEPZh/aup4Jff9aBuhJPH
MwhQitV7PKHF9o/cF9cKWMG/ifgkAjKNfbuRO+9GgumGUAB5wOOITgc7PLsfeHLeG8ay/BNySw8f
z96ywjFTZT70q/FDK3zBh/qYRUn4LS1Pn+B1lpaFDjGVoLraB2BMO9rwNFVhYWm0+hBFNiTyXSxV
cY2mMpzV0XOwNATZsYNIHPCAVv65Chb/8/txrHlNe4XEIdldCfE8t/E8KpX7hPkTXec4bZ+N4Ryt
pEg0RJX6zgcaDtKKs6DDRaJS+VLkxclGUJskME0IMxYNg+pJcg/pOZNCg+Pk9EFZhizPQOVusmvl
26vPW1bKeSCsjHULJwNxdpWrRy6eA5o93hX8kuSRiRz3DJ/gXW0y5mJbMs56HQNIPhaDCGpNeKuj
ydNCG0GonaIFOhn0AhrIKmdf4c9MWlQ7h8nn9+15wystym7ZQCzkRxujb3/86CDImeu4UnZRssoH
0aVjRs/nUiUBD7HS9Siy0gKUN79xQM2wxsvy0FL9QIrDYWfnjwBA2+rUhfQujmqoBGzRU86z+J60
Po6uYunAX+iyKZNiyk9cV9IBe1G8FaXLo3wdTZ3+6B0KWvS+9+CGaM4j+bvJhAbvseQDcP7kfod8
YmdKzWRXuyD3od1mCLuNX44vSto0BIKcykJLR05/vpNio1u/2+f5s4HgAn5bgEFwKlspFKLk2a8K
mLyxEVZ9z0cFFIIuh4mNBj1IbcSO6kdXhfKVbOQebjNXw6Q2RE2bmZgLsKabqykPqSNKCwYYsViZ
rOiBRtvm9MV5WrizvrXsVkyMBPHDzlNZk8S7NV2vJg+fys9/Mv4sier+Kl3iN+Br27v13nSvAiAl
vm0gyG90GikV5IT20APJj8yiXavQv2OG5uHGJfw3At+SeKSlDSrb3wXrObtcWe6tzpWJDGD9aFCA
DwMctzOkZitRG9XlP86Aw2P69wN2YM7XAip7VZJvgPFUC5T519ubo7VxCQge/1X6g7hjT7R58XT4
r6W2U7zJEIEgGJqy0Vl/7VFnunck8vebaUAWhSYXnZuIioYkcw+GKaycJi5ERRzZ4yvQX4WTVc4M
wBD042A2J/uxNsd8A0ozHIDUehIvfhoibqBq7xzsoiW3MYmYkI8/ZjxBX0a5idKuLISfhtoHgrnh
B+MX/aOMXvDjj7x0hWci/HbYIjQWgpQL2TSlpfP3voP4DJF2r2oX7Tzhq5mBLwu97Vln7Mm7rWCN
4Hn2X3wZdbZzMt3Hapx7+ju3h+vVCXJEecRELkIXYf6stAMbhZZMZlxLQnTukNb4vg3N5fHYvc+Q
w3QyIsmB2QYdHQgA7w2rFGMlnnMUmzi4NOccgQVt2mfocFuiuFl9X7SRuZxzc1As6qMBVrXCDQdC
i+4dkWKl/KnKKHw9qwKKJwLygWISo8Nd8JC24rrOdPN3P7+5r4tRRzEyr6XDoplIjSNhy2mHO2x7
ryGpgUKj0sN/XOVW0YVvfC4Cj5SXz3T5bxLntYS/+wMIJM7n0UovZjmqqjpCSyiWaZ6NcoyrWu2i
aX/b4fDBI8rkL3C+3ZSDWOtXFBMbLTLnoWWBgASr534EotIm8CxvPoy8TDeAdHEqFT6b4yz/XlBk
hM1EzYCaOCRLj9FqzCkeUfyaEeQyTkJP4anx1TcQYwRzZ7CwxbDP/XKNUe8HjhBc0z48JBVAf2Sr
QKTWKRIMiPul0qpFKUvkvO7dY1xjFfqUEKA0r9yugtKlsP9hxNOFAEVVzMKck54MnxmHvNVqH9fU
ANHB9EVr6nLNCko0kmx7FIiKHrHdMl3zrmq1sKSs4YtuQeb2UIMHN33eFuEdHz0opM4wTLysvgCg
05b0nM9ltXPvY0hXHqkAd7rUyVvLWTsygtLIiGc+1PvzeQH60Op2Wk1TQgtXpQc8QhnIWeyDvM75
daVzmvspDUA8SndGbXUVQPNHXJzrKVoie9Dzj2YGo20rotXjBmoUQa2v9inkxlJDsGjju106iiP7
Fj99HxNWhEpyRdQ66Zd/cQxgBK0RF8R/28z944X0KFlRNJhB8lvrjzJyK9nwF1K/PK8PvuLwG1AE
s6hf018UAeujsW348L9JQ1/Mt8n6LBxf7PHGoBTg478QBeLAWeFcMVU7eW/pwwWoN0fPrGzYPCEn
sWINC9ZTMxkx2vsqF2W3+QOOVGaQFQG4yqDgrRH9MaUyYpoCbtBxZ+uReZuIgpAf4OQDhrZLywxL
es7aud9FHbG4LrgKJz1ctxBunfWdjRJ4lLMx+hCsh7JyA7r2eqZb9ShPtZuiPsVR9GW9bhHf1mrI
9XfrpsuLeO2p18K8/ZXqpkaTE7OFxTHISvwfrGNvugpw4vOJ01XfTUGjk7r+ysy1kgF/kcq857Is
LYZhtxAAWyYKXoal+7cE66S9zTJXMYjuV8Z/36zIXho3KNW6hvN2HjGJc8xlcw/WBnQD73nuDefQ
lzovv8TbQoYiyD4GF6iFd4Delj1lTouacSmzYpfEg3AwMXAvTQlEjI8iWlOFNSO1WPmCEU8LcmfP
OrM5OfZ30hh+Fa1G1KQrJfXkZk4ZSCTalS8JDC8DI7X0bHwLBLXO7x6rCaPtqCajHHGlJmaGiYKP
tHVLqLFKEUnYSVJOjgDADqQYsdZgJlGguAA67XsgG8UtPr3Nmdcr4naWokiaI6Ncbp9AUa9+bS5j
EJ1/dLai7TN6eNPK30r7czrhws8bwD4G9Cra/PO+CqDWzKOOpn94JEdJrMKJWVSw0P6I+XCdQ22i
Bk0U/ZsZVWwysS14+CHJDCIBUWX29znh8PA2uqFYn5KPbi/yWx7QNGOnDY4t+Mrba5sdmsJXj46d
VyFa5hOaR65PgbwoZt8QwBHjERCsoUx7hFnmHK114Wss1n4btfljT10z65Xjq7sBfeWZFh7NcRY7
6vZPQGHGg26NVEYYJmIBVHZnyKRCby8LOer/jVo17wYv6VyeRuiPfl1Lw4smYMI9ogE/ELrpaPnt
frU6Y13KPyni1IeKvzQEf7UpxNCqYRX7+fu5lGJn3c3nsO3J9Yl+Cdo+oqHrIW0b1jf4SGCfGgNj
fGjOvMzz7zvbtHs0U+IuSkuClBkKWMBHB2JSzhD2/TIHbhNQr1ub3lFzg33YKn8fhi70ObxMFDPK
F5Yg2jueqQHG7tBJG8q0+w0cSmUsGhnXi95mgJkSPXRZRbOzCbjPcr+sv+pALBuQ6PoPzzjt1hhh
L9/Ee8GjqMz5sky6OpjghBG/BYutsnbzWtXenErl+kM0yGRnxgEfA5ng0uHaFFoMnrPe9hN3iOuY
zWmVC1Etjs27ICV0R9FYMATOEwZxu3sX2N2AgP8wIANmTR6ngUsh2pdbghm45Gh/h0w9v5p14+yh
lc6q0CXbdSs6NxnNhN9Ky3klFB2gzSN3Wzpi5gvMCIsWsmK0TC5mFic4ha6fAH1Rj4499/hA60FR
+Iu96KB+vH2DE+FWFIGgWMMnms1fCbW99N0moeagCpqeO3I66roVottiG90uvswbh04A4bin1vr6
XeBRzW7AC3RRzNCVHS0XH+iRDe54c3YsjhH7sr32MpHDZ9fQ6x+PnF1GBAO0xYWl87VJJuvs+VEJ
ycZy1BlDGRvNct+hsgXMKUl6MxFC5y0X1T7SaPQID9pedw+50Nfi2XkW99v8PjKYvTe/+HdU3jaQ
f+8fKS1ZFWTqqcDpTm2zbZu2RaDJtlY71OyV2Hp0C14jsxuVlQabk+zzW3eUo6bLk889QIe5Ttli
9dLE23ZIjp3B+rfymu1ZRRjJa1+YawqizJITd2fmfCDdX3wzJvYbXUuijRxcnVd7AcubWiJwGP7y
WKkx2umwnjbXHCiF99RyjzKi+DGPYc9U0Yvithws8NKGKzxqtCDd2vjhkrfljkB84C4Vo4rnHVkz
uez9WhO7g0HywfWb13emedYardQWG1+BKfT6vNU1G3Z168ercSOg9gw7DGjw3Kk3xOD7mQCKmMis
negEnQaPv64Y+iZuUZNTOOtIB7ZSMzoe/fE+fDx8aP8XOrqlVDyGM2wYb+WZSA+NX1TSIEmostr0
QHrzUMhIrg1PdhCrK58UD+1yVdr5ubpgtRX3p2aDVEpRkk2tuQTXpsoW0g8e4D0zKFkQjDfg0BrU
gYhctV+VJzYDoFHE1YaQI3GcCidRbbh7nuKvv+Na8uiWGvCo5g5nPG7obqvDiehU2EpSXLIX4TsS
XUzpAau39uRwkjlPe5IqtJcQM1OSBnS4R7GdLgq/Kgvl7i09sM6tqVV0IW7YOAQaIyi1LvW9gN/4
+AJLNtbJTyHDtaSsygD1XisawglgXYHR4MdF+G0MYFdG0spssUU/xP/OmPQjk+Nsk5s9j45JACOM
lW4kChYPgTdRQjT45Ubl8VDo8G0r7hmsfdRVn8PVJol+V2lJ/AMBh6mCom8NFK9uRMp5dVzmcWZi
EgRtQqrmLl3i/xdyppzw9G4Pbe+Wlx4+/gLE31Suvqxm4ViqNdx22fmT0gh+lFz/SqSON2OLwyDE
XYSJQFn5NLH+LzLUeRwIC1+bCZ42B316plaPLsuP0OSg7uZlrNDC1yy2ApPJ6E9QoJe5AktIJPgK
XFWKOqurEzHltmopvf+CaN02bm7QOhjxWx/Nx7wHyIvahe25YYyq6zDPnY1hadvV/8MT/GsqwaHD
JWOvssolpw1OBHp1BxKebk5USZH6bKy/JV7i/9eTFA9dM94uLx68yQ/o01r4GhxI88PcY4X4B08p
/UmpQsfLwVr03EH0cUEQhINR7pBBSM70dykR6ZF5KpL7WQGYMkY4VEzZ93TTA51JyUgs16hbAc0p
UN3QwUjOHGWmc9z1zkgyccVYyaVPSGYSY+ItArBFAskNiEXnQ+kRluZhKwdpF02MVaSvaWhv5ULV
PxumDfgIQN9W17O5p2QnLoidAkOth3pLZJPs2AV0hih9Y/1VtorU9esaqPi3YlJm8VoEdfYlKlGT
GM4EVCI++AaYE+ioDyDCUcTwLgpK8uG0SL2fo8YXgaaR39Ad5Euxj9lGibraSUQ5TkLes++m3Enn
3JjLtD8gKxz/hpZW+j33nfUThvA2uuj32pp7hEDBzpPivks2UPP4DJxgcJUEeH+1kMrL3ETN4GUN
2Ej3jRBq5Ngq8V5KMCz/VIlNOHUUkOuEwYkvafoxXtIRnNWwoAKcr7Ble4oTG5X/iC8qb4wwVgKF
e9eL0HuuhP4IW0qO8eKSJHKYiaDdEIXHHT59xkK/hSc8UCnuYidWaxNCRgSEs5mrVj17cySmmnqH
NlKkwIBLGAxkQ99KYK5R725tiD1yeS5Ky8elZKcHnqtgvPDUmyyYlYj8nJR8woZ/iG46srfjCKQY
Do7fbjThJL+5NVEg6ompV8rvM/+QTuvpDEPnFQdUh0RIzWUt14KxhL7p9trJQF1ODOGAuZAUTqG8
7xznF21SeE+9IKtNru9ZxRHpiWUhdhN0mkFZ3xF92Zzg7kmHtWE7TyR4A/LbCN3WlW+4wjZcc3YP
n/LPJiNVTUwZ93qmLp9utfhIKDPx1+VhWNiH0wYqxfOs85Ux4nbvB7mVs+9nCoCB5mCm2H+wqOtL
hEf+pAQlMk5Mb+K2jC2GTEpc035mPr2hL8kfaAOwMIqs4/4AIJ2Nl6hn6IbIJlBLiYcETKbF2ofe
2vsHd9Z4OlDqDkXJwzZVXGTw/YHwosrvKrkE5B7G4Yh1jEKreqIJtLgEaWRDhB+szYd54vqONLXV
0xR1Ggwirh5kAqnhNEnhlPnRqVT1qBtIu6+oxvGH/5eThilR15QhKjmj9zcXr9ojgMqTJREG4+Q0
IiucDXy8diFN0NFndxzmOkI45KZV3zUzHB+j2ekhRjvgFbOkKJRsaMGVFjfxx+fMD8TpQj+PnSu7
tjyerURe61mjonSz6qKXDm5RuU1WIjidlS7wwNc+P2SlmQSUsm2CpIMSZdZIGeYmlUJahPKXY4O2
cnyKSleFHcxMBu8c29+bOQmrBgJk9P229mbSFbtm7HZtMv+8S0T1OOGS4BDxI+vxLRUz2tz5jqXP
nY6B6M/8eQ4h/DgC9R8ZWjGiitpzU+IjQEeDR8jBEzGTiBugt16LxWNNV+YCFAsaWqndQ2wAft5G
R1gDlAVO/W2OZfIbsnBvF7gCkE1S0v0QSF43CcdqM+wthdE1YqPNYu+lfIPdPNOoedx+IQJ7xuhM
hNoAhwk7vjVCQ5HSndg5S4RR9kFnpkQMp1tsdtJ9t5y2o2bStr5apIIZP09tiImjGndK/IDR4yYn
WvEFZUMNNyrGO6tuHAbPYar5uhLgnppSNHgR1u6B3r475a/vucmuIHdm+KzVoUAO9+5VJZgGRz3m
H16KEBmGXO4XHY4rOh4GFv5uiHctKmjec129CtklcgTgFGEXbedQ5jMJytaHAQyGdAEMeaF1fv52
Vsh2PcxANrQBVmMm30oaEBkxj7GFvDqIzF8xIQrWdRr9XWFC4B0ng6+SBPzW5cBaK0vSrtzWXKD2
Kwbqq02JhoWtNpiW6EwayCnqFlGkYSR9BAwYqi6RAJbG9Gp5to1sCpYPAVYoiM1j03qozYZn4nuw
AQwFrnMHqVTElE7YdvuoJJLNn/xEXubA7dXzK0oCNvatnUDVWSiaOMpMZwLtYSXysgvwE6zq9w18
g0Jd7IFJfjoednHxduk6TDmDrD3GQMBkaneEKhYc3VmHso7LTr5lwIAg1QXM6AVEzfa9Ucdb+5cb
rm93qvWbug9sXgVqKAwP6WIcqMlllpQfSh8Ee0Rcet3TYYlnqPnFdI+4ob2Z+Lv+RDRxkRSbkN+O
GlLYnJRVTKDe1eoqkfnC6vCcYiUX+Wo8QDjajbZAWp4PhRTD9AyZkxny4qArDhrfzLiuv2fCLiEd
IMvJrcA7OL6HNCc1g5KL9Z+w7V3Q6hNxShdyNdfVdwCR7XhMToEkRF24qUW1ZyLY+MMGDTEFezem
4clpR5fBNsAxF9xs/dXqLQbddGPGPkkQ0nrqRGlQoyl5Roc3VOiyGpdvuZviytRwud8mbm/K8X20
oo3/ZQI7183AvR6ZtV+w4IPpTMG1dycAh8dl7aLSicE98fFRww2EiKDX4AalyWJOoc/nYmDyUOGC
pLWNSBWIhzlRda58NmD8qIXvWXe26ElG+JNDSeG3nPstrZl2fEIm2UPjyi7mrxGwvycPWZPUNkv+
pVMs6fmp3Wgns17g8+wnG+GJ0VPtgDItzr1GxRrSbnQbmXtvMLHkybQwAeAySIoyfBmGNhOfHYcR
eJAxXfMpY1fmFw1Dv0SaBp+jhD5agSumOrGzwsBYqUPLJoKNDIgz9H/696uEUxinP3r1rt7t8crR
5rnPcRcWzzvfVs72akrcXoUfAXjGpCrymWGS9yN/6myqyq+dyfvoVkDnoa6IQWxQyoA0N8VEvJQF
RXdHh4QrSgwcG5OKtjsOyUA28DAkGeF65Moss3iuG2Tcim08bm7phfOABa8b0WYPCvD82hUsvv8J
FCuElVkcEdl+tATQ4Z2Zb6TCzeWg4xvQ1tjwgxF1eDLVktUQ5PYUZ//GylPqy9Ya9ZE8jm+SWDxs
e1g5Lp6PgPYA4YadmmUuTX4fCIb39B4+W4Um4KwQ8IgaHOhud73gTEOM/dD8RcM/N9rbLWog37cK
b2NRoLp36U334if9Ke6bfFXTQPzVs9QW0GvCsCp8RNMq/m0FLefzAFf5cf6gEA1lxgF8A1vhdAn+
eUikY8WePZntZIncoc1CVhowGNOt4c0nn2GAB8E3ZjQMWhTiDjDFsEKmPfbTaadQjO1OMU1sHHXu
zMaSTOtVkELK6m0Y3e1MC6RQrp6LiAPWW7FMxHeuuXABIs9joHROSNLD6606acYpk5s2tybw+l+7
28C+mvT5F1dg7Jqydpb6T2A38wzrwXQmUn4I4ccPI14APFKkpMXgAr+MsehZHeOrIB5Y/4y4T3/z
XahkN3gLfL1UVFC3G9tPhwrbV6go1LhKxDMLxCOwjeacfpkJoST17iZl1qAdS7/HKeXvL7VRwJo5
xsDW6HCeqljcV9jMQDaRa0PMIcjrnLLwD7XHncANJA5uPmdMlNXmuCmVvJEUfRgrzz8Qg3tyCda4
zcRB3D3l6MUSHQdMgbyTgoAFw0xPQ5sVNcZL2PY7tH/xW7WFyHBRsCc5ckfwrTEPGiYBrkIf0EHC
uqgJOC75SuIarxVM+VTcUJ5wNn88L8bjFgmtyqA8Olt6QlVPZjwLzO2WS3A1e16Ht6g8fV5OoQOK
aG+OzOGhYsEt9OIgGNi36wx6gkmrbnq8SEkLcCN9W+BBD8LnLL5/6D1Ti1iXBNb3JTiL1g2Qe6/G
5n5XsLofc1czfxzmdhEFSYXylOiiurT52wT+PT0F8a1HzCCHxeBKttbYtaW2ORLLpq726Mc+zZ2K
BNUQGM24x5C1n7vakDZMgrM6EWZWPGUFVk/THC5YNCyqGcBCcfn4mY90lqmzMrsiFuTngThEJFrH
NeVuZu5g9ZJLMvatf1Zw4KxFIsNtQHtIi9ThbZQzW70IwG2ASxjM3dPHg2MTdKpIMremsVgh6J60
Yc5uTqp5P6AsyuR42nuoxExEG7wKPwStnp78orbpIuPBTvGYCfu5IMw+Atkv7h/+SBBBnXRWN/B+
146QbBYjH9jqaINrOgKiySUQ0rMRp9yaH/3xdb+EW2IYL8qEJ+RFIl3GAB1qlDDVhcXEKt0YRJlA
h0w3WA5D/qN8847nhv+T5+fjWDbYLS4z8D+3GcHdtRn5jaVJJupqHx0BoT63bZ/jnB1tP0Skboys
p/jvtpB2STpG0h2f3JWn8K9BNoWaVJf+dF0xjeqiwbMzzcS1cn0g4JQp0GILnc0iraxU/alOYGH3
ybN7BBISHVDNuth0Nm8zz5ptCjVaIZPxC35kRQscLyPrOwlCTdK8l3ORmfiLwsIQJB38towemQgf
g78Uz5Q/Hz+TKU9NSOFolDXERbzcwmyGir3wByG7yOmGyiZgF/1ckzEi/pXJLt0aVsgAU6iSDhBd
Yo0MEm9Z35LqAOtdpWtzyQ80v4FM5kdgKcj2T3VAc3BgrhSr4GB+ZxunrmtsdHcEOZOBJF3M683S
bofKmD0V3fqIKpWfYsq3axPnboY0WJetBAhCDW7FDkI+F4zcTHO08TIyIGme43mFcMVol81IS+Se
IBsMlC4kJYO4St7DW/Ok8GDutjLrIuQ/FZUD5u4lqQkIwA3O+9KUc/kFREfAT82Fo0CjZjJK4QZK
Pkxa1w4bc5W1zTOTPE7o/g/j4/PtDiP+ERyH5gKObUFKr7wP8OizjTTGRhknHQOqcvo0AD05e/kB
3nhpRvmsBMkLAWy2R/C40hJrZTukrcG/TnHCeTEBjt/8ZYD97g7tUYjl/VOGbncU/l5hFrhejD/6
GCokREOwgUtAA36n1PJdbswU0NTbcFPblTbke8D37jmECrclvNv2Ut2tBcEHIQar/viJn8FS96to
jUFsuoDy3o/P/zRM47htXGiSDTtMzdu7n0909J5MiuuZpK6GMl9T8DBsHyGRs2VvnZNEYiyRMIOP
+SChxT7EwrsRLJh27oq/9cbo8KO6CoaJlOo9tT/MYAI8vkhFDQBtX4IgzMzgaGldtKcC3je/nb7e
OQIOClTLVbDJrewWmzIc+/zdCR295uMOszv32lBuwg30S+IDrBxy1iE3oDZqkKyZ6tzLdj1znXZR
rWdXmvDqkty7gOwDxuZANhsJVEZDAMokgdsyFAiBiNnYdJZiTjzrt/sVGM5Q922YlcIb1imyH907
QPdEZLWyyHi05dXF1x4IAZXAXftlzfUp9BWva3Eu0sxvjofYnLAZJoTo3gp+Y3BA+9TgEhOACNnw
lkX/SXPXi4wNqC15wgpbEqRjJ5S1LqkUQWumVEzt9e5eyohBC4SHlVRWAVghzNcLC3pfNNCW3UcI
1gFB+vn45iTvWVRFH6t8cw8YTARt3nhr5sOCFzYnLUKkKoJpOjsxsws7mG5TbQ8nPvlpi42ARANy
y5FKJY+LMV9QyOfKKD7SV7SykkkoxC+Y2/w8CVfJR+KDqmx2n0jrwSLYkqml/o7WBqIYELbXYV45
HYTIYakrNOCDEKwfkmU8TAjE1mT9VHYvXMQvuPo1/Qu2P87d5fcyVHRsDEkxOeIOdpgq5XbuD+Yu
HS73H5FW3+inwqbecoBr/rhL+KnfafpjFvASfJm5viLs+2LwDqn6Kn+qz2fNHHDV0fuOU99M8bp/
G7iKeyD68hj2/mYt2SLWZSq/65Y+dlHShTxF3xdpufUDJMCr/YKgxzxJ1UwcriPU65lLkjL/XAxU
B/ITroVIbsZRzgMbQPRtzOvx+m0yxLDLkqe8h4z3W+iTsiI8F3y/w9xKI1nuSP7PXDJTnzADNFB/
uimLelPJ35fRmB6UEmaG81yfULW8gDDT4fq96a/4bdyFnLTL59qxAYJQcQgSMJGvi+V159SWD4c5
u9a/1vRXbmtJ6Et49SKUAk8t/lDCKkScDZV/kXT47CR4lP1Uxkq7We73qiPe9ZZg03K4wBmcZAoI
iCpdPCBCNtOwahv1bbMKv1HIQVIpQlW67zKrYARqEKdge9pgY6Q3OHIzYRYKIXVQklLwm4yd9C8R
CzbWeWW/iPdaSjsFHahPrFVohfaD/uLpHDUWFjGNJsXe6SkDLigZZZdi2tbN3p9iNa4pSq7KC8x+
zh6IuWC1wHzgPX5h+j5mimQVYXUWP0KEn40/4McH6E7ZLuIPYda+cnrbQ2MjNLo7Hap/z0xOfF8o
wwSQd8c6H/e1iuduxLIN04CBvafmoTXutuLx6lBm+Y+0Zthd4Xzw34lm0if6G3rvOCRXVTF+eUEq
x49U2VZ0UWUzaQM8YIwG9I6y/xK2ccyYs3OeQGJjywUlJl8bXa6ckfjgpHfd/H8gJZhtaXjOhfD2
w33/mln2/5HEddZYUi9DNWMZTht0JdmbI1mIiW9MseAlX55G3NHhCW8GVf2CLDZd9iy/5EvAR4Da
auZ3KeDhkvuTAo6SmdEh1b3NYvBo+jMaCGhHDXXUTICAvygW/wognUbYU8DtrTnvTom22w8mFrY8
ENsWFNIETKVX8MPH4pGKzOa1dadqUfWRszWsdGtJ+wSFkMEvWQUHdHw/ioNCziSYbwSR+eWegYrX
6/itWGjNd0P+39lAplBrioebKns1fMecF1XU3ViZkTCrlKg0UvGiL4G5/7ov54QXHQStAROH04mR
493f6p5xixwE+zLaFtoO8L+gN2vT9N0aMwclT7MqpPAeSHm1ONt3Fmc6A9Q/x7TgqxhMmk4zTfvG
7hDiY9vY01NXtNQiKQpFhNo/MZXDqHZyBglDYEV39mtJbFDZS+4Fp4a0LoOdBSoMzfwWtGWi6vuh
EeZ4Sx8D2QTLWSu124aY4wvVo89/vEa1ZyWG4xPy+1OQeCUrUeohHCGWnQdpw6uf4KUEydzzKWOZ
LHqd3wT7T8ffxfffOeabAJTLSVKTMSBB4VwVxeW+4numoGWTzR5ga4XZmlWws1ltWuNWUPPl+cz4
raFQ1YPVGpjNlqY1FNNaLs2JD7He8F5Y0U4niFyRQbQhp9bn+BrCDZ47Xe96zFYdrtpZdrv0kTyj
ImE/y9FMPtS20xr8Z7QXD7I/2af8UORU/oyarNeXpTT4x/4guPevKUipSaQ9mqU32WYj8egkdb3I
tQ1crQh2pHj++Rr5IBcotkB46rVyDEAgqQ8=
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw1n;
use gw1n.components.all;

entity PSRAM_Memory_Interface_HS_Top is
port(
  clk :  in std_logic;
  memory_clk :  in std_logic;
  pll_lock :  in std_logic;
  rst_n :  in std_logic;
  O_psram_ck :  out std_logic_vector(1 downto 0);
  O_psram_ck_n :  out std_logic_vector(1 downto 0);
  IO_psram_dq :  inout std_logic_vector(15 downto 0);
  IO_psram_rwds :  inout std_logic_vector(1 downto 0);
  O_psram_cs_n :  out std_logic_vector(1 downto 0);
  O_psram_reset_n :  out std_logic_vector(1 downto 0);
  wr_data :  in std_logic_vector(63 downto 0);
  rd_data :  out std_logic_vector(63 downto 0);
  rd_data_valid :  out std_logic;
  addr :  in std_logic_vector(20 downto 0);
  cmd :  in std_logic;
  cmd_en :  in std_logic;
  init_calib :  out std_logic;
  clk_out :  out std_logic;
  data_mask :  in std_logic_vector(7 downto 0));
end PSRAM_Memory_Interface_HS_Top;
architecture beh of PSRAM_Memory_Interface_HS_Top is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
  signal NN_0 : std_logic;
  signal NN_1 : std_logic;
component \~psram_top.PSRAM_Memory_Interface_HS_Top\
port(
  memory_clk: in std_logic;
  GND_0: in std_logic;
  rst_n: in std_logic;
  pll_lock: in std_logic;
  VCC_0: in std_logic;
  cmd: in std_logic;
  cmd_en: in std_logic;
  clk: in std_logic;
  wr_data : in std_logic_vector(63 downto 0);
  addr : in std_logic_vector(20 downto 0);
  data_mask : in std_logic_vector(7 downto 0);
  clk_out: out std_logic;
  rd_data_valid: out std_logic;
  init_calib: out std_logic;
  rd_data : out std_logic_vector(63 downto 0);
  O_psram_ck : out std_logic_vector(1 downto 0);
  O_psram_ck_n : out std_logic_vector(1 downto 0);
  O_psram_cs_n : out std_logic_vector(1 downto 0);
  O_psram_reset_n : out std_logic_vector(1 downto 1);
  IO_psram_dq : inout std_logic_vector(15 downto 0);
  IO_psram_rwds : inout std_logic_vector(1 downto 0));
end component;
begin
GND_s5: GND
port map (
  G => GND_0);
VCC_s4: VCC
port map (
  V => VCC_0);
GSR_30: GSR
port map (
  GSRI => VCC_0);
u_psram_top: \~psram_top.PSRAM_Memory_Interface_HS_Top\
port map(
  memory_clk => memory_clk,
  GND_0 => GND_0,
  rst_n => rst_n,
  pll_lock => pll_lock,
  VCC_0 => VCC_0,
  cmd => cmd,
  cmd_en => cmd_en,
  clk => clk,
  wr_data(63 downto 0) => wr_data(63 downto 0),
  addr(20 downto 0) => addr(20 downto 0),
  data_mask(7 downto 0) => data_mask(7 downto 0),
  clk_out => NN_0,
  rd_data_valid => rd_data_valid,
  init_calib => NN_1,
  rd_data(63 downto 0) => rd_data(63 downto 0),
  O_psram_ck(1 downto 0) => O_psram_ck(1 downto 0),
  O_psram_ck_n(1 downto 0) => O_psram_ck_n(1 downto 0),
  O_psram_cs_n(1 downto 0) => O_psram_cs_n(1 downto 0),
  O_psram_reset_n(1) => NN,
  IO_psram_dq(15 downto 0) => IO_psram_dq(15 downto 0),
  IO_psram_rwds(1 downto 0) => IO_psram_rwds(1 downto 0));
  O_psram_reset_n(0) <= NN;
  O_psram_reset_n(1) <= NN;
  clk_out <= NN_0;
  init_calib <= NN_1;
end beh;
