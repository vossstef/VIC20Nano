--
--Written by GowinSynthesis
--Tool Version "V1.9.10 (64-bit)"
--Sun Aug 18 07:30:05 2024

--Source file index table:
--file0 "\C:/Gowin/Gowin_V1.9.10_x64/IDE/ipcore/PSRAM_HS/data/PSRAM_TOP.v"
--file1 "\C:/Gowin/Gowin_V1.9.10_x64/IDE/ipcore/PSRAM_HS/data/psram_code.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
h8tPCcJ1E03+nzgm+FM9FxZfwO/+bm6hqcf+bbahfDQ6qsmrOfLUHXn4N9rSAKqtP7dKEj7BnFH5
fRkCyG882rEfzvjw6IpEBtf5qZBfSpatCv13ZI8HUu1DqjNszHWCYXt17tmgVDfOucVRNDWJU6WH
BTL8pBqEPP6Yd1zT3xY76ebgNokqiffCRRVSn7i4/MydIvDcgZUCjXdjyU6ME2cSnb2ihgxKdWiP
YJuC5CykQMSVT78I39P7W85Pgf7LE9dwnkO2hlGbYXSQdxk5PKMyJvwpb1vJyabG2TmPMM4105h/
h6yVw4KxzES2XW7aTcAKjlTz98EW6QTDIY8fqA==

`protect encoding=(enctype="base64", line_length=76, bytes=310448)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
RlONMvlwz9n9vxyIaj+A6rtm/2/kJabTfvb6laHHaUPAvzStb6iLBIh25CRxmNxsEZIydPFk4lVR
skz7mNWkcbX72hyuHSg4fbqledRXRq3J4l+Tk6zlsOvPyal+L0cZJe0l7OpEb5Q32AOBYvN3/0nu
JfsCwxhV96IQXtuzYIZmRh8UsfvYSDLf+7Er7AcYhPsfjmVRZ3y4KmsciPi9Ojw1ZRvHKW0CF+Tx
pEHK5PDZd0Vtge72xwuuv8YZi+lKsEktuCs5E7BMKOYIIO4DQGBimIU4OA9Hl4Wc1eAgYX5/AOqc
TqLKhnkLMcsCZzkk3Re1l1JkTaqUvdjz98HNEkM5Px8kw8BNVi+zK2w639VYm8R9C5HGjH1iH5E2
ArwKNLcNUz41QAHUaYr2EmBwr2cQqDk0lzPeV58QGjSAqbMhTOqX1Em1twjqadh/6QIb6eqZxclx
6h68KVmWBAh87brd6b/JsegNgOC2nrpdmOGF+4kMJBT0BOuX2mRb8uwjbfK0JkUvMIW0v/B0k788
dk27AuUioQw93YTe1ZCOImZ/MIiKJRux//G6tHFSctcqwkVfl3KloSygJYK/nEMlw0+PcZl0LRq1
ePBoNsnpswJGswJE1pOKZC1baJ9OXvnAYrO62lz8gvRTA8DTlTN9xE6PCM79isdmER0vwUTAh4St
b3ddD1LiML83zroKWdl/SxJtbUD6vHZODLKbFd7KJhV1s1ab6CYmtg7iUo6R7wUwsSmuOPK2gQxm
AJtzpOWM+0bNl4Cyf+miR2pg8NweFYWgZa0c1zRJ0S9SO7NYlRwsSFiPG8KnLun4nfwbpynYHn0+
TfDb0BoyhzDxKQaTgCXBHCjVQYfqeO0XqifJh4vulDa30lm/VZqwIqFkKh6+nDx5GFvFmB44aD92
tV4bq77TIJOFUvTrlpNe2Wmxo5mbFV7nwJw3ZFOJVsxSKe8kVUwP0pSL5l9+1Ck4P7pMK9x+iQ8E
VQJAQI3SMDI2866h8eQE6JGETx9yKV7VVy+Tdq4WR9bQcBW6QAO3ZiTF555lgWJ/oFwjvnSjzjQx
JesP+DWcaOGUcf8o69AhE6IoVWKOI2idTS8E69kPRsCv1HP2D7ZdXlEOglWfinmZ2QyBvYYe6A3L
Yt+a2Fl13srZ8tPjFLgovc0bJ0R+nwcMWBl1/VeZD1qisjS08OKMiAW2lOH5DZr3gkuKfNCrlS8C
wSeaE4SlejGGWwnC7SmVzQbkb+8VA6RwPXGu+UFk+u3QAGHahT18gazytcOWv2Y3LCqLLYrufrL2
TZ+TlStLBWqKksK58hN7+KDnaRs1Gcs3qenItmZuih35B7iysOsmIlxzynB4SNaCIrDOl2PX3vZ0
TWftuh50DRqpZwtG/st8wcf8iej/iM2O/ap0UPZpoo/ZfMrkwpTiaCcNmeuCOyesywmSa3d1dfEM
8ozDIzEiL0H1DWDiQb3z47WqNrmI8p7oF7qbgMfT4BwL1tdQyljpSisO42TPwdwXMTubIH84+BMn
hAsuYct5P58M06cdW67pNvufFFt6K9P3jM3Z60LNRW1dPBd/zSRNvv2cw7vrI/ERvusvdziID663
OBOCgPJBVGbFR/lql4Mi7MBvmlGpbmpSwkGdr0NPENVfr2OCBrk5XMFkcrwiR7nuyfbwUHCryAC4
cm94G65w55DWZ7g2y9pmbwQNjk0hjNoQ0L9AATbV9yS+AGESMafIgjcQKdXQmfI+b718OyBgTJh1
Z2jcDD/vnPMOL/Y81GLq+DN7QLIsaSZBsifie5bGCTxMqJMc2Ty9d1LquxYmoPzaSO2S/DlSJ2DO
OEyLu8m3n0GjuuOIZhlnrbY7nGyNz/O4Q/KqDfjJI0rXwq/jltvkAcbbkT8OkMuErAq0RV387gL6
4ycJnyN6Z4HqBn67hhRI4hRdRBScq+YI7mCPZiPL30ryZa400jIJVdRCGVrraU97ad51Nc13NLJx
gqda4VynKzQkKmReLfm88Yt07SAK9xGT9mz9UqDTUaZo/m5k64kqVNAlYtUNOo2Hc8R+As0ooirr
HwXLn9e2YGzH9+yjKua3k93cIbrztixAtOJXs5hSQrDY6BoNFTZFui+2wVMejHdwHXKEC1YVDpcy
eMyEUmP6j071ITSyD08GZUupnPlQRgHbyOB0hb2+7JTouZOcMe9fdciWqq6BPLPVkw9Ef80xoGys
De8LQrjnu07NbcCP2ddyV86BFeh8oYzApjxmZRZ/au1kFYADu+WKUeQQGVWNfh3MJ0IkdwSJuCrs
K0nqCtQVzfRTtHVJt48BG32APcDpwpAqj+pmjZ7IKLbBElsJY9uzlO8203WXGQeQ4kHYTWGPIVqq
4I7qXtdV70o8WRJRqP/qBPO/UDvnwREAw2U7BOChTJDqGPQjvXlTh1ndrGfvYDdBOV2R7JhvmZee
4X5Q6+T14Vkj/wDas7pssE4oKhmqoJSr70Q1Nra4Lb7ulL7H4jgpP03g/rgisG1YIE6D7wC1FIw9
aKMh8Wgf+EXs5hlJx2uAWvqucpt/fUmClvcgMQCrej5jJTOLJlEWTHq6F87J6H6zpoprTrrJhChO
cO7VM1EI1n+iKFBlkpCyAmo+WZ+Z2DN7JLRTGYDg5Maa+9qOSqNxplG25GVPJLOWFgP5+UMDVaej
heF81n0VAx5SqxZkvG7eHBJFMSD1z4qf2FYGFDKjbt4jSIAbPKf87YO+MOeaFjR+Cg6mo5w3CuXQ
hGQStuuJ4JkJCiRa6nFz1niWA3bpLinBOHtFrQ8CfVSp+jtj6jpLaTRtwwxa0gMt/oPlHQC4RmNS
RX71d9dYyriO0CfZYmGjZjIqMvhCKhPu1gGaFbHumBUKWeNhzJG26pWNjGnj9yX6vpnNASh82+6o
mvwk3uYFXXM//WhCYK8cXvpPvJ5TmQFJABP2oVNtjA3aNo/Vhl4WJ6CzYxo8umDlrSI0Pbz7aKna
Sp2t9P7x5lReIKeGAY2VBtw92N9kIUT16WI7Y6DH4TU5uwNo+9g60rZCk0dfDfTAK5dFbm2s+gwK
Ze3nF726ouWMXbXIuAZHkYC3hzdJjceBkgSMWJmeqe1olmcF/mHHkmDiuksc5ApHDVPW3BSARYT1
4UwEhl9uSHvGG0vilcE8Bv5XxQ7ENWPypmMxUzNHUzUHuDRqJWbIehJGPAk6Y2FXP5mqCqO93i9e
qyFWa2mylgQeeOCIMOoIQ/h64nw2vPxf2YIW+DJ9XOGiVFXW3kdkh/Bi37SZsHzUODSWUSUcadEo
fSfln9+A2LRF/maf1J06mjBQKKc1mKlKtFqtMbgEk9goWc0lrWo1thUUf5MUU3NeD4CylrYXNHc4
zU9SrwZP6JE9IYv/nEdMN60xcbFiN6UDYBQmAoNJRm4Kjcvk01otD34vlQtOGua2YXXtO5c8S7r1
PdSqN0POB7coBSkNNcgxA/Py7hOb4TZSsmdTbwpgOcKHfqOtH53B0pmEp/l6OuoMdxkX4HMIpXyW
KI5E/ovo8j6oNjDelHo3aZR5UM6FhHHqZHHj3cfdyVUSwrAaupLl0TW3Lh3r16z7jCAKYwmEZDUE
hgPTqD8hnUS5WNSu0sTGHDy5xxPVTeaz5Bn8RhvBj6qb24+h6cpYUR0hWcMq1Kz2YzvIYDILHdOv
LEmDqqAQTBwo/koXxuR55qk8ELPUTl/UCbraTqRq/JMcZCG0Ywbq9oXNoJEO/8Zcv551X3NN7rrj
uXwEZeMGGn15vhe1m2lUlAUtK2eJH2MyCz/mKkKzd0aKV/jODZgts3ydnw8hn3oq19hjFneBuQu2
N2UG5bQr1sw2rchSHjNQghm0twYCTb1x64NK/EeNC7zwNreB5dmCHs2y3Xyc14f3oTl9dUDQLqB/
KI0GWVAiFFivFIffCvY8qT+XryH/rqr+12X4u7mJPoN6Mwebku2ymU4v5GOLHwpmam0HvI/C79k7
vf/9K0Tu8ZHQXg626qnUbLn4/srJx00aXUpn9CDskFqvZMTn1GS8iUQu/dDVfpLu5M1mhciA2B6l
Pt5cQZqFN182mfnomym1xxdu/Q7GKL9MF1/+0PuInU9VvWGLrLM2+cGdDPZOh9Liw2t9xc2/xJLl
wHTQNYFxAYhN0qlTSBSLyNyCNndTW+MMma3qVth1TUUYD3PNLaniNUZBtkR74JjD25ETqo5BJOdY
k7rbU9G+qgGcV0T1t8QSeneq/gYOWx87jUZjrDaaXb85zODmWMJolI9RUj0FE0hfH/gzuYQTDAtC
SPiM4rNlUEQukj3AJH1YgNlnY6jE05Omy8Km0Qa/OlZMO3IcxU9bHpZcNl+FV46tcvvjJSyGY3sd
+ao0vgfT8CLTSw/fuaHs8aw4HLy0Ki2ruRyfIWpr9n5eLhg7diAHqMfWggYjaXvaqHlTD8WvgJb9
ecC22FD4AgnVmkU/4NSs+hZ2Fxq5sz4HVEN1AlgzUMViRoJ4fvsreYnMovBhBb5bR5wwGU53W03w
BGMLwqbpxed6Hb5T1WrtRccm/omfBEMuJP0afjUZvVGmm3I3MMAPQWgjgrdYdLTdIHvZHFJfRnrn
hopkvE5yDpSy7EIuXrAm2FiNaTJ9lEtFkLUlIBLJ/gkpWAoulpdenv+Ar32KoZDcSy/jBkuo1w0t
K7YqSzpyjp1RuuWJU3nGTxe29NOe9FpdQlspvVqgd7ZguwsJNZNzUeVDtOHthvMUbaGmW7v12kOQ
Z02Q2PX79l/n/s8WjvOPghQtTvqpNSgc8NgSVgPOxt3RkMenArHE7oOhuyEddlRAkZtqB4zA6Yqv
FSM2GqanyxucM/Z2iDCXKIugPYzIunKMenU9tY0ykiEpQIeeKba6wwErcIBW05dJVVq1XQ3kMkrI
yw8apX+ToxdKrYB89BZhEbWlTjjgArBheaAzKWfjNEVig5mWCuK/JkG2+oFmDpCUJ3vk1LduzhaN
Hb4q/qmjQoMX9cmLfGD/R/A40CWBf/JbYoVsNvRu5f8ADiVCMnzAHzUnqnWL1TN2/sqjMVNLacHb
CIzPGYF76acXn+hukWItGcTnvrN/1FrI+CRDsAHCtFqTPKZnCMNdNEuSlczKjoq5XrjP+TMFanuC
mHEUVZonuw47djd8Kfc8+SYspO07NKwe/c5/zi4J8fnBaM8BOPA+2aqUgqMbhZRf9IszIH2/trIU
Ed5roFPdiwDdwSgnqqclmBj1rRCewej8t5rw8GrzD06aEyfsbwvBarzoHRjXwLGIhEq31mUXmzbu
N7pJcM7GArjVNhRsAfnuzlgGKdzbpxFT1uzbQxa/mfmr5l/7gJZi3FdCraYGzrWEed8Zwgym/nps
2Y1Rko52m5K2SHiqwjbNJ+UyZzAR2cZSV9pZE9bUFKORQYKLamNAxWb3FXAIe3uGc6zjX+wNAZPh
KSjEhavCCU0T8ow0YwbctG/AakDXHZg1twnw2ULOgFXrDSnoTQMLBF/FUDr+2vdDkgN9xrH1eptt
m+JF13AkZKfIGbP4SupoYJ5xRdqKod9U/Z2oTrovSBBODiKoNZmZKLuWZNbxzfNxVVrOlIi0eNCj
74e5lyK7x8vxWKYHPG72scdLSfdKf8A47vF8EM5J6RwyAx894X65Qgmlugm2458ctro7TB0Ji3l6
3DSa3tJBz5OhG1c+dtkj7lz4TFYFN9LohoS5zu1BdaPs7/UyuWlDfRpbOFqjCPFqQVeNNw7Nio+n
uWbhYDs2JU92cwNQcAy7gXejusJgxngldBHIzlkFRKXYGYMSF4B7JBm6RUTR/+BkxEvl9Xv/VQ/+
94IdNprb3GxQ87evqcpLVtS4ML5kjrVgx6m3K6/wGTe2/8oqX9RhN6tRiw3UL6/5sRI8ZMZRNx5H
OVvipkWLlAykDo01HFc17v0sKYfKd8wALugfK9+1qWbetoMsDqRNRdWZYBhJJb9XHDKLoVF3HKgV
8NDP0DLdIqdZp8MFj9nKa0xhFK9TklDdWwl/8SqA6n8569M3bf400i2HnU8HtG2bMCyYw4cCrttm
XX56XfLnsFofNvg+Kx7HTJOjMbWzVVaOPAHDiRkP5Z3r0TKziaJlKZLzZIJtVFWUVh2sKigJNk1N
hcQpFXq1l3QI9ATxJwg029v0p/ulsdl3lOoMdTd9pCt9C8DcJ3MnhQeYyyftXWkPnE9FFKTz5ihU
ZlzTN1AaWqVr/NDtURBLThyIdXUwAVuVWhDioDVldEQM0dfRmDjDfHYO0y1VlZ5vDoYJlRulxVBh
+SBrE7FMiADWXLMBfAJzF3d1uH5rtJt/CvptUjxb0LIXbGzJGxNLidOyxGbsuUhQrRul9bSbXWvg
qFcPjmWhHUZD+dez+PJTyoJCKPeXah6cZOhiX+Wf1Sf5ow7upuD89wo+v25yzdqkn1MMFgSqP1eu
it3nV9NZcJJi1rjDbnRyJAbYIKFQPnuhXE8pJum0zdjveNAda+TjqTy5ZUJP/QAPRuyn+hAeixkr
Kg2L6qQTdApGV4xBU3zIM3+Gcr0DxZq5AgQqLGitvAIlxMPEabThEAiHhMAwtea1U9DzVe2cprBx
331hShYTpn0r0VC6EnSPARe/8BLvwboEjoQK9NxSZ0J5mOmeDVV7kZwIqScvPXUipn9A7DONJy4a
fmK3Ff78RvVqBS1UO33Bo3oWbvu/AktbM4D17RqKboE0oSvsp2YV2I/CfRO03ZAtb8cVS/sx4Xmz
oi6mR24AX6Ahq+69691ZHINX+6MrPY3uKfk4Zg3PJXnvGtPia+rMbmJDowewA14jzKpAsM6mxcM7
OdDREO5DbYMG/OFiJRx16tfPf+lA4Zei47sCLGkTJ9XJRhP6Ant5PUHJJK7+1VyCXqgtBtGHAFjk
t4ijJZVmiVO7IqH1RVL2FPoMrFYfi813EFxzx3SGBuo8doeOUAj4bbZXw0U97KJeM0IRqjXseIUW
rYOaUV7E8raTAyoxyvXu64L+4493/opDmNjTKAjV4U7+9ZaLuX6/MVct5vTEq+A7snXd2Xk0uNcx
Jbd/qRAngvhg03OfA6TstqQ3B1io/XkAFSMjU7vxMr4HeWIKdcx6LU2spRiF6DtLSZ5fhkhOj0HI
PlKoF/uqhYv+gHzhzv/H5yMCkONSySnqSrexpiv8KY6YpPoKq39YF31PJQt2uvahRHeMoh+DE+vS
qGy5KgJXcHf0tAMTsTwKQOk4h4M19IkIiMNdxtp9vJe62r9kRf+jHSIHksBUm3FgfZTtpRmT9z9k
Go7cbVpD5r5mEMwVajeYjHVsh3dH+2SuhXoJSyhdkHPWovTDhxmn4hyaSyEPD6KemwCRIxUQtccj
ICxXjIgOwL1CggwX0nX06JEiCbKiUANWUK5xe1NQ872Red0qFgkahuY/lVkmUd8MDmZjR+3wshWw
yHLT5C5PC+GI83fj1WtM8lUt6+e/CQEnVgyu+uigd690leCStSUEQ5Hp1Jv4d9dsYI9+BGNESIrk
xNelAdlDUpUSXZw3PbBa/9I6dfAN7AD0j/YflH7usqsWub+bvRt4xlm2kCvEcxqb6xigP8ycAc2U
wre2r0PAmdzbhWNxPozasQ8ToeiEEx20orVkfiLPzw32JhG/xJRtFXJnDy6gymWV0EiPEN1LMWx5
stsOhTVeTamil3ttkGFwitpmuRwrQrKXd57N3FhsJ22/43XL5bT7GD00YQt+jKofJdxPa2XF+Rqf
VJ5AFo3Q+vdRzIH6ORkCqSfq2cAcdWljGx9Azn+B8CQ3D8dn4kuyeZ+cNCmRVM2v2htVowgN2UgO
9zk3Kcvx9Yvv2zPhL0q2fVVcLZrzTu4KGmZde4sMkg5JM05I9U3Oo+1pSCC0DiotmJOlDuRez6CY
49N4WLAJK/gh4GJmaFT/KQHR2W2K9WKzVd7+j35L11SkQCD0oGqzMuFoS/sPqxTEg99a2sXUr8CL
U2bcLLPBh2QdcWa1JqdhMpGzfBPdrL21+15ulnUv8m56d7KmpBqy9UhLOZEit4JfL9cCPfmqJarf
dp3UWOvw7VZJsF0Ei4fnYF8zMJvl5TDVqU3hxwM9ctiv/kfbuOKMq7AF9gBNi3+dsMqDTcnl6rhG
y+D42CjAwBE0msjPd77JBQZZ9aC0JyjQJgltX4ubOkRLBOFZap16WEN8QLPNkgcv2i3eyuXistjg
Becp7bUw3HYLxbujlqidCxmapw0XCzK9rVdE9tDxk5zyEbGDFBwz0qHzTzz3hIIKadYx6uHkU7o/
ztPrDjPQsX/cM56t061l8EGz6bScDoF2Uszj6INxnD4+bAhMkygevE8Oc/YX2cT1LQx0yeKVAIxc
a/BeCaq3gpkt8UPMI8eHJunC34o35rfzwr7fppA4pm1LaKcZ3XVW5t4Lb6B4NeYrJsiKCBiZVHa8
Widf54VRSDFUfIz1SR8Nx6YLwYlGU9Q6l30LNZ/LFGi1fqccoSkUg5auKwjsJVVxd1bLcK74VSie
VCQ2P1yhHS7kyP8Gqp6qDhYcoAnzOLqritpyhjXwtOA97cqCm/TsypP8O0xnZMMdZijZBx9TbI4r
Tw517LkFha1V4XcOq/qzRQraQuWY+2GGZ2Khqbb2++vBTewSAt1cifi8Wq9DBnl1wPpENOZHMiM8
T1Ez8j4IC7a2iCfghdEkg0LGOLiA+4CEMzmlVd4F9+gXC8mxRgkdbZ9gyy9kUIHfwj2yZxeDSHjX
cNLTzlertc95LakhrU0lSPPRlGH1/zej+Juu/PbalzXQUqcUvtSX/v4oKxgkG4hEpvYg+xGwj7jL
n0wkynb7FBUV69MtdV4pHBea5X+TDfK7xG9+XLn++7WklMp00hiqXfV2tJDR7Z82fJojEyMtvlHB
N30F2eIp0XDav0QAgOUKZuk8sQMgz3CMWhVYrhMeeDECIkTp/oaAV9TqLKb6tGhytoofyACj/rGq
fDm4QEY8AfmfeDCXoH1pzou4Jp/rC2nBwJktrEhUg1p/2+xtKcufyqpWbWRmXYT8N4d48QX9Oxva
x7SrfFfAL/9MH1WsrzOY2qad1G7wH+ygc3a0gw7EnEE3NM5B378fL5Z16pvzBvVsRLDF5w3ptWLI
rPLoWzK6nCsqqowU0tUwJexJGtrBgH7qMF5PjNlIDT6RdB6UBnpa4Y/hSgHckqMRyIawI6O2WrAa
aA6bZnnn6i6FTHnf7eTsjzxUKOtj/ssv8eF2oG8o8aL7JenXmJ0QGvA4ASmDTGGtCgu4nfw+h/L7
m/S2ZnoLZWIq9qKkry+DSPY7UjgsHaVfbafAxUWMpYnvvEX6dbrjEdzi2to/6E9SwKwZbojPEkXW
qIQxQCoJ8FOZcmaUFHkLMzhKtM0dnMhE5vmUU0G+pBc5886ubF1C5d2+joaUHSwPnSYLC6//FnWn
ZZqzJpu8QSVZgIwly7D6vWxjFAu9QdZ78vnxSbayDhWs5dR6FW32FuIoQjTEz8W+WkFSOzf0hVpd
Io9Uci/2IXLM91LSZFC8oSOM2qN9yugbjC4bDcg1gJp5VMIx6CZH0vtVVnXRw5gYB3O5x0thloxX
nMaf24n8ZpSdj4RNWS26gOeQKLvXTtkrhrnXKTo4FUwjdWarL3thV+nglW8kivnYy6NJ5Pz11MU4
lsozRVeY+u6YzLQXr8kQIq3J7fJqrACBXEA1Iv4bZ/TFUhD/eKR9SEQME8+kzhn0woSos8rOJOSZ
JFYZVaI5OCJxpy84SH94H/pNbSd5F4eIwW7yixt6b3zcxfA0nIksDLI1VW0CGUuB6PjFEC4eqCBP
/YpDLR8IrVPHo7cqK9vVkaDRr5YzZkvVTkqt/3iOgqhvpoykJ27ZByUk/RwhgvE40dvTAqR7y9Oc
8Sf6/K0+7Qtk4YNJW+CPeU5VrzVsb7Ej3Qvx9ons6N+RYaaEFmj4pZCwt+2MitUGKIDid4wUq5+g
KifdhzbTKkIZoz4WvWHwnJl5G450nHU6SnWvIFoF7lFJ84iY+X04YIfZ8UbW6TDVe+zri4ivMHXA
xaxhy6OKVNuay/GlDzZAylQWdgzwrBEEzd5xWvavJ0fShhlYDtr2Z0nliqTecpqmhv903esch6VL
/cppEm/sDTe4urr9JvyI8uti5e5d4RQWLw/JuGFAAP3X9yNSnCiHZXqU/uxoOk5aeyzmJUO/4vq1
SNvBA/jO+iskoowYvfq4KL51/JVy3hIXS35nsx1TOMZ/Phu+IjjaXdEZCWMC4b6zLFZ/ZqYQ12TR
5WrbqBZNs8ClSm+1chZNDD9+Jn9MbqYy91llJyEGi5hUd9ZthNAmKunc+5pv7JbGr87AsgGYEXLN
Hle3thSalXCpsD9W0YgFt8o9qr0b2BUymJqyEjMdlzCFiW3f+bhCtQ0J1qE/VfV33RNXMSk93mrH
ZIalXEtyBu53NJQGoFEpkJbMqznRvp5eL09e9X2xgya7Qs6wpgtNIUL6ZinqAwziDCcu91K6olci
Jyf2w7G+P3+TFdh38tIu/era90Iw16jyjS6HaNHVmwX5IyRzmx6om6dH3IMWdymwrLA6+aAhwXKL
8iMm66R6o6ydhKBpMWFQnwFuIuJ3IwaVMWmZxRsavdTyzdZd8j33f/MGt8xVMQakudoSsUdsdvm1
Pqz4LipD8zptLSiG8Fdf/Ht7TAzjZEbpGnXJlmqE4A5RHgeYCKP9409ijFQW9gj4rj3YRxmnmJHS
//x6iFpi+jgOLzf12CZIQbMNta+nQkgeOwyvpdhCLA3xIYLgQ1LCkyVQ56RZk5N/3zI3kAENRhsz
8PusDQyycOruXiEI/QMAaKNtB1aYBxUh+z/gQAP6StojeKo9rgi+WxhvCTpE3CNysc09gayPN25p
7sfcBUcXIrTSusC4Th2HREe9tCvRxLDCNdemmoA0Y1AduS+9wMCrSGpRhLzVOGiy0IKF0/KpIq6I
NxDCEFeZysScePTjnUM2jdrQJPd1hOC/6Tuz35TBTOCWKS6lOoYVzjBwz7FdsazvJvDvSwZzq7tR
MEimjANXwX/N//FBayoYKLZeW4dspYfWS4EJZMCGuv97NuJuDrc6+qJJ0t9b2tgD4K5nshac1XdI
BfeS/HvOmmw2uf34ZCe8NnzdrBNeXMAW2I0NJJVVAOiz8RfW+7e6edC7/hYEHg1I6B1/UPi0VKt4
wGKTMqOuAXluRjNCfXMphcwnAmBzsarvh+dYas418emCuctMkK449KzjtgORJcZ8HcQ4RITG88C1
weXFfiLZnDrt7RwSRTnJosuhdoyzllnqLKdzQ8j7pIL2CLg9V4btKQlxfpUKmhIp3tNnaYs/skyM
qBM1ffxlVVuurl7ywdb+33P2RGG1xkEpqM/yz7uje83pX9/+/JStt2Kkd53wTFvwf4hX/1UwNXqq
DEUFivGpq7VPcNi7zSe40Vuvh9PcYLi4Xv0Tn0mz3AuFLRj5PCRw8bX0ZJ2fOZQ6PQtHYxNuo3/q
1XqRx7V57S11M/GvTXpKGBpkWoDgiij4smPI11JykDTMpjh85PZZlBvuMM5cK1+JZPCGlIAtdHtF
n8WvoHPqeeCadhOm3z+MOVALMmu7IEe5RJjZn5YdsIMfphkTFFDPBG3VK+0MoPZYeUVAMofdl3h/
ICVm1HDiGIqroeX+p4K2XwAlZek9sFZiCnIcyyYPAFgj7pIfmNaoFLt39b2EWApThp6M2wkKTBkV
K6n9t6ihlFpInPMO0wTdW4Q7OMfZaqAjv8EO5anZrzLW5fJt90RvbQZ6DmoAx7CbHH3k9ucpIHOD
y/r2WSkRiN7/1UoEZ9aGSjLW7axnzkTbXZzl+YUdeRg8FCY/A4C6iiVv37Ix/kiBNm4T/YBVoVDr
fIgSX42wyxSfjPjbPX1OWzjExb8KtzMqyHQr+/rGyLcG8hnfqcIQ4XT0Ax/PsBrjGqR7spmLd1Hh
JIpm3fVNcSNOW64/ooSpEZ5vjVcAhFcHAvWmhcGArpZ+ac7XfB0QgbKA6T5B397NJkkcUjGxDe/w
7l1uGKGcMV3XuMphRdY/wUkF5XesfxwiddQua18NRSLgGCT2ZIPuCYviGwPtmRzftvrK2qhflJRp
HBj7Zi7YGSXC9m0vfDSKf+3s7WxFGTn8+P5FWjWHz2ojMlcqRMkRcVTcNT85HArYk1KX0OHILGcD
KqjD3t+Y+uNPHcSSunhviAG8/GL21M0uBePSGFfYQahCfQ3AKr4IT7slLO1RGyXR+6QyphiExZL9
6To1X374kyvGRGPSsCT4Tn822KboVAwYDc3wVc3rP8RDts7MjQ9EqGcD6XbUgj2q7ndI83SX6igL
v7/SFmfPY+phuFoYG4IuIc7q/o+Id7g6iuAvnzgcV+6dhNiRJsxxQNZe5DT/xb0ZMlS9EynuWkK8
eyjPfuACT/uw8IueXefu7A0LscxoTdWbt0gz0GFx1HxSZDBS7QoRH75luyFJwApIEpoR8Zft2GK8
ZT5XvA556K6rLq+SnPFwWu1WswAoJihxIb5bIi9HFz7iD6FofbYomL6Xd9JRBk3Ps1bWBxPUyk7j
nHNYN3EQsPVSt47aYQRS3R4ufHyScYgGM5zOut0yxDk4PI6WD9qsPA8mC+zummtQ5sQQ8/6QeuCr
CDTF2V8yArWRveXXKdSzVluXWYvBOmfrgzgnFypznb1i7SXMB/nuU8+HytKaWMxmWcMJLbOnCZe/
go9kd/FZ/w9IngkGcHlgd02YqC0fZdbdZ7PsduUE3Dsc/dQLWYFEPgH8jhcdpnNV75l9k+bQWHXw
sFzrMR+T4SPQC1eCiMjXZPdpmadS8/tYz9+j6D5Dlolz38Ijq5Nb7exR3mSVUF8sGfIYweSAaxw5
vJIgMS9upJNrl3ztferZwQKGr/qVbpQvRjnu7142M5xYkTyEVsgyVi23E2HGS/jxFntmWpM7vZ/k
m7qzqn1w+TgYxcjJRvrOEzasueJAqZV6zcyYVKZLu5qjQyaBU1+Sx/R9GRl9MSZwv/rUW8VZkG2d
FfBYiLVQnrv8T+XvDc5IJJr3gL4ogYAnup+EUNEiGfjDMSqHEGwrNr6Rf7W6Ym8nqAMmeo1XBdWi
e3xJQZwzAWhwzMjClAA8uMeVI2ArPnrPKFvccu5dsFi9PYel5JId/GEmX9zcOkChy/oLnxh4GjZB
CkeJQNTN2zd1iuJcmULAtA2SEs4nYFnoVkcCropChBYRC9F3Ku4Dqn3zhaT+iGBb4WQhZard9R8X
1FjvaYW/rnuJu9GhpiYhwbLTYrGCZ+Md0CmkQASs5k2H50JJOwp9m1T0BSohB4fcldJVU0ko9jTs
ox32NrSnD+/3lUZnzLj1UGLVkvk8j6qcSsmMY46cv+PIxEL5xyyAW24UpA+G3T71F4er5HA4Ph3K
He6LlF6DVISAgEpPkrJxpemEZGPiRRu/i2AYFyxRjfjIOP1HN75yJa0YCBgpDNlyjyfCblt2kIDZ
pgRRPduc9Li/2b2eIP5zpLqpQaIrEOT/EobPAPdZu3lJidVqldEczQoyKnLSVkVB+e+2DUzZ8r61
U2owEcdkLNGmR6F7V0+YWNL+0961114H+Rfufezyo3Tuf3GS8bCxpxHOP9q+08VKtfphJQrwjGBr
s9c3vFBvqYZ2lCIDBEhIJkaqKCmmchcPNh5ruTlVlLA8aIviSBUYq5P6CUjtxzv9uCDtcmUitvFR
UNwcpQzVAMCgTYo0eZZCGJ0M8CMbexOQrKdLFp5Hnq+a6mVV8KZoD7y1ZQh8IB+02yc3DHF9ga1z
xLzwNxB5/MN/er9z0+DbkY1i4hqmm3qgMRiVVFIHmyUfzHEEKc6gq3oqJ+vZaF6FhnhQ3veRZvBm
OyGMruegZH1MN4rQFpxB7kERHRrku5qQEacxu9mbhmXhxC52NuACBCAvJMH+uYAUK3RlPauNziFq
KE06psWjMN72SJHVXyqN+zKeykJSUmXyxr0QgpdkYvMNj1LBFsrkavCxOayf8VNyNyS+aojmRvBQ
N882kOosEpoKQ+VAS6QVcuG1/jQnuL9TZ4ha3ds3uckGPUFjcafBvazkzcUOK7QYycovFcp1hQq3
DZQs+BP5BggTT6wkIsaOoijJTgngHIi4Umo5Qi15bmCmPdFt6Ulu2LpCCA/r5/iBFGVO/Xp0cu+z
0ZZTu+2E4FiwDZA/RCbC7j5loan+NLgrzuJzvo9qbIeSHwKFBZAtKO/TQsrsoSjEyqSLj0c6zc0I
NcS2lWASwmGbIcw7G7a00HrzxvsMRN1WlHOKMggT4BlSbxkUSIDVV5EjSucqvAt0isMLmZ9VwIo8
DbYvSOX1PYRXIu15Ux8SsaEYbRIBCD58i9C21176u2ySk2gUfVvg931YNFSCqe8rf0XHUAod9X4l
Is2lVsMCf3BEcZPxPJdbiU/dKg43jQeAXXSJLZBudLOV6+hgC16Srx2AFs3MYqfu70G0EYa7lTcu
Pwsx+j4UiYPfPWygoLBWNksgMCHDeTbgWsSugXhnixSDjoas651k57JGLNS7smiRWYIp7WEPUKwp
UvUKIbep0QZ3EhSlnV4QFyJxh/b1nFMHyuj66VsjrotV+LuwyaraBT+LivIHHIxVDhoVLs8kFTPn
axRq5dwAI8PdHLEANqQ3Z8Tm5W8h3kUZLHSC2LV5egYFyEtY82sPCW7WfHhDwMIZmRun5dFxiaeo
TIslVRp1GINZl7SyEW8UHdp4kHscwx+QjivcAz6L6WecmGRDq6Zl3CqvYYwdSfgSHKkHoeVWz/UH
uvo1wZEeT++so89eLg2UcwzVf2s68UgwhsCh0NkHocmmEHZUsW8mFypjXNIJOtcmVtDX8SolXfI7
N+KiqcQAhX8xtgP4tifYmPvhQfDEvArUDgV3yyTpo0IcokaoCChduM13q8tDpPJuwNER4fwWKaR+
VaHIY5g/LV6vC2LjUkxiw9oVBJvjLQcM2y4gK6BFEex769/XHobLZR//5CasK4g2JdchFc5a7l8h
ahVWRhnDJBh2MMbrBT5TCamWDF7TK4W1+MmLkWx9AcPfMnmTNsRHqEbE2tAyo5GGzzGNz5hAtpui
8NjEJzhdITgfMuVKd8UXqk9z5AJ5WMGMNVIPc1rrJT+i7FVMirHTcCp8subgfx/VrKR/p7Uw+TOs
6PrT5i3FJvISuZz3YHb+yRbxRAaenS3SkYkZ7X5v2POvRGhRQ+pn4SV+ukha5S2DOMm0C3SMHSR9
wXsedUHBUS92YCm/ep26iQaEL81zhKk5gKoSeImDRReiC0iqYkeQC0LC2ualragPrSF1ButwzUjJ
wKYuTBEY3qtn5S3gn0PhH8I1K4+KDtoSkYCfU01J5vucerOa09Mv3zVEgnkiWIeH+bEcrLO0osUy
7awZ5OotzudnAk9I2SjQWnzUTcLnKmwxHn8l5NA+v728NqA8c3MdKwxokBoVH98td+tyl3z0q42A
S8g2Q/mV0sACOANI4gazO58dk2Le8/tynxm+AmDFubK5i/Mz5KJPGbSG4TlO44PHbaSHVU/AMXWk
wgTPcOvoJo+bgua3TWXcFbbiqwd2bj8YMvCTQ1zF7TN9QxJfAolp9ecXfQ/KLqu3LqV6pYOq0B22
1griJIPvX/f5BAGaOMgQXMivHQI10sCvymvVjI2DKUV7h1W80qBtLdOgjGMy1/+YnGDWx8fktO/Z
VX37Jc5kCbjRmJRZ/cf7tlf3feckyWTeB9qKS55kP9qWw8BzzfISXz3caoR+EIjgXORwgPYEJoPL
VeBhCTbMWxI6F1wdOZwQwaT9ivJ16YbHG9OH/CRHnmCNxrqRQyHpHmm29Mmiy/yMHyYf3WKqHc7j
OyQowUn7aaqBNuZcYRoGO6JWGVg2zAPA0wfkuU7ImDjLGyfM3pIIU5YAbmJcZ1R4+hC4od0BdeNt
249pm+8qjCu+Erw60vG9KlC58pH8kpvOeEEW2OVOIJnWBT+ef06hPSN6wZiwQCJAwcPWnWPU0OCm
1Sdds69bJDH6/U89Xa8oGEuSP2XenqCHYH3LZKFc1cSgJ/e5qjonpNOR5NLpAdWQgRXQJha3FsYq
A6+QRbg8HFk8408i3xa8AO9TTkUS7NGWisgeUj6Db6F8GDHHELXfXZPAYGMeNtzDI/FTKKlrTdMN
T92buqjVqEEpABhRozIaYhG7gQXRuPIw4aCWzDn+2JvEmvbPsEwcGK2OYq8U04Uz6KVRUpUU3OMu
WpEEbS6niGVy+Vg4FvlmqqaDDTDbjrCy5041ze09YOTwS3M81lfHlbah23iUe6NUsytm7xMtoiI8
+8LJ7s6zamFCW7Hqi2kUP474lBh3NIZEi17ufvCqYTdW6W4LOeIFJhDg7Y7MJOWvb9FQoF1/E0T/
Q5qYvLpMNXvLjSWIsHzz2We/rb3x4eHWHPB8DiF3A4YiyjeBS25wVLePYKxi8RwjIxnet7fZX04M
vsDL1gv9fu/HLadi6+mzaPAHtMc128MxmwBjpqZPh1iQg8yWyIUn0ruf/FVXofY8Tbq3oGlrIXVh
ppkIhueufU0tEAnjv7BPY4wHRVkSVekDahRuHuTrLqF47UX1LbfaWGlVCcCiS5zHgxKiCPNUcqG2
r6133L8LG53xSEbkWVO8ffBHA0KYzJyiKCH6cAokdTv0niV3xXLzYQYXmMaFOrSgmHosYsucom9J
ZQi8WSv+HfUMUqhv4Kn7E1N+pLi7sLsxlsmNPona6WVEtAdCpwqNr0WsdCPQx0NNEkzodz7ifzz6
xvLClxRiirVlk+SNe3OUH7qye3YockS/IKkw/x65ULGDsdbmNIT+lZG9zxdsuZLKI12bNS5S77Hj
4UGVueIBmwzUJ3ea7zd39+stH1quuGtCnoyozrUDt5os32gNuNOIizoX4QiWxxAh6BO8QJ0DMg0g
y7uiHNYc338uZvjc9lkShoMPA5d+xAUyqdGvTsSwogADWJpdvuVeZ+beJh4q+nc4GpKH0rvdoeJs
UGtl5t8sNjFE/TCyL9O4XiLbOBAVab/vI7zaZ8uOGrj4dFve4HcHmo5k7JbkSrQrqQ1+YdfWipXY
gv4foU3pqJ/mGXAIbHPLtmHh+3Iib8CHZ61zbbnAOoAKG0U8rT4WRuaBPWkZOPOtLF/gB07/cYoR
cjN396ZDistltp/2XuxFTz7SewgPERZ+w6TzWRGRMFrLDeZzLWCYk9CqFGKQC+fSgGvXOy3RZLWf
oYtqTtzjLiaBDb+SmjjZDcgQBSYStH/rNPTNms26kOlJAPkwqIsGFVrgmOR0vON+il5eR6KnW0nw
RBWA1+K6qTPcSXKsbmLAERKjGHNKkd3XL7RGyWBCmG0p8wJ7CcIhr1dPebKn6Z1waIj16UDBt1er
sWbLk2SZmvnN05tk3b9WV6sLd1eNUqMUmzycGEZhB8woyiNKjs7LQoiOZIkIMpcEaSFZl1AzlavQ
AXMmF6UXzz+Vd0YpdjPBuo7SaEB2r6q4QqGi423FrkU1sCJkVKW9a0RVY3T1XhqbNF97IPS60o9j
qRfqvHA39IYQDZTEuWm8W8CfcsmvU/E0BQH4GMKHvRmV0dwhi5MAGbXWSESf4geTE2+U5yQb7BLJ
BfEnaKULZrkuraOpjozbIAhUt99aMsIbp6K9ozoomCTVtdgvf0H1LCOhn65rzkzw7Atj0NmZaumJ
SBHs5MaGp3ZaZDhdVuxxz2o6MJtg7K9d+PGsek9q2k4oS5Q8yJ08UkIMSHyPfZ9rbjIVrriY+Euq
KRhh7RMkcLRBm3/0weWpx8YTvEUaVpSAZiRQsVxtw8sFYeIzfoeZuYmxanypnfLm05Fu6/+V2bWf
JVjBvP5R8c4r8VQy8Qi58TIoH53AIz01IxekDLy3Jw773MRREn2AlyZ0ZMjQuo3Qmg2nw8HmwqrP
46bFshWNengWLXjFhAw5MKmWw7ImACz87sHsqi7MVK0wgBWDiqjTu3fkQjZUC3EUYxltiChJFD1X
pAJFc0l8ueMpmSaiyWuU8fTjpplHlbzMMYX7SpQG3fZTXyPyYpdleaLEWRU0msoJoQouRUQlaxpY
U0dRxjNcHzq1d2H4KrBYD1iRCzRT9D3i3+/9NdzBVEqRKrTbjAmnf4tL/hqFuYBFdnhq47KOC2F9
MzDR2Ox+igs0cCCZR9Jg8eSO0GYpvAKnn16F+oRveS3whx+lzfouyIfMwke97FxZdr0iIu6H5Jlc
daC7MeE39Z+OyZ/s+h9+sX/u/yhAmJP02G2qsGHA5rKGIG4dPoNj7peNoEWR94tanrWOegLMGmNv
EWhaFz9/ailG/7jR1+nKfiF6oS3fSd355so96lxGvtxzYq1sZksVlQ4TraBmXfy2S7iVLEheMPKP
CXsDfma/dZdkH4LVdGWY/p+pVCppbYBa9PY5bXJIrtqzp/r34PFf67jF5ydT7kIEyQZ6eUQ80S0N
tXPTskW+QN5e7rZnCabUe/TtRk99+dtdkgXdwfbrhkIR3wihPK5REff6LfBTf347C/ScewDT4LDk
xzrhpUcChwpdC2KWACGEztYye6wAIzMH5/QOmd9K1mx+bejEulNtIf7xvC/jAKnTJ5fjoEf69vIc
70Ybl8jognsZcX+uoz5oHxj1cGxA9VdPT9E99Q7Ha+30NBgQeW801n/nEwdiGTmRpANnBjQwkyS4
0Z19mQjPgnmn1HgChSms84KYlvuFjsLi0mb+nFlIu58rHSfygpUI5mfHYS6Da7fhtSMyDi9u165B
PVxY9ZWtBZGn4dd7gET2Lx11SB/M7IyrZ6/z4ND8NZ1TE4nF40kAqkkfE3lh2XJDrVhlpnlUUWXk
CXCpWMEMo/LGkehiHcEjEspNYEnWuZ0AMECZLUDL+zHqimiRQDO3dE7kc94bHmuE7u5jAq1x8r6O
YHldzj/r23tHzaUqSd9XZSscmlYB5nEG4qkiQ5lcTcSy/fKQ0P0S8SgA70VtahC8RpO0RmHgiwhW
OzihziVWtKHk1+cm6zitcVw4jfGMZsPF7vSXE8lXZsbgUZOM9pNkW3kI5OcKHVl5gfJnq9B39dyM
8Gl5VWavZcPp7AwJlwKcIqWoGQgdIJCYll5NjRM00aSnt9E8sc3+dyFqgvVUmRY2ed67OKuk7vTy
YQVPQ0tIwf5ZvJNjp0nbnTtNAMLDY0Wto1LbxuGRQ25uQRbwKsDPqDncYmEZu27Bmns8yycIV/wD
4o1Cz9JC6DxtOhJbW3cx4rhNa8huftFsshprZflNTHYD97NOyMf4GdpNH4iIJcvyzJfsM5qVKz6E
iRjePviQapCt62zjrnaKEw5DPw0YiE8sxxAhsHMwXW1ZyXvbWSlPpMO6IG8OzQCDUyNjyNzCrGvJ
hJYUsxPrwHLdiuPVOp+is1UVGYOW6AIxXDUAdvrn3Ph9270ahuAUktfvj0wtLNcxhYJXaotof0gY
DQA1lYRUMkJIX/R2wB0JK8snhJ61VIvTFdJaqpx+Bui0K62awWv1LVr5TTTDqf9nso+XTCxOlCSz
MzNZ0c84HfNNSlwHhVNxlMuMxrdq0zt/mlVuajEqK/BwLOAjRv33qFfvrAgrbAdT5veMn37rFF1H
2xxOPmnBYrWaHu3+GZE50pNWNkLKWwRCAhmApOIRbhkqcauC0Kd9RZU4v6vSdKomyIbaFXwldOmc
1QNoixDKUPqsAvN0uan69rHfCh2iRk59GyZdZDIn4GMZ2dce+Fnct35BL7PhGvlTnJiWYSsczd6h
DrkvTjqsfzqF9+mVn5tGrlt2q7Jx+ZudLxsrBLHFJJLcy7QMm45lolnD5SQrIiAnGauIbdECQ21d
JPARzmihwHDQ8uuPs7bMrxTKTTauWLVuYkSDTb9711PVi4ygfeFVw8I1rYIuAnjif1HvzTSKhqMO
mVSu+EsblyuQJFcr+nXoFelSfcWzWDu7gd1FPpkJrUYZPoUbfoWpixMnPVZEd8MUkCl5CRKGal/0
1R2X/dXhtJ3jSiUdkNF0qCRWhgESOVtqQBcXnaJZu2fJqZDnJ7queSvWqbnyHssgSeeO72S8/I3a
HDFf6Y5nUMVs0ihGfXA+MrQxi5u1ez3oBr8HsAdGAsa95ZIAjdCZ9haJZkL0wC8TBFTBzpbzQ2vb
uVIK5HxmPqD6VH45o/6x9WAmvAiGez0IsYHcksu2eK9vNJCGl1HSMYNm9q0nigCXgIX0jA2BUb7C
1Jyetxnjgr+FLBhmOHT7sc9TI8TrzNvNBi572ap7vC5Zv+gdtJ0Yrl14QKo5+EJgxdkgad4c6UgS
OM63wv6uFtpYMGjShIn385xg+yYK+4ctoXs6q47SKqe5JSZJlA67FD6X39K9JpPDiwc1LPQ+hDUs
j12EEa2R6e3GpAMUXdLD1kMmOwiK0fc6doRuGlS6t94ToeCsx1UhV0VY+D46iVL1i8Hyi0gOLAPt
DRXSb7p5m+1PbMJRUaHkTsVQm1E3EchfvtURd2FXRUL3FRtyZycNAv6u8lzMuQeEtruYAE3eTNAi
Ed5cDVQFIlD+sZxcHHpGGyq0QlJoA6koxiWQMrmDxniC/mzXLn4VXOr/nzoyn3I+syZKpkE2mWsv
NHJvvPJ6UBhOs3BSN1QJipbh1YIcKADgDMOAHyjozlDSMNUjBlzTcj6a2LK8n4sALAipQhAFDW3p
lBAyTy8FOJ0JBs9Dqzf6HfJfsa7/Y8UR1mSCw2KL45CdO2tHU48aUTS9xReafazbDMtqV6Vsv6Sw
+1utOXe5jy4vrJUqCo8Soz1INTNUP9r3aQCOcCdwoyh/s8zaL/cm57I4B0r+yEq+P53XJxbU3jnj
zGG1MrvpvbEbLCRJPnSX9pgkOsvWOE4a5C1l+L282AHCyZ/G63z7YlpCvEuv3AIdlMCwDe76DYpQ
l1ajnX3y/qPQph1OFG8245a4iElgoJEROfc514j3VIhr9tgNUer6anSvaz1zlJKsNQSaQbD5CS93
TNjB0E/0qnppJy1OQCXjzQ1kp+txkC4PZRmpgINla1KiJUKMNr1FjWKsiQ8Rl82jPLepYGZpfHEJ
y+fvNLZFNIfhK9sBJSTgidvxDRBZMTiiVus3xBnx95ts8uacUHmzL4C8BWVcMyokqN2KxO7rEGEP
4s+6acwPSzMIWZODcqnUioUijwFXHmgQZlvGiXu7s4TAVrygJAO/c36uSEtxTdSLsQYRrjOe0tdv
U+lb6tTW6paPfvflD7ki9KkGTBxpa6e7OGzOt/OfUR3c5xyZgbLsMDkswzC8WgK/4MNR3d+oBSX5
xEgnvJOkf/8Rmpp1G0cZzgMWsTywilEdAe5Su7ugQ7rEdxeN4lsoiE0d5Yi4MHqWzC/eiKeOMJdn
5JeWkNdljDQgAM6eayH9cGKpuyV4+Wq/lpkPRuYaQJ2sHCmbkc2K5RWxg5Gv1d2KrZRM1nUC/4Y2
jRXzIUirZ+mlEEX4rpngXt82qTNTNl56ApEjpBBqHDx26YthEc1jR0LONS0Qvpx530WjRV3gE2i1
AFGMMGBdb0i9yb+uQ2mrRgurOPIdrzf0O7cyIHWpcQFV/J2aG+POPOu5uhDZSrgzBMWV0ZBk5toL
hIN0LSJgV6scgw7wFQTSP13NZWOd2BZ1gBDQGeoNeLrUhdSI2B5Y2eg7qB2haKs4B4/v4OW9y1D8
RhxqIkr4QMF4ImKqRjOqVIiaZMRPsLchnax8lyoRDhUptNtBgINkL8Pksix7SKdDQIe2Suk7GWVU
+7ejoRYPByAkjltknbmDSC1ytTf91lVMX4YIoWXFlYhOxJ2cT3nE9J+68hs+dddar44yLUkS8eSy
TRjuI6Xci2CtOx9QKYGhwdPbTXuPbQ9CsTSSSU1MFxhh3Ho/H6fjIE7FpnHXlGtsK6p9jNVo8hah
mkzeBbIRKRA6x5lQk2+JgARfbjGTa597LyM5O0Iz93EiAX+VNK03j5tw4EjmNTQ2JhteEfOCyT/K
BWbSusiIUFL/w/3Ho1AS1OUue/TtYwXpu3g/q60Jojb7TFoMOxzYWICmfWA42SmoSxhEuro8QiUk
4Gm111QJqrUyf2hp6vgyCBLatF0gEzqHBM/9DCbtMkuB1Mop8remFnP9wEkace1RneRcPU5sm40b
fUrcDzQBLPJdFpqUHoCiC9Ev+CXW+qabysjrro3/BVc40xO5tIZIDHDRpipK86B2uiNHRzG418KW
TK3HNfmRsudqJ1ofunklDcPcL3f8kOWrHYK1aP1in/cvNvfJBkhYfsRl1v8rLI+YZxvYPzbh29Cu
rhW1hhFPkWZiRMt46EaN7P61LZou4GIfHOj0/9GwlRdiQK1w5VTko+FldnmWBq33OYs0TDTU1rcO
/OrBKvuHe0eQfoIpmoF2jxfGWCh1mBIa0OlNVD3xRi7YFCF2T8iyp5gK3KNoDJzTKq2TPxdUwz9u
SybOOO4NK561Xo3W7GnntQDI/ux7weGd5+mCnF5aaKRWbt4ZRt95zElbz+bio3ddnn9i6mq2uVvz
Wwio51A6ZMXzXFsO7WrM/iYLDz7OlLVEuf9okUoQQvJ+fRI6K6wIR7th4gCnOGzws+ngXqVtgt5E
xGNa7zvZUSgNEh6r0VUz8dWe2ts3jAwnzdzPQlKgY7yg/YId5rsPYnxp982mBYoNt2EomNpUPsD9
pvIpms7cjor2awN4tXJ1JVVmFBxshFR+HA+ppQFWyFF03ftDeTNVQtLclCdBqnD71ki92UDKewno
jgDHzRqVwLrBW7b1GUq7sUDIjpXV6l1RVYjEUF/bfoHclOWDBovNY8ZJKUijt8ZMuWsvj+F9mXTt
eSM1HjgalNAjwnNNHjHU4uDhQn7HwD2012rHP/4JuSnhEatRLfx7VjGXPsdNyNF096RTIpWkU9o7
g2X9STnBp6gwGbLc9ucg8aC7Fs5W9twwBsUP7CDBpMEToqUelcIh6qZNsFe/N3qgKQVUgdy83KZD
VGFNFyc6LaZOP6L4zWMKL8c0Ok+G7pGsj+2VJEZBy03Vid1GozDtwKlorHCcHrYa2n6wNOm1FRYm
oiYfQtz5CR8ImaBi5tvHJ8trjHCBGbzqhsaBI2U0/TVo+0bdidNRfcrZ5pGTWH/T5b9vnFUF/LZG
q3J9J7T+3XM7Q0wBa2IJv8zTW557OaHoRNxdwXWm0V94uNW4PP5mkvWmK33CsZq9Ipdjuw37KWUL
EN0iuM+lFfWfpZ9YRte0xCoFQWcwjZvtnMKSW7MHGPtiv5F2WKaHqyE+GxTnsrEn9s6pru/swBlI
A/gE2dGEPq4LNxVCxm9Enj3/EEMbCh2qmorD4WIYwWYQ2VEFZg6ZfnvUjy61WGNODeHBwqkYK/MI
7ba4WeLLFcr9AB4061HpeRx/FLsFx3RU34r4nfNLcGWXICYpRQFd9NpENLKbG+UWMhoChDAMcb3f
0l5MvSISIlJMWn2KtwOsIHb+eTV7qX9C6jh5Oy6RLYUYSLSrGZYLSEELKDCnXSVLa6lScCmOp06Y
TSoKoi1HHLyR6/kOvola77f3dB+eAcnq3nuZxU2XFzQFXA69uk464BIxQHisuV+o+bdmdOxd64Cw
NephmGg5n59s0fP6e1JVi4ppM4lFnGztB/O60JiTeBmG/dabnY4+fJDtTReZuQXV+VtD/SwbTN5W
Y9wKiQpAHRSTmisgMHmFHyBifgJvjhgDClj2wVbq/l1GvUBZN7tgLC6sYupUDMj3Hmor/ml2QUnM
eJoCUa87bDD5FwVYIccgnsUYCL3W6SczgEH4IffcO1HrIZ9GuUuYJsGJEyc24EqgElNPS2COF3bh
Aa6CLZTAPFitf6Sz+NEm5UOxJb5quIiXwZ6eJ+D7P+6+0syl5HRVsBBWWktvE8WSU8TEI0i0omPv
FMV+OuXUKQDEztE6FAjvycat4eUn2IUbX1msdT0qS6fYH3POiItyBlamYaK3Etr07yIop/XgpXDU
n7awbQxpAIFrXcemhNoYvJvD+eiB1Jcb4dMWGJHBz4V4lSZFrG6wUtRhUBIH9aw6e4vCMeJbdQeT
+pmY0uuABDGeNgiwExvjHXUPkKUsJycsGhPOlucZBzgP2dPN7dqgjk1bWXMLDsgjZWyMvfvu1ktw
e7WXtRFdupQ1BWWsV1SuP4UZdNINS8JUGkA6D0JJ2Ko/OXPjRwI0+Ju1Kxvnoe2RaIc9jhnWci81
GX3QHTFjgmQ5a3CuGLL9m4FSZBMh1MlW3Tgd4cnhbI1gZ2B6vvWpMNJuZSY0OqOR551ZKHxMUxfp
IcIR4hLMqCybgC2Ti8t02CkVTf7+B4tWIeTO1oMnd5R+ZDsuExvtRds+glCVJ9tSH8MeuEl1t1Yj
7jxNFbidMC9uECrapN7drQAzh+6ekEkbQ3xC5YRSRwwWk0dN+/l7TBMu+5kuOBlLjYlerwCa+MMb
UHM3r7eikwKWUXzhA5LPhCmmgNvSiGoZTklTBuJlOP7NYvI1cye0AKDPLuly5HM/QxCvp0vXk4Ag
pUeXzrg/xKV3DoOqk9E/NzpDnw9r8SBOYsAw36M6tyolYzhfs9TiggrLYCuN2rjJJ9oBr8rkHBDG
IWrEjNiqTFhuavdKiHgPONEHB6gvo4kPmS9N8HZKaJihKxJVeQ2Vc34f6zaPsJcCG+eQ6uUmr/fl
FMeyojF49PAGrNNQwGIpQzZvP77lbT86ps+R77YruVBuKlkdhbt2r+U1BQ1PpbS2uQsv08Oi/Jnt
6vbcPM+Qd74czTMaTeXtvtAFxLA2Km7DxJlORmt5qUGY3gsoQrcRr9pjlzhDXZ8I8Y1enVjttZnW
clGt60cu8sWLMpyhVLgWAYDLOep6/MwvrciNob9Nd5THuP4PC0h5OJu5OhFcXChaORoddkoLk0KM
Tqa3KPCc924NCJK1/hBVE97sNHMXtowpVddUJQGIXLIblb0rAfhRzGeRKs6paBcQXf+t0FIKckh1
chSt4S+2srr/tY11CFfMgMz0IWXd6MsSgWfKiqBtDmzbZs6U/vhAd0DiDRMkmFxU/kTXD59PTw/n
Wox47BQW41PinV0B+JIakqWj0aJvdjsnOBS7LCi1BlkartlvSsnRQeWxOarji+Zu1VnzYPKbhMf+
etSc/SuYEzGNKZNa/9SIAZAXfAEaN2Wa4AhFei+oRPJKL+ah3i9Agmexz79z5Em3kNZRauuUoarW
EzhMTAGmMp4A/ZWgzAFaeie1ms4y04Jn93wdTGEcTDWH6ckDuOX68YEFtKj/zuxggAVJIW++E5g+
uZobDWEHb5qdPi9MLDq4a+CmcX8kg6Msnzs24Wfp8CxAEMP420UypLc35MqHdF7Fmd98rtpjIS+R
edtqlbd4CHZTJBliA2x+npouH1InalVRaxAtIVgOYjqg+JdAKAQZCX7690DBT0XZz5Q1ThHrKanW
6qsBP3UmpRk4lyMUbdYJNbY1e8GsL48NgAW3IYHRZhTPj3AHTUZy5tQiAIUlA51WYje8/tChe1ZQ
208SMGxOgNYKKttaD8k7xoZloP0uD9ns3oSBWswI8wbT8VdgrSaf+mh7ptsp/SrCe1M/k2xvyDqi
7eHtVSdatBAP+ruty1RtOsUipvqJkZxA2mAJz9GxdESAsGEI7ip1WYVSIp9gMwdk0bvDNVQWM08Z
xZ7kWVMi/jeLxarae4a9F8WvpoJM/T5S+jsT4OlrTJRrj5FOC/bSfDLHQWYUfu5h0OTcO3ncnVbW
tGvoBbxqu1SH5cDjoEZRqVO76pVlmSLSz4AJv8t0X6UO1mmKjwKTWf3NeHJqYTJUsqT3kqz9EcNn
XnU5YOWX6P00Mfxew+PenHviggr22doN+Euo0hAhZvsHJHbPOxKOBu/ZIpzw9o/raR5U1hu/iDQj
Rnktb94mA+HfwIm5dzO+mkFHS9yLWwPLGD3JMes6mvXEp9pao+7W32Wzugbq3PV43D3zr07xbOle
/ShWbiC+YjTavunl4E4G9UJw8VMNWV0RFEg7IPth7UCDDeQNFwXImi1kRYdAhPRQ0Sn958sP/96Q
wJBgWZODP2eK794SrDH36dui4RHYpH2JcO3FpvnxTysvVv3eSw+5F6mM7o7RZslMhWucEblEH1K/
UDoaGrY20IXQa2fC41G3XD++n3xHMuVgnRZRyXFOCeRE2OIyEgiL4flk0M1AmKqAZM9K2lcnLnuB
Zgi6UpsbD/UmGhhGUigAqJRxihfPdk6nOrA4VBoZirv8ZwMfgkswnatS+k1WcsNiT9BIA7m/8Dlp
s6NFcOL8CTfJbKq9zpoy2e86yrJREakHO1aS510/5Od1uYKptHqZP3QyrpmFAhoJN30VsIHgcrVM
2rUn1tzL5IO+Gj+zhT0gFfDPwlJmCvIWLNVv5nDypatTnZQ1Ur4LG/LnVA+OylZaO7MBy3VLktRI
d7Bb2Z0glPo4433aus5PjdzUApRjKrOkU4z/MnBsJw75AUFreQfFf6AfKntFBUDfukdX2pU1JVKK
QjDoLOoeIYx9rW/e3VCdFPbdFTuGv8g/+zz1ES5bOOgdqYLy07Eb8QrtGJgztyuEr55gfPNaK1ga
Q2v4YEXwhqd1iGYgHHUN4tvmV82KQIeWPRaaz+X3OgTwJsUpYb/iwqEkgjZNZRTiChA34b0w241h
TREfFVKO3YeCmN4V+nH2mgMZKg/2QqxN1IuA0kdJ3jr3to5XzVTGSdr6I7yagTs9yP4rehmDfcS6
Uq/gt5bLRMmHX/EVrG9XrzSA0NXHoG3/gsvJMHIuJ+eSjwhk8kPEpr0FImmbhxX9SasQiAOLf1Gm
DBYpLlQMV1/ZooKIP6HOfHJDfDMWD0Rit61pF1sJAKPFag4kdYnjiQYYWeiPZwOFDISBdMN/nl0M
RpGX2ai0+VK5kVOHITRU06xDqYN/TnFJbWwIh8ALy8PlZnaap1qrHDMYXIHsyG6ymlFQ79Ef4X1a
Hk5fIj60qTcBmQ4msiw6H973CiZ0PIpaZzJ0da6zSBKwQrewvoG623e4/eRnauPfDZIWznHyhFrH
oHP+29ou78f/75QYv4MXyCTo27WLhLNuJB4XJstq5p8vU1DKBOYhzYHEz0x7Vxd5NfuZK+/YqDen
xaX3m/sORzilnhxSyixyQs5HhIJ1vZmFlMdpEZ8EU/OpWSM1XTeTLOQj4UFNCTB9MIoyF3o3rovR
3RWP1WqwzBc7+xtcf42Ku3Y/DNlHmIPEBTeRdc91Y6r3m0S9ylaj6jajCptmyeSXcN/hcUWHF9C+
E3dXpYQXcO+K8En5v2bO1wv/jyL7Cvgmf0XkWjhKc82zNpxGodDXh5GKMkpcGHQTjrTooZsAjkHl
1qM6sVfXl+aCBSEhVcvsqXPtEHoAZ7ARlmEsXSQ/uwZZ0glcUdZAti1fz66AqG9j8cSbKOu8RsaJ
RMXplZbYeUpbFocOaCjJJ0Jjsdx9QNHBhY1r/KZQdgygSlvaApFNdCI+byBwvVsy8wz/Lf5HQQ5K
HwKe7dTNtFConihlST4Y3D4VORW2UmZJTpy3pXDW8+eyoX6m7xCJbhDBcsfD+lNGDBDBtKHUlizF
4UpfPsZORn6dLLtABarwuLPhRpk5KhBcFLFmD/bhRUi+PEnhrFlKW78XoXOvDrMtoricYJyI5oQQ
wXOD08vF5X5YvIke6hMuhI+6H5OEWxRav1bLW2TculfLMiA9KfM3huyK+RG1IQxE1I1orkrqzKnh
GbL8aa4goJRcNhQRPeErfDvmakfzdxy7LbolEbSV92WsgUTljNjkNOg3zrSvwNOLXJtTfPOiE6dv
1twXc//mVg2D5S8Kh17LDYapNrxYrfAYf1hyuLqg8ZqJdp1/DsyaJBrmdS3Fr0XSGPOYxd0jirSC
szdXxmMz0+mS97JY7rAbZ1Qa7jhHdCscSbIj9WmvYgYlVAVIqtYEmxMyYfdgCCESYIxeNSsULPmd
BMUCfjSacmawHi8ozhW3TJvd3YgBfGyfizB362pc79mMZzj/3hj9H5finWwsd4WYq0W7q3zQml11
sqGCilrnuBSW/ScEqilGJCOpbfGoAw/jfgV1D6QsAg6GQj64c/A3+YRoeHwOPiPN+YuNswbg2ZI4
WmyqfHR2Qa7KWG6jT/lVNBrD0D7Ansud/M78qAMOOG7L89ONkeQyS8eP3xTG7Nt39cJ9YNdU0853
TQKCAuMmTj1Vt0KHNf9e2YLhGv3MfvqTI5bya5cq6URQY5i/VBOjBTFZ7A0u/6bMRlKfoKAOxadk
Bi6SuSZ5iUWBcBslCVp47Qy630LPP7rsE688rshn4PHPPZ6GARJHhHJrlpfVuit7yB/bOvIVBUZF
I4tqC1q/dMFsM08X+6Isp/UCrEJNko0y+21sEDjuyBfm1ABqvBXFNRGSzQ5SFn82OnZJGJDPwU7P
AJQyce5TWo29XdM0oUJRLMRAXuy8qxHuXSy9R7XM59yAt8aJExWPs7wbmfPzzrSX8MercBn6Pzf2
AYNzte2eGUoS14oFGUnxKxi8aTdRhiC8WY+Lw3lpQKhXmWWHN/9s7JLs8/ZYnTAyf3rf4ha9sLry
NPTQRGLDjLqJUjuycVkIfTnnp7gFVZxiS+d01ECC1QMfw7akMp3dEXMnBDefot4M+iY4KMeguKpB
jsi27+enfuxVrQ+9e8BZs2krZkCaE3Ubfdi3ILsOZvvtKX1rvMPm1IgaBIaSF0AOhJx9DNzHyWeM
pCyHMirXP9H+QbPKqlDpNvDRfzNIdiq6myYaaGYc/zsZCOVfDiR+tL4yanTrJb52fb+2FTzduiRK
6nu1YdSYG3DuBwGN4UGsrcpKoos26YkQNliG/KQ9z/iDrbhUVso02lOllBwPDuHRJ89RACdqjb+5
q1Z1Klh+V1xglckY5S3n/oRLWzvPoUeRDOte3H+BmyAYFBKyBA5pWlK1+eG8w8sYzwcZYgjL+KHD
jR/rgRFWWganXEwUl5EQcZI+O5kuUtHCsVKZIvr5W1EpkUhC6I4vm2eggo0mUxlbW6b3EaLbjKt2
z3vwutPxLWHf59MVQc3D8nr6b6qozXVIHGeS9zEYQb5r1gOdtyuB9rBpFowfzUpc0qZPOv+oHQN7
Tz873PNkRGp//9urmOA5jTvTTZ8vbRoF//OfJWIYKqZ+ShwHMfFn9NxU/JYvgJlh1yV/n+69LgyG
QHOVLYUzraauMg+8AH8DHBoEiMp4t60BbOouTvCtaBo3CSZLZWgsalMumyy+p6CVOD+/0GFWjpKN
IyYx2GIPaJo8moLPJqGU3kDekgDtTxVxBWkiWmmRq+C1+0raWOdWymM9fSEMS9zhHJari7mb+j6c
3G0+m79PlBOXkzCdeVGLWVOVzo9BXsx9QYAspqzRFGbhULNsDxAIEMfzQIKrgslTiy2ZJKlmO505
J/jz7RRdK1onF0b+EK/TfT3NjnIZU5iqHBgqXEDobJ5d5ZBhqC35J+WDzwCP7+yH4thjjC72zo41
t7XxqBayGLtybGyPWaeg96GVJvirAc/M9bXMdR3h7WeKlf+pp7MmaI16OLxKoTAi/L4l1zd1bHDx
RDDQPmMCgMd2YIlWUtEBlUm5G9iy/WjdeDCzpqbsdANSx/7QF2ZM6VH/rosPJyZyNrexIsp7UI6F
KTBbCH6eG36/nQ5sqZ8eZq6WeAgcil6m7gL3iCwLQMjdJOAum6zWaFCB2GrmWq1SnhdgkFrw5ryt
SnxARLH9SWBwYOmXf8BgEhAgLg/rCdofJBFCeeXw6Y7ehqaNNWG0F/nNaUEMmPwNNrE5NgmjMgWK
rqH5ilhpmyDoNXpFv+t5Z1Z7ikto6a2eM0e2Tne4jXKtNpsJZzPnuCNQxjKyXbtaQxSXEeSwlft+
MOZvRQFWm10MlgrJjC41uVngVPbBaOHIuVgUXLMJ5KYlt8t9++wvZCnHBQ5vt9y1LM4tIRHaCAiT
hOgMUSH3hkBVO6M+SAfM8K1SugLn6kOlJp/Zkyd0Ke4keQClA1bMmJEYhhyS4qYArCb3nIh7IV92
jY75TtPzgv0VXYlfazW3hOjij2azgeYP4y5GehwYWqs5qQAtoXHRxL71vp4FyNfpg/uaeOeDjRD+
WQNOu9FXIgjhCFEpjzIj0AzN/iRH7GCGsQ3+FfqBZN9C9CKjM2x62tDcMczEomcdecAelwlBL1ap
0JQfLrXT/0WMSa6Cw2M4ao70PMVkINeWNaLfUrL0xMwFaiFyhDduprNHXAHODR9Bj12w6fti9qzw
wkNWkGsY2dK60ScQQ0b6JNg/fQ/bxz30d/zcnxW2ucOnDPrlUP+eESOsvyWFQ34R0EPFG9VBOUyM
cE1kmWmS5Y91qhtSd34hKYv6jA/xjVsWP9siwwzMKYLQqRknF4NT9Pb7jnzTfYQaTQPrEjvfuuEM
+IVWQ4/0bzfhyxyJsR7xinxZbT6MY5US27AYYy75GAIzDqCvpaUzFm8zCXt5g2wAVVCZxqJeFrLI
kPUC8I5oiEWbwkMhfPBtpu22y92ok4QOd/6R2nLz0K+OhO7aSYgwlZj6y3rgjHHBODalM2N72Tur
Bw1SKMdzVfenDF9lGXi4ZQgXSLcFplagfOcF1gzNSJjOPd/3E6+tR32VV77/tPW+C8PGrhby/LhM
l8U5odADk28OAhlwIsWW1/nRzfchaqKqx4cbp78pGtN/wZtrePSpsyUkE0pBCjT0J+7PIR5YYPdz
G63EGu1EU3Eg/2D3aEGNQaGk93X2qBJXpwKjsq3lf9abMtz/jo4bJFj6Oapq20eqQWbZ7Qj2ObpZ
fhsWTJyOOeuDqdsBPUW5qn+z8ebNXVypNoRMeZgHYO4Gp/TZkFateT+Lxh5lDml+NMIksPYbPieJ
nHnRm6dx9cHlaM4Swjf/+l+5WT2UogLN8Ha9jrlIe5PF54Iq0o4IQHTe29DG5xBKTBWxMnCQY1z/
uiX9H4WsvQod0/mHm07dzycineRP2ZqTKKZiDc/NvqBQbnUvpJe3W4bs85xS1ZNByvnz0kd4LEq/
Fh3GeKmwWueXOCcyHRp4P3dausH2NepkEpKSHojweJcE+kgxvgPFzn8R3IIl+/XoeNykI8FXrhy+
N5jkNklRFdydlo5TRYFCMqGUw60FXMFnT5GsCIqXBUhF1AhDKWP9gUPKwB8SC6P2visUNd19BiYL
DnsIvIGWOUfvQvOKILafWvc73HxiK89NifBKVPKBo1gVg9oP+rUcNSusz53x44jSTYSyATrZ9xq5
bawe0LKSkDwL5Qqs/b0bMWNDbSihEfWlKRiYUe76wSzlXqlzyZHfLfAwG1pq3H0qjvrAfPru995S
SAr0wjOOrz6zy39mv8ogIKUzkOEPx2iax+MNeAGfKgAVntfty+bQDPLNqmp+Jy6JDzKQYPB/CTH+
oIg3hnzYTNeKLdIed0ercPb1gB+geMQYBc2UUyFInrKdM66Q7CpjCT8We9RSQ1LH/JdEhjn5Q957
htz0pD/yR+bKyQ/3g71ZKLp5yGOEz+jWGLd+KVkncBnFWkDKsZF2pk/Qo+LuePbd9N7Shx6EMnKF
YmekdTteE9ST+gMlAoHUhYC/bq4WZb0jLBphrQbN8vWtrMgkGyfH6r+JkL0mB6Xxxn3+Fpraa+iK
x2XF1Psx89VyIPpwiXHElwy2XzSl4e6CTuCrCqouHghZ1QSG9ymYjWFxYc1FgI3YecpVh83+616G
lEBrsCblnFuJiDsmjDZ/JZ7Vyf1TlFOwM/Yy7ubHnOmjeMsLb1BfHKkJ4BHlDg117J2WuBPYJFJz
s2jxR5rgBos2pDtFD0qMAndINzei9Tb+M9Nh/nmPr7dn0JSwjmvqOmMXNZ8FoBZt0UjecPIShaTn
4+E4B3GCll7EvrQdCC4sNonZEITeYFKdVwAGR20PcGtc0VJf3m0Mor5CfmGLbEvw4r2XdKDGXMxc
iYvoEDctltuy0REzkRvcM2FX8Nx7PL4koRnGGC+3Ce2VRvPA7vIkuyNNcII73frzivQ2xelTmXeT
HwstTTJd9ptdlh+ChvnFzzB/XHq+AQQFN+GEgx0XwoFmqESO0XQyjt8RO0lCVLvpLKPp/r1SKlpZ
EFv/YGR1lWuKcz+Y0Ri6dffvm1zOZJ35VnokfLvXm3a48hvLCI5OO2406CaetH/qYR5F4BA4RNH6
e0BFx3qRY9R81fotrwp6w21LoBLy+wDFDaWaRn8nTJMolIIahcAXEiVyd65vJbuM+ujdqOy0DrXd
uEQiYFTgtr9FHSfkSoLizibeESbL7NqmIS4+tl7APgOK4coQDuOy2Ca6ldMKk7V1NTWnvWS7tGQr
gLFA5raVu09pNDAV+S8sUMA3g3XX38FVI4SwtTDfdIbYQZEfA+xmYGKEKzo6yWcPh5KemZ4d0SZp
8/p9Fk26kScICvDium6WOuOzSAE+WZl3hWbAVjdTK2SzSxB82Oz06sQViHVvG+FQDkc9vYS5knoW
+Zr1zYgPun0xalQ2QVdu/gh3jrTTgDSK1F14I7s5GVHGH1kwJW8C9OhtWy4BRdbjhUDxcUdiBaJT
v3S4Rv4uJagm2AVC5Z8l4s9Kr/IEDEjHS3dAkq6uTbR7FnpWZF4TmUng4Enx707tmlmw3ZiF12bt
5gX++p/N0M412K9H9/iR7KEFNrBB4AOWTC7EDE0wPMWLUbWGzJz3NT6TLqU1QOWfLj+X98cM6pXv
r+05s4V25lxgJEKYmamVkF6XpRlikR53EcT6cCt5iuw1vxaSalnRgUB0tmXpWP906iMVlgBPa90S
N0jBFe6JXRxta/S9lOZOkS6j0b2D15y8CZ9FyhydsjSpL+OkkPQQsxh2r0sqItBFrA8s9hgcm9ze
MfIWZpESj4Hp58JFC0TinNph2yHDg4LqhB8KvS5XN9xhLjLj6/x/Ngk0LCtwWPh0PM5H6+0LkFDE
Jtl5hO1Dlc9ZQKluPG4URpDCMJbofhdpjj3qw7PMGDrfu/t3h6znVlJE28Kty5wKO7O525xis7Ad
OaCVTEVJpSXXSmbn2gq6hisNWjWl+2ou2nBWOtoqfgTFbUDr19/KKlDLRn70wiWayDvzE13gqZxj
O35sMWic/oivkcxRthk9G9caX/E9tnumdynlEHyWdbHJvIeEoqsxhO1qk1CoVkZCLLxFqRG0w8Yn
yvUElUVT/nxPemIRTfk0xe5qHZ/mviD3s65p+/gUKGIRI6/96C5Ll5b6Fo25mZlfjg0PIEKpIxWT
7g2JqTWjnjzMRyHMyBNl1mtAAbVYBRnL4KKihmQ6uarnF1pCT5ajaZXdfnv81KZsbo0TQw+uLL0Q
Hc4f/x6fDbIF7ewjpnAtSFJfpkJasb98qxbbj3TACi6M2HcLxv0BS67AgFFErivQDBpbNnbz4pml
xboNSRY8yTzrZjsIzNLbYQB/b6CDAe2TOeZZOCD3Ysxh34XT1kjWlUkncUz9/qRWmtwZwUr2NCSd
zd/lckVBksIHBk/BOC2Ma6eNLoKVuNloVxCzRZI4t3BF+NVvJZhJRa/jskUsvKNk/K98AJcqO4ZJ
MkfOg3ude+5xn0A/jhmYXN7yiEMked661bqX5Dh9kw48cOk9BqpkGmjAqzzp48wehpgX3deKfbMX
d/hcwxdky1Irhqa+vytf8cV5TVEbDdhlC8wsHIiwKpANUKQzy7Ke1aymFs75+So2KcpuqvTTtn6A
cpqPKluM0c6Zdby0WoBdzpIBcSS3j3HsqJG76/nBzdNVB+lEHqOuoCgUPk0s29USr5qwakplesgX
CvPScnIfsIH4v+Rq3OPtvFOCSLyUKh7IDOilINh8+LrK9Y46YwOleOsh6C2DGF/N9vNAqjKc2JDy
EwNiIPuSOU9gdkM4yCnk5KYUzA0eR25N/1ohce8wp7Ne8bX91LjX5wQsYwEDeTuUfOBuWDlJRJnG
KznSSGVtJBKh5+74E1NJ4iW7wx/Gv60bKIeN0KHlws3UJr30rn7FCM3uHrHnUfSmfBSUgkKeybSL
2har8yyHqhivT/ULe5OcWWW65Qx8P4Nhv23+KMk62ucVtwmh7EFAnLPLC5dD5SuYOfPtUzl2Awte
9KFyIUT28eYI5yVkYeOCOxKtfGWsxHYf7264xmE8Z9ICf92AKU3G3bZib6/OaTiFX4PygB7QyQG6
oXOS9lTiHLAJjRO8NLdGW0rxD/VKbVv8BMjHZdsTDE66z1l7s++kBQInrw4OZVBhbYrqfuBEIb9i
bhOhQvedVm1LADOL73nZxreeGcsFduJvc3ekyXcthLPIMydmgVBUJyuZdMPKFmvMnOHPwQfsPJtv
3vO30HSMi1MdqyQNCPxwOfDGeW8X266f6HPK2ue2Z2TnoCwZWmlfU29NnyL1/+9iiuxH91T+Lct0
MLbjKmHI55xXAyw4a8lqVTpBn+R8oy9tXOJU+VRt9fAGbiGwFmTYp0xZNT/JPj98edSNCCsrJJSw
bJiYJbUjX22wtiVKjA711lgE9LWO2DdTAFoAIbNbfayAm/oKq7eIFzl6k+5phWz6pNX5IGs2AhXd
sy2V5Wrsd6zHvUPASqcZuYVBNEPjecgRd0fbKzatUWFAUR7zladF+CLpyfACM/H/f+w5E8hc2n4S
tdSKS67NQoDHPKnYZvN4gd6pP7kxT1rIN7C95FwylL5bGne6Fk2CrNjjADGT9u/L/ZJZ7nL5Tcak
7oUt6SxQ0AtHhGCEcZA43yRHoY/QnpAyja9Tjeu189hYPjj3ois8Cfc4bdPFrtqJKevE1SZK1k87
6CfCkDgcZblKWMftT16LFW8ZcSmkHVOWr8afg8wpbu5nl1rLe0ok2z3tIkWPQGhRy0xzrsSKTtpV
NMumfZenqU0Fz6DUwxMPp4qMpQLL5QjRs/hwv6+17jYGM6nt3Ka0aNsGG/d9kGD09QEn5sp67BIt
V9loo1P29Uj5uQ938A8I6F0UfScnls7fX3jB9oeQcGBUkhjYxF5kvbjGxMjpo7VmUH0lHsN7mvKF
ByKi+p+eK0Ku+Y/JX1t11wXOsFUfiH6rByYx9hm9vWzqm+3tmfi0a/JH8e0/DRLagno5V42eR0LL
OcSymo87AYFrO/wbsPg9jcMgi2RK8R2jHEUDbcB99aSomq+dRYG69yLrwNDD8u6Pp40a6a32/vp+
26WkOlg1PWRWgQ5HKqMd3js3Xx9s4Jj+XRpIyRNksF/QQTQTV31PID2Ur/185ulPpzYKKBgrW8oM
V13g6Yk+gCe172edVY+2CzmZmmiD1tCOTrfPO6dg/Vwzaklbgs8zvypJPDp979SkGjzS8RQJZZb+
8phQ+3n00PRD4BgMwqMW+ynEiYvdeo1PrLV4IW2UQlDZuEIDAeINgLUxLXkslMutEekFBtiQWV0I
KmTIC9sAwCpI0//6z3HbnI21/Jb3IIe8eReMER/hHB8zE9aEToV6OiB4M/Y/IVw+0Z8QEXWtp52N
1B90XwrBRiW7/LrOoAMM70rcNDTCTywN2AbJVzDLogd160tRUDbhBojmMJx6vtNRy9iUkdwCBybI
HLTRvwkipfMSljMEUcR39eJ5AUxmc3KJSl5L+qpnahu2BXcMuYlCL/JA3u597FU7wWusptuR9GJr
sz03KLSPQNG7mAR8EmM02zg4yO2wO8Nlvpi6W5fSed95QLd/SxVntoofZxFNoipDBKs6tpPnO2rH
Yam4T2/QiERgY9jDcon+ZcNwNVhAVcX+CnoodZhn09Xrm0G00eJX46S0VGkV5460ekC+vSCW417Y
QhnU7Ke56BU1JQD5+GamsEm0CTm6B0EA+zQYRB26U89pSYTuBnO4WLBa4YSk51pJp/I9RcXVUgFC
2GiJUGVhp6LmQ/orLPQOwr4cyGC86CNaiwVW83dlQBAgNcx+lHQmQYcdoFqHDeHTNd9Amvys7pF4
h1yjZ3gUD4usD37XZKraWX2Juk39JuFesX5ZS5wtvrFGE+L+IR9uyCPfWbWPlyCaQw9bzxHy1J8l
apXFSo0nb2rW61/nvLd+kOYliOvj1fMVd8dJA8HVnZhs9YOTRFtdVkQW92wm+sib+Eh9x7Z5hpgQ
KM9zi+bVYXdoQPTmyY2XMnrzDzO5cLrHrhYFjXouhpTCT7Tcl0L0cMdl2dxDZt9qTJPJ9/unwW8Q
9+aTonNCLu0PIzh3a/KfEMOuz4boF+ijkRcDWddZoeG3viUxub0KL9EgSUAsg+QM8+5wm88NtVVP
PgD/48AUXntLcHjDCQqhbsaCbuVTX4EvXGuTOy4WGqFyWb8WdkM8TaCHlwCuQRwSqIhgC/FQskCz
FDyVtTeQLcQqFQF6m+yyid3kEHuM/8c5cdtB5vZLJRDEMwWO6d4ZIVtMkgnbAzU8aat5slV4jSGi
mIgqRKJN36ugakW0KYelkdZbOiD8h3bLnfbbYGg9Yic48tb59ry6o33YyidMH7GSXidNj0vz30g4
gJCpjeSZVUTAX+k7kc1NYUA1SNUmSsAJHS6XnuXdWzIOwACp2LyzEA3hrTXouNhWtPccBOs13/FI
TW1EXwGLOxVnDDGUscNwAMRH9UmRQTTV5uPvosktQbBRPPLE54ggGjp7WlTvtn7nF81u4/5TpAhV
cTifO+o6lof/DHKgWYjvrq8mstySfA/7ZGHP763KaaPC8ae55qhLQRPZ0QTIPrOIdrlRx6kkOw++
MZpvpBimsBAEVMimZNnMdx63LJIeNXfWjTMY+UtxOLYamNdgGRkLC9wLll3Z38LmHMlLN/KPkiNR
X5KhI2VtD5yRI5Cuk5fBXfPV4xW70j3H+OPl928EtSnqu22GQyTOkZqegfPKl26kTS8T3KPVNPai
rS9yTvAm/y5ZUaCPJWLldH9YqT4wAwPyhzg9ZfkZoncFtlUVQfdMMwvyO15iRUCaDM85IKrKeGxj
oz7/qmdjRx48JKQRYGZHBvmsnSmUaBZC8bHFvPlvBSmLUjf2vak6kJ8CGApjUCjSscpYGZ3G8VpL
mcwuhUy5suwS1K+NaV5+swX5fuAlETZgNlejCrDvCPdgDOoI8Q2dd7dggKy3MMXBAXAECEm4nA3K
RcsKHP/F8vruaoJwstGyTGfYh2e/9xpiYjeg87a92j7cqhIWbySX7P+ncQ4WVwE1Nu9EVPM79IR3
0Li1YYjJ2YxqQsN92WFst/DF2/udZ8Rmql/HKIK+5ulDUUH2X876Do1eRGSweYbJm3s9u0kXX6iL
8zNvQSK9GLuQmlKQSF0CXGcnCWLxL/mULA+0BrJa49zua9+0K5qZrq4PjckumDqKLhg3bNx1J8oq
48PUIrjaBjasdCQybUHV47eUT56GzPUAX69snzcUvb+0wVQvkFChpJZuNruEwaP/fXnHCTuomnC4
6n5ixCjA8ZeKfFK1qGzR5yBitRuE/+bLkRY8q8MNWhKHqJdicH/ws13JFC4f+TCI5IOvn7tKaMVs
yEW/xS8d80CuHR8dmXd4CmcORUZsxtv/2EZLwTjYSTUExsX1Sxwp0IZYszz3HtIkYegYKG0MZvnX
JOKzuG/Eo6I96+i0FjRAdC5g3w3A7YBNsGC0K9Tr0dzc+MM59eArUlIOya58dDBypmjQH9YOgzwr
Fpx6L7aJCmjnqaj+/PZvxk2HVnmObxLNBy4HxDrINFsYxZIhzWUayHXUQZyhlW8oPTQg3BfdZBOR
RpRmZ2+KTUYqVJFQ9dBBBY+uwFNUUBv1SrLHtDocyxw/KyTwp5vrxnz/7YRxTfUkrUAchMxAwhz9
DhJZEfZTAtcxp+Fssj1tAaq2OkuAWh1pYpWnPq96/GKC9EuKeJOkx+lJ3cxyfy0G8zpep08Zqy3G
ytHmEjLONMvWwo/GuYkbKa/qbwoVcHJ/xokM3CWsplKpCJ4KkLc3AYDWSZP9cwXNX/TtDnDqF3X3
IesKbuo/5T9xKXHpIFVzjZ9ycThGpfBbMMiT/mOYqhEDnNYxFivkuVEXDblmqM9Pgve86GkKKY07
I0QTYz2NX0HmJ5vt+2IP6M9QtQRIuB50g64OyYvu7Bk+z0WfKiyVFFqMVBP/GOwQJKGqECseY8C+
Av4wsVtbPrNWjo5g0aFYSMACDwd2NjQaE2b6GKQPxCAygypzXIkxAlBMEdwGTfnMWqTRpS/0/ZXj
5z1g93osApkrt5YkdtPF8isr9LzndI3OT8KDyE20dUshwmmzMZz4MaFOX9yf4ubEskXW3tHwqXm1
ytjQUAV4hPFOXIJi3ZJDWOZCzIyi8Ccth5xOZ+m1fVB1sqph5sNRfmAzYpsSyHiIIKMlemOLi72d
wpeWdbeS6PHWHXRL9RVMWQMCyE7LWm+sRR6XBczfhbxG2Q7yZ1TKS+BFTjtZjmGwFdnMp8mbHVBw
XHdJ5gkgCvnDRuThuh5enrpgGMgazHuvgNzjLOev+pc+Oy1wL6U1MCKuuqjlElT0wMeDwNzKb71H
fx3iuyvuK4HsYO/UVbu0/+wddfFfne0KDQp4C3dqNfTrMN6wgK1sZRbAyv6HCYfptmBs6gGsbil/
VQVqVRCbeN2EGhZ4PJxQIoXSSw6vRynAgRp7Z2hg1Uwmc1Cb7tc3Q96pqKrj3vgyqFtkUAVj83EA
2S287JRUw4Fl/I/ORtyFdcNOHEBMf1c3Y6+kEkP+nZ9bCYMdAj0L4Vh3h1sXrIiIZG9s37lXlPtv
gzM8o05Z7SAzvLQfi5vHX4DhKXd1SHIfSJ5xND5TMJFEM89gFy+2btFtA9fqKBCrXZtqtx6Tc0d8
5razuCeMogy5XpfoolCTX4vRltIwV73a4+ZuC81KGdi4snwUMFlrilHAq477oYxA7EVZyQNGmFyB
Eoq4le0aoDoKlU+VcXmucyYtSWBXXR8v4rX7O1+vlnA1NAvQfKNSVCYRt/7uuYWHhuZhse7BMUAY
6pXY7S4hrjyVWvVlaoUFm0U7nsDrhIQYEIADztNG8KeO9o6v182gOFDOa438zPtMaB0COKUmVPjo
l/8G7NLRyK5MBBHxq95pgezynrPKcjCiGnfelrP1RHjn9COUtH+UMDFERsF5cvGTwU9PLZPo6/WN
lRm3hJBA+OoqKDT8ZfOLggf0ch1ZYIt09lstgR7SOKS+zYbgbAbQtww6Z5G0KWGdKa2S2FHoIDUZ
gbkUhbVwnQZXH/XQSB8h0Hk8jIlG142w3fCXCiDpuqP6cCUrqejrgjjoBWtSI+9RuAmoVlUQt/sC
HjpJN5bt5mQLyAUqcY8Poh7DpQ4vTDSq52Tc8yyhhJZHXqU/5tysJkACctrmY0bXFOr3I5iXin+1
ZEuEndS1DTqu9yJrSZYuVexxHkvs6usMDNzGWVazfnbe+lt0s7+pBCh0KpfjMfLBnR/XcpC5Zm7G
Rf/gGq1gnnDlVbF1mSnxK4g9OPeI9Tba2SxQW/AkYzcvG8vgxDWR/RQ7kxpVgkk069hr0ddO5vQT
ilILywdS5V2CItDBvYNQle9OzDJ4pRo82zv4UKuBO22zNEhhXR9Km80PBIB2K1Y1iIdOiPZfk0vM
vyjUvL79EvAS74Jv4PtTPPMrUErV0F1mb7DEN8MvbJRBbFNhPBy0owXkxYsoorKNCSyrruSXKb4r
9uvBbDSp9c/q+u0Ctc2SAPIP48itKHo1Xq/Gv2Iq9hHhEg7OKjKQ0BfRT2obh0XJjsbdkAjn7HYY
H8e2jcXLYuEImDzvCg07Aos5GKrrZke42V5d2B3aDNbDQoXjrKINJQNrIWYbfrLkSYUliU1xhHG0
1mq/DxpJ5N4biz/KV6UjBMG1IfO1jRtH9iD5ctqwdxhKePIbPPStEK62oF6ksFKxlnPc7jc4V5nS
m25pHP2duCKOLD5SpqIbAmOf/G1UZ302Klac+mAw0rR44ya6kRNBkSx8ybw+JXizJCUSgkqlw3Mo
ZgjYcmzYlGB89pL/GIJrDV0c4GRs5G8NdVvpUp3vvWfvjzxrXcOo9qHWVAQVRBIl/e+bqwOACc6k
23Pkfv1SVlnSn1CaYAKhtFo1Nu3LVNhcW+tTO71aACUbY3MPDm1UIVMJv5L/Y2FKZIpdV6tT+Ure
teOMsfJoYNGsEyCW9rSfzgbx/zzzlsAFZ8P8lReqsXZ4Vt9SesWlUccID2Af4pt+rs+wSz3LMBmo
607yLJPJyC+nCP10b55wN2Yj21oPZ4sVlXI1G8nuLdyMgfqZXYf1dKzOGLXRpWozGeR3QTN5AnUE
LfRZ+5wHC9C1N+dRcaM09hhwRDGRN0zzjyCJgfY+Wor940UKKkwisx2XY+ksNK0SINPTfgTk/JYP
uvz94tCuUx3W4jEvjZaI3hei4RBEHHW83m5nZuwv/Za5dn/TiJeOxaIFwfHOv4jnsgoQdYgWBiSW
YleWvB4kPYyLfNNunP0Phve7y8qPh6wwZU5fmQdJnpfaudjn/ho9vsnjraCsNb9IZMkzWqTvHk4f
ZN9LQbi7i0EkjA9e0PjZOQZOMJNtsrQv3OYSLWZT706ATdWXK9aNrLbsvGtlizBELNgMdSy5LRaJ
0L8Aq6yqtG/EpgckPIfm0hef6t6O3Gc1fNgIptSxulaJdjsjJxTE49GbTTw25ua4ZYXBtCrdleuK
HytB2ud7sqVDg2GCXfIbxG99ek7bePZH7TWcRtZ0XH7Lc/StYCjVRe6R/Dg1xa3NGEvEkJ2wIgUb
cXB9jlSBKRDwXRoNRDVqfO/WegxtiAtUwkXCP9B8jeOoDLnM1QYApch5QdeNV0R2tM3RgVi3hXFz
OyM4Y7+m4rRWnD3Oq3Lg1T3Kzr2HlAV4WR9ZyHNqbxWDgD99kvxbGzptgnvuD/G+zDwd7cABaVFR
xaVKrfc7BccQcA7gn2HPTxqhSrPRb2UDvD9NZZyVr3+KPP/2bc5TAbLT6FuE3NAcxQL/miNzHEG/
smUsOMAUX+GfHPg/FNrHWM/TFqP24h6JaUwkEJEFuydbA4TEBcDOYmjjTHXgKrbwfrVabdIDeWjS
cgXrh/199Z+PFLgWU/W5h8R2N0Av/a2Pnwpnsx2sF2Yq0AK8wpLaOCq3wmekvt+ejqNVDJheMATl
RXUf4URKURR8i9HjvFiOt9xGmV9PeheugNjMp6uFrPVraikIRR3GSVpP+GyvpFgSDPNYjiSRLNgg
QlbMKXVGnwb0YaEipPhOf4N4hmyRALX75NMXnCFx7NWdmstuUQKKjzfQuPc2hmzxe72E0DufFM7I
668d1dwAsuij5RHt0SonEma9GQoqptkBpwHw41j9qo8z3QO423ugyM9krcHCDRW/BOYT5CFhPPTx
WkZyPuHW96N9t9e4Ho4SmnUwL+NYCD2nia1JgDhrljPn0tXSlMlufx118icrtYVVaxuZcMRGc22g
nlW+AY7hcBwHCzMj0rvLUwA1D87Jjjl48eOurOBV2Ma8hM2g8/Fwcm6wKGHnBcxfYqiP+aRhKKxy
0uLXUYOW5gVPiuBKypOZaPIPVMSIEp3pKYdbwKukhuG0ab94Xm4l61WQMdLKKYtnZc3EhnK1QkyE
A+KGOnIQ6z9j5oVrJBSEYBuj3ei4pWEIhO5A2mml0Xq4/LaCGbKhVjI8Jn/x6tMJye4Mrm9H8Q6v
nZ7t2wmwSM+kSm3y/hMq+ikgf+8IZfM1WoruFWPUSCkypid8UqGG2jONyjMQRvNlwWw6fogzPRkL
pfaLWTgQ+LJpHTGY2Jk6eoWms/N2JW0h6i+h6yMXuK0VvrFNTXoorW8JViM5muiXO6h85FcoWgi/
xhG4gZfSOHHYELFT4n/CfKo77YZFJ2veMeh6R0RCX/tcnXkPC98rVmVUTca0HRvZ97VKo9ZXXfip
R0FQfvHZ5j8cE1qRtRMeNXSG+f0UQiMWDIeSHV5PVcZsoo19Yz2HCAxuojHe+wKN3AAINJpwXSYZ
drs5MpME6qEsYC2HiNoJClo03pHXBKEn5WTzi1MfWW4kgQoouKfYrtDBSuCRCHQ0m5soIagyk89F
VrupqTa7t9XmGIfmyGwBENBncGYd9dBtx79TitBZFYi/1ugC8VTVyBs8ogFjk5tTke5rSW3vI508
XPLiUpdHVJEj9EvLKB0P6oh7YYTEi1ETlgrqA88LQf1AD5xDZ+hsyFJZiPd5sR59aZC2V3RNAG83
p7tCn1iLqE0HOc6U1mXv3KyhGi1O/4IaIIt/Rj+lJEq7mxFQwI1HAXGTcXELKzTuy3QnDiANo4ey
n6k9PfvDNs0+fCVo5+MHVJRTVX0CF+1b0OIyR7WN1G6d9BXq9JOdNEEffyOUCzA9Aw56eUNZvgnm
cfmOkS6X+q2z9izvLqkCFbxdJXxfmsgdZSbzCTnh9zMKOln0TDe4goEkwnIn6Qlpm/Sin6d7qPKb
CSpB0Youn7zzB+wiLYaQ+f6xcMZd4+/M2imLXTOY0TvoZDLD91YY1pk/c/6OcT4iBjqe6F0elIFL
ccqnZD3RStZfTJwXMcThFl/VfmZPcO8XkBcxzYzJVv7BYzhnbJH9q9B1UWbSEmQzH9/qlWZ+q4wk
Ybbm4u1w51ywJXLZnsQS5Dt6ZIjlRrKCULPKokEe5eANZ505YpF+YRz/CJZQdY014Vqr8Jd2zMz+
S9jYmeQKt9mTyCOTz8JPlPe1zGWon9frZ6UaXqgg2oeq5i7gO+tPHal52axzKuUR1yC3Y1TW1+me
8Vi7n2BJYCOOkN+2Q/fTTBKVMlvQyi41iiXVM+diBSarCBky7HSt3CIAO9bmwAByGWqWNxioLm5k
zQEKfAqZOpuNUrvXCyu/gV5hjSKoyc2g1Jev+rebS4HoqDBKtDAPc+QdbvJ9oAGXuMBB6Tl+8Jz+
e7DgCZ2LKjWoyXD/hD1yhl3Dw2Tpiv5dksTV+6SQ+qCSX+9FGyh0P+o0c2mddu00Sf+bASeccj0o
0MY8kzNF+6HFbhQULzllEWvnBEzmL/XbZ7PNP0BlM91OXae9uz/IMeR9T6iP4q5O5ehvtDM9Xvos
EAIYloij0TjSCrQO3oV0b3sZ1dJB8r9TVEh5rHufrwDNyKVRiudOHVFwBJGB984AZU3QO6Okgol2
RU7cov4//garTh5iPzpCKbqvsKSUsNpaO8K1b8dCL0gppBVQ5R4WHA0ZcbSTnGTZcAOqXLdqKT2x
CAdU2sK7Bj8bqghs9r4HSD6i8zbbv6W6IN/JW199/oNnbnvEdwhq2cV/w0UVT11AmzyMSyGQ2CYB
+/CrO5JrSxUtuRXZYt+uiWWD3xmkV/2Sa9rhaFSm6xFNjM+4GGfutCO3P3p5eWiL8ItADs5oyzVT
xid7+PI2nSTWlpTKzG2lkRJ2jYXGha1ukBf2nyo3BeAJY2U01ZD6Y/eP91rfRcpgVOtW07OmF6D2
+e8l+0MRtNq3qemGIhOUizsfbbZ4uwnIL+U1BzirOIjiyM4WDWrxnDiGFXfyzSB0cvTYxxfJOHRf
nCHgAzCMkI0z9Dbp7jYbM8w4jycqdPzjuNhNVFxK6NSfAiQNtm+aSQ2hnWuvqh1fwka7zD6GzbFI
WLPKadAF2rKW8PmNCFijJkY0l8goiKbi1PAhELav9Rp4XMv+ar+o4zRjENTn2dc2DTp4lDHxZVbL
KvwOqPNyzEPZHRJD+ymac7havtr8TT8P0KDaL0zSob6hL2VF8qYDPmrqeoDc+oO+PdL67CftIxJQ
4WFODwf/r7TI4J7yGzJEfhklSQUXp4WU6nGuU1nZZHBDO+RtG3Nb7aO2Y9VvlclA7VAmvnTc1N4L
dT2t9sgf/p3RhnOPovaHmu3px7VcwoHn58oaJWCYf2ds0UrZ6Z7QKQ+L1C01KkHfJn4XxD4gLcmo
zHwSKzwTUJZuwTOwjap3GyaGdExJGiwAiKqT8wQ1fyUSPqUP7c5vt6IA0YZKLMfIYH/ia0Au2R2A
CKjYYJaKwPXQg+Dbf3+RTrcOs5aqipqxN2hmtQWWcxTyueb8r/B25ASf+R7VuJQ6xBPxGkBy3zsc
SFsFb4pJ8NeGbByMpXHRmRIbCLwZoGLsZSia5+1/ym+zPuzJH68/fZM8IGjKZutfMzM1yoro0fZ2
Xz30v/BypKAlinYIZkGYy8tN4dR4U45Fqqgre559sLjceavPyNU8PQWg7qPdboWz2lRtAo9Y4ADM
bEnD+Fa79Zm4vgoxKAvjejlalWkh5GW5vt057uxbqg5Z0aNW9zpUtX1RlDquk+MrViGCvw+3gI+f
Z10aI1pFrUjwTdzs6j/iyrrcfelWTyk2SKoWs/STACkXuIEzaVXYE3w3Y9oB/dux90scs3nf3vOn
MocutorUp1ppSQ0Z8suKwmb/gUnqq1TVFjgnsuQ7npoFLFPjAd7G9jsoZze17o09Ye1DM9oa0/67
GqPlQsU5FUEnYcx7s1CmaU91qBOIv5V+efJSj/OHB5bfPQJgw2ZPHtev4wcdSWIwoqFFh5UOlkRT
nMKqaq3MvG5U1bNnbHFTPZ7s/tXdGJJjyBtX1+evDqr3D0/mucJaKiIsPr/LIVSyJlan2rFrZ/Wo
erz/JW/Z11SIWX+XlFw3hAm55qd+mlB7XHXIv8mjklaphbJwvxtZ0rfW622IaB6Fd/XG5J/WMGDW
XGWNTK9w/bswCq5GdI5HySc1a8B4xoSG6fu93GzbkBVgyf1xsTad+9JYsfHepieqvlbxeybakNKF
a+3FHqda+ey8FpOzUEYuTk5+nSJRXI6FNue54na5GL+JQAaxz/EGhFeBXCv8MMU3U1rpWidXTwbW
M5ZRW3tJXMeSG2bH5OprnZadot6UEuarWC48J0iAECNqXa8aRM3/gVl9qgSVL6IF4Q21cdpLyNFp
g1h9u69vDtI90ZHdJsscgH2V2awsS4xRfuoFQwiTbidrmBHrIcaXP3roICUA0904E+2YvvJ8tcgE
Ej6592GIX/F+mi+/YTd2YRb8JXsPmq/nEcmd9RNhiS0uKFhTnCdM7oq3QLNBwgA32XPu7UP93pGP
GEGjFVm0pjptkqQhtvUZE4rYf6ij0yCh3PFzztaliyBzIfsleIe4O9e22Tdfswvk3CuJQ5QwQszF
jPX9aaKu6vuksgZ2/RWgQIQjbwwMAQdiQU0DzcZ1m+H9w5qkv9Euu2B+QdR0mc86lZag0Rl5Zo1p
K+ywKM1oGK2CV7zwOk3QtgJb547fmTsnl9TxlTgU01qk2rkwzMz4IEj+GfW1ub0r1u/jwRgnsA9n
GOEGFKqGKQYgPY3rs8jjxs1GAuzJ2gW6dBNKQp6o3+3s8qPe1xcIg2YXINY2Qcc58lLno6V7Zwyn
FuQKx9Z63gXXF9wQkG2NLrqXROnw/dFlVJEUnVhcck06qAt3xNaDvO/+SGnNjpDZFLlFoRPhN3Nx
5ZAXSDT0flXpr0DCNweqiHRBRZHPVC6g/pTPj8uRmII6YUn2Q5nmoWPVscV32bSro7Lq+9bOgS3T
HEMHNJoGJjwdFdEM3mEuldS33HvZK8NRsQp/m1q7bMIRlW2FeVfXVS6LTo934Yfkmqilb9mIMjMg
d2HtjabtZIaoES8EzgffnswJCvOX8JiDblKhjKzu17XWsLCQSHd0x5DDjTo3q7VAkvlvntcxtPbn
kwH8cSZEBzof2mHvwqt2cl4MheuzvAK6P6R/L17ZRidPTKTbiPYF/gRt2W3dhORyet/o9YeDZh9t
j/qdd9GXBJh8dBnU0zWSCVuR87Xu4zWndgq7oKpnb36suexp/kskdyjHlT0OAH08HRhlATIe2ZKM
CA/0f+Z9Uwko2Ks6KfPp0fxw/bV/JLcfsoZO3Y7bZ6X41GkIL+mbUbISRiYtJ2ZsKDDk5DEg5bC+
cLaFMSBcj97htLI/Q7pFTBZ1SqXgjad9RqG1ik7VgkG/VjTY8IwW4Xs3gX9pJfNkzSBrkyvohDH/
w+5RE2dV6svBT1y+LHfJLWaqfEgoBxoY/odCx8BgqlpV969hNROTNFknc2Voxco2fuwK9YItS3fi
A0O3L1H1qI+HWYYZ2AaVXbshtBsGUUYuV/SAkagx0Tu7iW9qo0HHll9d8ichaxzqS8p8MUpmgyoz
AIyZ6sFKVlDghdqCKWyDVT2DNQG6UTmyRScNEHHtsntFRFK+CAU0YDYm8CwFJexFC9LjGbIcFVjG
+ZZeOuy9Qpft+qJdGXGXSGoOfHkh6sLsWD8gMD84U4d62YBt66aFseH2JbG6oLNsp5qnmfBadSpu
6pfb1yXKT8WxM35zGkoD9EmCIR23LhtZKIB0lOxyseYTtziG1vSC/Tr0+aOKy1Q6RADAFNFSkFtE
F5LvtfjywX3C9W2s9r2ypm6lt1a24DKNVK92slthLoeaw6No8wcMktagO9xAKK376iSjhVwffwsc
Y24YOZWhuiSN7eiK8tvtQUpVM3CSae0C4VwGNDkCywty0G/Zdf3i8b28s2GO9iIv7WwJJru6zf9R
/A44a+D1uFeH30hiypUwLcXLh1FpCykGIaPsbd9zaVycIy6adSRWZPY7EmvOxrdYcVjJ+hcDxJ4J
lZInC3QwiOVLLXY67gSx5Rr+OHx9mVjvkWBqsxh43FdUG1Jpz7xVY2uYfOlB7oF6vq6+LoZBvbjy
d9Fwiit3aYqNa7WkMcx/P7QpLt3MpO1ZAxZvK27wK7eIi279qz0RjYLm4bVk6WM1vpZnR3kvbPVl
qBOJloPi3ch9+1XwQGR6IQmtv7odK2mhcHfloF12CYoS/C0SHdD7NZW0z3v1DVGrnp1crmuo1QLq
GdTKRKqpekOiEP4MrSTdjrOcQTIKzYvmZJiSfOMfM5CaN3WtBFuD8u1WsqwgokbzhqbfneQ1Dn4g
wO2aM8q/h3/jSE4EmBs4lk3ziJFcEHGp6oQdCvzN3mGg+vYHjSdA2YW96C8q1iS0vYfNZHaZLvqd
JMbVs+9Dl3StV0ww53h/zmD7KH+yjMVCKuHKPnQbUnOV9HpkOYBfZhKyGoo1CJvh5aQe/9BgYXZQ
fbhaQLHoMBCziEFifqtnAEHAWWopxN6paj7y8Jizq4jJfwCPtTsci7cXE45u7xKZ3FtXZ0+eELvW
N2FusL6pKEFov7Q5dfF9mvVrFOa4u3DQUcA4SLEUOEA+HI/oKyhJA2nsY0yYdDfYKV3HNBkTNLYY
TgUl4PYh1LlaDrmlpWwn4XwXL4Pdrw+QBphI8r82aKPaqM97rlZ8n/glX6dH6AprVW4/WM/GNVSi
48pyA2rmfarqNaCLsKnryJ1610KdS9B/p81r1ZdVtGNzUS7D5M960z4RvqGSVbmpw19HXvAbczzk
XbGTuw1qPNjIf0Dx6+JUE0MFZkXOyWs8+LtdhR2ed1ffR/toBZAIosvLEYivQ8rEM0ovqXgSYpSe
nXlhEET2ohTJS77zj1ao/OxiPOdBg0fjkjy+KuplVKrHPmFTBGNDaSU4ykge/7HQJ/otnTuOdulb
KM4Z1iGiNscpOdwVGqsM84115dWdg4cX4k1aimJOsrl07RoXOyOcmNcFjRl1uL38xjXvEIxVapp9
G1JLP8bLCQhSY/PnOcfU9I3GqFVyj3JCHdHPFhPY1FIxQjrlqKpfB4k7x7EnHkdEsgn2TE7R3jtt
g1WWHLUKJyl/pBFv+GNuJMUNUZ+MiizanpmRt/tKFzNjFj0YOWPM6gAIVjUch3Y4pSBdI/oBBQWs
ICPcXJyyxdgRzwtmFDftZ5JpkgRVyUVPDiCQ8EPzo61+07rcBaDNMc4upMuTx0ddrhxvVmkfemMd
z2iZxWLwV1hX71Yxql8rxdVF5g/KBZmBvHmR3hHeUq6eK7TDZGOt4IZnqN4M4W+3dYrWLG8GwHQJ
9QmaS/r60e6qzHlbLjpvCWd9WMNqps0HAO9+1N64ms3jN/zTqmBRXvXo3/gc+rtDautdrPK5uc11
O7jP06htkGkRPV4PYKagA1+4Q7dehi4b3rdmI8GGh1pcHaDbFDScB5Ruzbg9t2Ro2d2FnnHhn1K/
p6Ce8Y8R0JM7q51iRFni+gpFEyoivgGYfZwyBSVBvlHVhWxVnT1Vgo56Y1hzG3mDjpOc+LhmoXPu
JnArPYNtlA3BHzKAUOi3SJqIRXC8AVVZefjLPZarztDvcbqxt7ylApeq4yDKUjaGjSfZCpKTAkIx
2FUpR6YQow9JZW2n0nmaZ328Pex+tM8p6mdLEB2qeqy0RXWfrJrrgIprbYYSbeeQtT1+ifawEXXv
eZe6aYiLCgQvgl3JnfFwDbdkI7r5ebM/0ZewfYQd9rhXYBFUmMlSuqp2Cb0Hr8KHNvxh6haY3p9M
LygGFqa4gzP1HKwmppjdZbiWQjmYQvEBZYGR5YOVPzZNAKhbSbvbsxjyWrBEgVe6NRyzZqElymSv
hZHYg+Wj5/6bNvR3YYpl+3lPUxJ7qkqQI1INzD7DS6ZDr1jkrOpakS1pQi2L/OATZFZhvjJpB3Hp
ywUd2OydWVS/le80hbIhFa+A69kvrjkUnX/0j+vFFatmM+NRnBCI8IymxDcpcyPKoJ6EeWPr4Odq
RcA0oX6laeQGZWb7hF0TedyWl+hmEa8vJQiYIGrU9wvWzUIa9ML+5O3nE+jmXM8uv/1wkWFUYhl0
O6lnPJ9rR5mdG+zpwhQ5LjGAI81F+ngB4aM6ps+KiyucjDlbD/1/H49BmEDm5+qVDJJXIEj0smJ0
hND072IjrrQx5/S4esKhLkmm5AARBGQJ4asNu9RSwvw7zVDTUxyhcVcVBK0hTp4YyPxl5z5CrIXu
EUScxkEWDyt91x6+jGDpAQB3xkrJN7nchljTwkXRNsB1+BEfPWee7D59eHzlRWC+VUnB0fQAj2n4
lVxWD756m/H84GqEcwqlhF1Mo1fg68PmIvYSnxASuFJpfu1PMxwkk/7jm8BABu4Uqs3kDWv5lyZY
x+YIA/7nXUk1HeVNHJVeSdmq9VPCM0OULDQq+8JFYXVLDuu1tUIjQIFhWxknX8FecDxeZlbJrkIp
EoAMU6FH/zxS8IClolqO4Qmv0nmSiuDvK3D4MgXPSbnRH7e0i7Ac7Siz5dsyRTIRvprs7nYwzlf+
w2GU3d+BLfEmFgJxkn5yAektV5tvBzFE8uugosutL/hfnBk/ACQbpTXstzFRn+qLN99Hgfpob/bj
dIFQNgIQRLK1FK0MD6g7qAcsdUEeKDh8fX1cLch/ymjusugs6qMysRkdma/M2ROtLnKz3E+iKHmE
NOkXn7QRFbR3DOwwwHuA8NhwzXKmw9AlE4WMzYyZiwyfenN7fdbK6liO0Rlp4VZoPItNYzGzV0gm
Wy9yIc9NVGVsYjRg0yUxZArWf86EDXm4TGTShtZqQdRVbc6+YcU3UzEtwGrXFeXUfWE9g9uB5qH+
iph7cJ9uzbNJWazvAZwzE3D2ZbARW+UX5Nd+Z5LHVhTW5Ghjcl9cDla7RwUU/JOiftyYefOf0MEY
vJVOhgSdkYE96Q6x42Qy7XBytSeiCf12J0RqWE0FMwd2vwJqPKcaYaFhXVlSc7IM4iTJPHCoglyD
sBhSgh2cMqrlXIvnO4AQYEKePBJs6BnxHIif59ayWN/+Hjj8jKrr4SRY1vn8ZXirsCS7TsiyoZMh
8pTG6hVqe70kjZm8h0F+b+BB1rJkxvUyBjeA3XFLPj3b0NUuurFhuV2xtpw65aj5FO+d2ZziVmD8
dMfklhEVDy/DOlRa3X3WzMw3pPy8p94aEd6chP14O5YZEivIuwTIPYVRdk43z6J0ACT9KmcRGMNl
TiMjj3XttgYyGUL+talbZoGQ7ZHJp4X5/KbsQl7ZBZv/nAseHLX5d6Ndg47yiUWxy+2op60e/oWK
e/+umoSD5aXIE0Mxh9j9UbHnV1e/530UZptUb8qsr508DVwZV37o3Iw8PMxyroPZqu2OShhCALc/
wWpIB3nYlwTqOtLhB2UOwedkWpNJ8LitrZRJNDZqy5gGs1fzhvKpiMM8ubm0GDRSCYmzcY/2auRZ
gJUP9JEr7KHERzbemqnSr5m4yueGZlQOjfBSyhUGBTyMWP5GGaRMdYJ6p9LG9msNLKJXB9vxGaPJ
dhPQiG2TDSk/FFqbiFEhZ5IrZgTYtN3WaS/L1R5nceT48s9pUxJIZ6j9WcRoQr0bUwjU4a68rXwE
lfI3NGcKdG3uKJZsd6sFZOW5w3c6wxM6GGb6kQyDJU+t8tJYYKA0eYXNh8LGQww5PVsmGMFX83sz
3hXj5rFLC5gumZKCOcOTsOzy/Tu++ip7On3EyLI7bCkApWlorxKX2dsvudPNR9jD6c/uDoyiXU8r
fR1j5w2Pl3Kr0VuItYqBscbF15/qJSsv2ibOz2Eijopoa0IjhdB51neFOzoCEH/Aqij5HxqWZslL
+pwsF8n+XxUOmwvs+uDQGQdQURvFnY2BLLOFBVcZqAFI/hAlOZi2TlkUpjBtFgIt3LgH4SAKFVZB
BHONYlVFujTnH7tteG2e8do1TDtmrSBcfLhlDXeE2ciR7JID2jen1zIK4+BMn0ij+/rAmc+HArrT
fG2VaMTQY6pqDBeW/znuRr2CR9JVSfUZpKDqoitc9r8s8bZ/0Mc/DpAtYljlJ7GCYanmkp01lMnF
K7l7EsG5kfMup4WK3pixadegqXO7aAg/I56e92t/AgQGKJQ+4JP1CQkGquAqmkQwHzBAmOXuIHk8
+28v+aHaDCdsXdDW96lkzqosGz2BsoUUaazsN7TbWT4A12f3X8xlZ4kybx/bfmkzIfoE7T2H82wy
d6wQqrNrfpTsrQ+Iag6xpnST8zz1WjV6pdKSe+0Rao4ylRM+uI14CnySAKkZDDhJ0HZcV8WQA+sn
tzGLd8rCog7ig2oifPoLjxC8p482fasH7YeE2qwypNgtlKxHxFQCw1UjOQvj0ArNx8RIPXEauMOX
ozwMGVGBFhC+n6kst5/nWl2xa6a/opZJ7mJ6igGzFG680fWnj6cLNIrF7o3ZkaiwXo/6dDbEaFhy
qsQmNnDoFoYQ2Wtio3nix5G//B+QM0ZgKu2iC+6h5uAm6FSrvk1d3kUoDPO11Sw4eDm91bcfvmP4
W7rUpNsB2utdA4xmHaNbilLNu3A3PkLnjmYIzOt3WGB/QVhYM+pCKtVOQptkif4jmzCmehy4mS9m
hL+2ZPePhlVifhjLmooWG/bdbUkzuMQfFd9tCTdTdkrINp1oCworYH23MH9npopvz+YYjPk0juyA
NXLCiEfYJ38ly8CJJpWG8TjvSwkXEaOOmyLu+KPMTlV3re3hZZ/WvaVtqtt5zg0YkpeoRBrQoioa
W331uCws1QgtwkEKMuF855PuaG/nvfof9ls8BrkDS7ktvoJvpaOqScNJpWMOmOQidrpLWmIbw12i
ZcunmZlQ05E0mJT8TBJ7o9Je2igCdsZueJOVpo/CODpX+g7mORAOYbOTOuyi4MhFdVZYOhxqijku
N8rpZ17MPB1/y7XsX4zzbyoJ3d4RYBBGvV0Z3XSlotKfM5V9Wgfvka20KiauSNGWIuVAwqoJ23pe
626Vjwc20G/eX4GXD5HR4H8ESSZRSIMbwGuiO6zNB4ZRuL21/DFGfge5gkUFzMfbWr8AwihmKVWc
elEs+qH7jYNWN0oe/XUnSB5/mJGZU69Q3fmpP/d1MyX1i2T3TBCR6k/9Or6WH/SN8MoujFkp3dWQ
6Bwp6E5l6r5/nmodxqc/nlxPkdJWa6R57GoNceks2lSIV88yRiKrPm1g75q878zWog+D6BdP6+TN
u556jr59yjpjR9BJY2xOw50ugt3D/anqn2Ks6cDzFh80Dt+dphBgwN2+ibr5zoH7K3MhLETkbC01
6+HCPgLJ3t97HjqrqZkbVjGyXD1ORww+c6BmZnWIhbRWcpxIb+j5wFkvC77Lh7ArlCrJ0MQK4XS9
m9MYJg0ErfqIUDr/mV2yCTwLt1pXDAHJZZeMEYrlbCJVOYrfvF10JLa2mONwTtX6sXFyb+1IVTSx
OUJ18bQVBACnff0rdRzH8cyMSvPnkRvOht0tqDWTrbBU+CMeBn/WTt7Tml0f5Fd+8hffv4W4mg5M
8wAUXUc5xkqxamSUSdfHS2Ma3SwnQTNxgvpOwAtM2HpEw+VaV61R5jb19ZyupKof7yjq/G6MYRjj
2RwgeMC+Ptt3ipPNGpxm4094rpS2ijjUhbYgzrs92Yqys7n4/Oufkcxk8k/Db6M8gWQTi6ru4kz1
lsy1EC4iOmt2e+qWycP6/XkbKFvtg+/l1aRGmsRQghM+Sdn8PnRbWt9ZYKR/i2IWAejI7gmFqxTm
doK7rFNKd7ATo+2tMX8WTzhO2TYrGCp9StS6ncX+GXq8e82Oo5QbMSgSwM3J8L5MaChDD5zRdsLF
p8ZR1pBlIYJGs8eReKRpErAzCK0igsEANRwjAXcIDWxhw1OmVs08X2GJfua85ur5D8OVkczrga60
gQ91/it4PVTggQTGF3EIOA6syhVnIecqP9/KnB8u3FUTUMigTtLgVcvcjzo8aEt1Kfj1a8jN+fmf
0ofhB3un3C6T8KW8CjT7R0eV72y8bEocjB0prvPZQxkNKbQIpzG6c7V7NTpiB7jWLF3hA22dSVNa
7+bUnxVqv5NS/7TdlvoO6AOCQDXt9otYHObjBOqCewYMd6CYBtOL5+VQWMjupgkbWnLcko8F+aIB
SGNlOEGynav/sJfg33J6+NdkYueYYy/9i8vzv2tdwrimwWlF+pfmuKP33dKyQB2d0MICRjYAiR/7
jpDkMuW54pF3pfAjFoHIzf7g5n52DoBmNdMMKSqNnKZzt0V22qH1uxCEkWEFOzMGb0mW8t7SBV+W
2qOJbSzSycm9M/tDAQOz3VPIRwrs3MuJ1c1jH9U7Z6hADUArdiN37vqXwTfiWXjuGWr7aTUlrXl3
eWWKOjjY4t8dhCyc+ZkXTLQ25vsoTQsrPKxhmoRzJnkMX2k7HPRqZ3VlQKyCHai6wZ85/z8wTLnw
GeHwGHZA+TqGfmhRyg/CI9QJenkNImqSwQSfr3zbxqU0eM2X2DMkO70wFYTih57PiTJ7pKngvuvg
AozLhmRRnx1Al6x+n3YZj2lyZRXcrnGYIH99HHPaNE5f+IwjHOFndEv8VHlC1jqUZL3ByPOec9c2
2bKLfh3LVF9gpmA9NGHm2T0O3Wh2v1BU1OSC30taIzACQe9Sfmpxkjzd8bDfSL6ewefAsm/dvn7M
JT8a5ag/6lvoVJCEjysKvuh4dkd349LahPZVmOmbhVN66rqlar7htsQgvIYM1LwH7/nbQxQON1wf
U6gsRlV9UoWoaBw5+FDAUv5zOLirxrlQxslbDM+TDrO6gAbrHWNBBRssXU93YrKkjtsT1f9+oyvh
B5MMZWknpGXsuhz31qT3J4Q8Lo7wvPC6dXFd0go8NLCg8TusAIFDdiyaAR75HO1raZwwooN+jxBv
u3uVFcKtwuLToPjk94aM505euNP8xYJSCTmkJL1G2zKFoerD2tutMZIog4DRqw2IRYHvN26mvL6i
SDOSXm6JkpMTX0OZoZK6S9IPNXhV689qRm49mPpY0zX/K/aI5UOm7616JbmMt0LV0K7H6tiFXFiu
1dnY/Nl4SycBlgiBmr2cyFObkhLsurnqWlLKXZ28kxSd0iT8+9wfID3PhZVeexs9MBxJ9/NzWmBB
p23+GEd0PCZyq44+cW4UxyONPiZSrmRQixW8Z2rC6bFEWblRt78roAhJvRgeLEp0s23onbAAQcIk
vmeZMyxDL0aFsjlJHCFBniMyd1c/FdoUfoXSFmMVWmuNeNIu11x63fdzyWJGVbaE8TaEo2yZxl9k
BfUy0h71WuC6HqqjKI/+Yn6bXlRodQrZmWFsUnBeGdrHqjU9BzWCsu8dghVSZ/KLeBr6dLXTGfZT
TrRffoyWFY2UHMJOd95agPo9GVm+Q8lLImMki8XK7kdO+/XaMtZWmRuiQv4wer4gpx0UEOizuPaD
2fL7aL/XPYzVPnOC1x7jemW7KNX0IxbDq7fmC33iuCXvjBEA86WQnDpn63WMMRPVl4/XVh69eb1k
C66/jvTpg1B8vWsI6itOY8eiEuJSAer3bT5N7oB2s8wYiEAYHTMHgQ6b7cDsrzOk7v03MuEBgmwD
r5DVgiEZlNJtXEPwnNRZMbAk+TaIW1uhrBtJkbIPQI34PymJuiPqj3QDZqrlps5Wg95T+1P6zYAe
3uqvAyxmfe57yf7fg7tDi/UK9vn3fopkLxrspRN9uEbEfzqqIE0GeuHQKa6t1RtdyFfH40qZKqos
sMManuZZpiVntv1an5O7AIQRNMEI2QpDGM2TLEZdyRiC6Jqy8xnrPWbwL8Aq6gunGjQWDBrPGW5J
WO+okdnsRIWpur7bCEaRHdVc6yP/8ncKjFoRh0QBmUM0dilj68Enz1krkSsbgVz8+oah6+cFUVtV
EdD5uLnBNCoGAlwSg2FZmGs+E4SqXbF7wJVIr5cR/P4iqYjbEn+fqJt5dUuTzh3nuFf4aWhZfg8a
USg0SbqWQXI/BwwG9zkNZF6Ewn6+DN8231E112SuVx7gJ91gQMxYKJal6S72ClqTYK5ihprQeIJ0
45SliVzvVdAQj0T5PImtOOGKdKh38kyVuDfzUAskS/1ZEgrhY4C3LLCQawbnFzv/EllHQE99AeY8
7CiRg9TabEyfZ9mC3oMW6gDcTTypytBuOK6uSmuyOYqYCTzoGe3EvaAbaHVLoLM1N0ySjXVLIzQO
hD0nlNQ9SM21GG1DsBTxlAmOXB+Cz8FmM6Po5213ycgmARJH+KlFhSyoxX475uw9fNkFds/pFHRl
Q8Js4OBfdilcm01g1Mlx+qhEX0c4T8cqqLZky2ywrv+JkPGfjsbDGyFI0/4kgq94QF85nUxGqBm2
9p3nfbr78MHeSZodb0AG/LSR2Z/pa5DV2nnXjjwyWUZTuhPh1e5D7adYfs9vRTcaAN2mNhlcrvdJ
Zu0mR3Mf1kx1TI5aPP4v+/5Ff1GWvIhwWPsW4S2HpppuJ45TThpg/MrUI63TCrd1A1Bv+q4pClGr
5o5VecczM9dKKVxJtx1NfI59eMaWsKtDwXVpUYeu68msovsDCvyb6M1IJId1ASsrGVw6P8C88NSA
qqOJbbG5oRJdPOJ5QL2BdvbrfiISirBwiH5EIHi2JugL4RiQXf/XJa4Rf8YJG22afbpBrBbKMH19
4cP6gx1ntUR3sqzg0ARrY8diAAVPiFhqQkpxhzHxtUBFr5PMBb88r3Xko6ZsUilCIbzn0spikxaH
VdzC+uzBPT+PT2oEN/KSw7oryysHIllyMltCO8NU34zKFn/nknlWBLSU9LmnLaYADq4t14ouVBlD
ORCpRiixnER6FTc9bIu+qki9BJlWE+a0n3bHBu9oojYiTdYovAej+TmEO+Gvp6vhPoCDLL95BMeD
LtbVih3747DAvDTdCyYqvBaFqb7HOeEwuOLSzmwevzF8XrNpC+XPm1fJqWSPBX/cJrzxv2qumNc8
yhRYL6+iiBnVVJrP1PfybEQELkws1HLRPHuTzVohKeG3kT8McUnaYlpFqEAYvKPfORGPvKFX+5U2
pmTzExLiHwMjiGIMvSltoxolYoAubJCUMMmUxlQmNq3m7MtL0p9du5y8rUJwb1kLwuXUUAV8qQpe
iqrH0prVQY75IRACC+AlaamG96b2pNSuMWwkmiRKMmxVemkaR0ik3zEgN1Iwke7vZZxP8Khlhlmt
0z5lp45hBrix+Jmf9GVwuwjDYvwt49wUVIfVp2QSlPF4Hl070JHk9Z9/cGWxGLXHthpYAThkwhEL
T/181vOlXNh9zyQzvO8c1TRvyFd4CLfc6ZxV6RADQmOegsULuqp+jbgY/6UdDuIDMXl+R1oQYUpC
rHlF/n2hvqBU1wKgUkIvHwtD43jshHY1bt2eM/tq5Wj/+DAbH+BjpkX8avqqtCP3rrOQOY94BBiZ
me71CCHVLPs2N0yDeN1PSU/zGkXRPM+8p2QQ1y14ODJQvD6NWgQVfsDO8UJkwStCmjVWfAM0H2IJ
VqQwJUK05DCW5551iRlKpByusdcbU+i7LPNkYng5opjt+8pP9hipO1a7J1PKtzjnWP5JpnZ2B0O7
qGDkdzpJ2ShNxsV6TqIgd0vGvElcqzN6byXIzsON714ygreaeeHJcRC1UDo1qdd1HRxKc2krAUtC
27uuJRu5uJphVc8F5YMgF3yW+3TMRbG7FYn3clux+gdx3AiW5LKrTNxHULy8Nx+NY6NCfhvczy/g
f0+XiPrb74kjMRSYNQOKBDxVsPnid0bih1WLYkaUZhpkI4Sejpy6XHQ6ICQxv2RWvjMyU60gLndV
ckCNKiEdAp4vHo/mNd3BLyijNJfgIidVYA44EDvS5ETR61SUde95B7d+pbOzRWoAWaQSPVALShxd
I66qQLSUdJ5bnJA6wqLg/R+Ohrk45ob9StPa7sVKpb7cJJYKkccjSaJtSZ/jIPxahkQdkogecjMB
EgsC4D6//F7M/IQF+b3I4g8zSGh+SIlJDoaSPThejXZHCF0cdBv+RLrjXHapyXJzyK6kmFtzJiPB
Ezwg4FSmGhNPOPeHD3ITQXEjrCpSHjMkdbxfVAqGqJpLdZvGcDJqBa64lf435+OgbN9HvN7CiewT
c1YTQIZSdGjedHBQzYgkTOGLc49aTqn/fucEWLEvopVwh2DCd8rwW2lCYEJI6iIEqP6Sn5Zseonh
lRp5HzYEaPZ0lSad49aD8g9URlHAdlasUk90sKUhypiJHtXAd1+JMV2dEr8I7qJfclZ27WVzU3T0
BfC5OVHxSIHM4GHUkojkhi6B+PpGvMH4yhPMovOs/yLIUDyVa2yzm3liwQ8NbV9jSQvcU89zquN5
wRE2QwG3ReZrJk0qukpv1kpwbjWY9TykA8bRZ9isJz66Pk6iEZDog0y97zjEEI3amfqgrtXU97nJ
bLRKALTTK9qthfbMsRV9GUna1AIiVAs0VZcylnf/LJGEgLUqaslcqo7s8cno/5cgT0fhWE9pHWDY
tB7YLfSV9JKhizRTy2HOCRvRIdJcaXzl/nQjlfiO1ulKprNMeZyCBlcTT7FaQoGvewvbUSP6jdjD
ZVbRgfJHLasJ1c+x2tXRRv9+eBZg8woAvsqtxO3eGd0hIg6Tgzr+FFMI9JTTVKUlXllgHf9zMtIx
PEY6TxvcfTYvKowp1AWeJZ4EIbPEXFKNw0lv7NTfZrthLT0ptE+oLCQdP2QGTDre95u9BlRzNw8w
LcSJHEJ2WBS5LyTGB8ReiErdjc7g5n9gKxQ8WXmoseSV7evk8pWNqu5fwO1HXg2YTIDijzBPmBuE
NfbMyIq24AK+Hop1ay2O/swBhz9wH6Wge50f6KJIvNgsSMZsPHJpKqSfhijXIgz9hbT5Ne1qCtxW
x20zgfi9iQivYyqaJjKmTcvrOeQhRFmS4p49hRZhQpgRfm0CXEpG2/rrxWb16rMcF2G65/FQWnfL
T/jVo4PyRrwnzVSrlkfeXWBxVxsqah5zzS44hGySdYR0Ew6YQaIJiyvqkITAq5lIQ6nzDff7f8QC
avUbveuZ+3SLKLre4sYTE+5NQRncaEbHavq00/GLXSLiBovyk3Af/PyhLb0fKUABif29AHYPzpJp
aHN2It2GoyG3pAb3rUPlRqEpQVK2wHasf3f0v3AuOOu0gErCYfPsTvv4b8aRF91fO0IxRqSQR2S/
iNuM0ISQFpJaQQiXp5VA99xcfn8BpJK4GcwuIvrJi5L7gCkXFQyl/TfbPPnmzWTJyI6PJHbMOaNq
XCI4voWjFwBEQ3HnoMbR9Ur5lg5idVJkKdOeaZpba0CHNMbjjqJq49sZQCnFXsXFJs3QMls1YB3W
8Y8arpq+84kaynD4e9CrtZsJXoh6FCcdl62QeMPtrI8nGTlCGJamiu2RQlpE6rv6fK1yuvQwuqJY
fugnPJf5y8Oga6+lgvv3zQgSbMvm1s3aC09e5iG53cuOjNxhi5JB8bMZji6c3XBZtuRIIe6+4Pw9
8P/Yr0O7dsv5FjWCK0V3eL35QKbRt8FdvmLXmeKqO9zfzMk6sHRvCJkISqWOozFcuSiCFLxFwl1P
M07EZriskruffbV8SkAG09hB1oJQpLFGht4+GgY2BRAM3bqV8p/l6Lm8DTrat03A20Umsd80vTnR
n6cjJzpwjWF//6F5S7HvFZv3/idAAeZhUsOF26/c9/UAOn42cBSwiudpW6a2x5sLtUXHSMw6CjHa
KMvvRzktv4sxYecmwvwTiImVPM/wdX9r8M13/4lnGvWeE7nnq68AJuAchvtYOgzHC7UeQzUx36Bq
D3ouihn5iaPA6dhT+Hxg7tyMZ+kwQs/ylL7H0qw0gJDXKDg4eRFx3ONJAxcGwwyVKbZyXcapyBbK
TMMeB10Yr7gTkMWpwiNr2OpwYHUCXO17+zSUfGkQMFBzQAT4rNDuLuypeZAPpYLeBdgjye/QkdKT
EMDGlO7l+/JCpui8NAZNQZmp+VxvTOTfWyKD4rGoYuo4RVyrplntDI8cu1I1Y54Hu1u8ZC8OCy9L
sLUKNMQIj7tpVbmrZBtBY6D3NHBWLejj5JaW7ACNl8hlptKYPTtPquLgpPB2ABNKI+KIqpnnpvnG
sFVkSstyIR+99vT8B6H7P5cAniZTb/zM8ECE6AxPtBewwJoQXkMt9NuoGDAkZmYXjofduzspEgCl
wBxayvMKEiLuYAFiwZIL/XaAXpLlEUTop8I6Y21AWrsEDI2p7fJcTT5ZYmZkM9HbUW9woWEwRey+
HseXSqLq5Gi6b6IAdH65WhSTT4YZ4YjzkNz6lDh1srLcQ4SV+LA3g35J5pUBmtGW7jAUja5ldxjc
Ki7RdPjMX01FFUDCxWSjsTolmA59/X3xcpRhRELAdswbkpd/P5HdUftbamT2Ptal/00e3Py+0hsT
I6ELZYDP9949dUGcWzZElaMA+4dVXUsoPctG81MhUbJ+koxiySB2gUZwlVrIWhM7LqwRPbgybVkF
HXESSM41dgwijjudJC2XH7t7DEa8hV0T4yYN9k91cM8KGrXF7OWgNMdOMUpdKSaVziK4A1fGdgXL
4RwquXNcP8kKJ6WAMn4tBdTBVbC5PU+fWIn9bfPyBGpN1A7JuyTqF0SLg2zbkY3kT4UrhEWjB8oN
YvxAM0ekMsryGJ7KGM5nkh8UO8ZK6w9F3mq9emoE2uTJ/7rO71KkYfcqTAKj9Y5pMv+GjNZkQKA1
nDYGlh69IsDgubJZwvmsTa+v6RdvWUsYG4ITEBLaQzFTKRW90Kv2feG5jhebNB2PO8/EaJnV6J0d
XsuUA8IyK+2hTFCFmCkEnCso/eotICxGGTSzMUsZlXupoXkp8xvkq+Oj9P/xNNjaLN2fbJYcvL9J
fy5SuTetMEDtgUNCSeP78i1V2saHCgaDaO6ssndIwEZNhmJ1oXBWBOB4EVlEvb7r5m58CeSdcx8w
2zBFTN+xaY0TwO6uNMYaAHQCvIjRpE8jdrA3ktKCFanYMMb+3xS6AR46777Ny1agw7jfKtwmWE2l
ktzkmTOQF4AnHqHOPyFZf3LInyp3Qwmxsd10C525o+mf5yTWdZx6sjk3lCsTZEVp1OyUAMweFzeU
CYLK/LBtwQS7pSDtXvXUrwE0QjuTdu/4D1IRVfxKxBaxDcgL37oRk3JF3xhWcpfBn0RXll7KpjH6
fGnOscYc6UHbKY5wCAMS18WJoxkLS3eGYdI3wCbkQ7K69VpBrACW6aMBvPYxTDE62SdAcbSjD3pW
SQjKEPDwLaY/jvmQgUeED9TEGiMgeJF6URclGKnmZ4VZtIwjRK3dVbltmlaefp0ni7HpaTLbFmU/
O3wWaqEppzpO/I8czb2cduBAfgQDN41tfNWsxLzHNyBNBjSAQ1oznNQwoNRC9eJtNIruSFzF6u/b
CQ0Twb+KCc3DQ6Fkos0csSg4W3/dESdSqoCugH+s/1XUqoElhIdOqw9mZporGkty+IQdUH/BmNaY
hKZddkLalJ4Ch08U+9uqIt0XK6VNhDyO3rbakfBYcp1JVJI4o+YMDRaFZtTABk9abZWDxh/kCAy4
Fu50xIO6Vmsb7qRYUQQBPGavMEEKMHmK32qIjIAzxXaX3x3ZaHO2JYQQ+/RInJTpruYgaJx7O4rs
7SNM/h6twuEs0jBduMEOTm38KT46ut4Yxz4Rd7QhEOT2O3OrZMLGuk4FMcIwf4ezkj4i9IGQKrU/
FnxABDbTCphEO7aKgZ+RFFN3a/W8QBxOgA7W8csokDh/mGCbrY2g4PR5dX7IroZt3CqrdREv6Vey
uJvWpUddU/r/lljoiSToAPZgGmnf1Gz9K8a+aGp8G4WieBX+7M3SfNRI0WTaSIh5BbhKs9IK1yu9
/8lNzcs2r8zcZ9m8RppATnlLq9JE3G4Lb0dJDrCJIV0ves/xzO5wD2+liNLW9L8mjfbzQtmLIVAf
jAsZZKdvyEqRmZ6FvO90igYEnOoABxICYiqmRdKmYqwa0dDsK8hPOmMDEuoAwP+8xLkvxM9vshum
81s1UexDi31ufGR2grVE7BhaSzT2P9Fqe5E7mVreX3C0RDK8+onfHX3U0ErZgReW2lYf6XYV2RiG
Wqei7kNtxmdy1ZJRRxtZV3VOqFsWGsjUV2FvJtgnB6R5xbEJbbd/xdxPUX093p3AHsj2kBRuXqeH
f/O9Q+aoBiHYGuQrATSS6ScSOfYu3efVObdY5uSjca8Uz6452Jix7BJViOs1RMCD15geBhuAZ725
xrjasTWmrMd/oDoCmT1pKZsaUt/jwn/6wTTm9RpodVRnAP4RuLqPDIhupuBEWYKdmJsJSO3Ctm/9
NwX4VTzTHrHvmgCw6G82NVMjXYOcBb03/KQT7xNHSGJqkQAaiVuhV6n5ETsNfMpQIrlVlzw5Nrwm
LatXawUo90PZvXhuxX069yKy1K5zm9xp6pnw2gh5yKlENI8WhbybdiaNpyc9YlpFGXAPLLZPmG/U
Z9atxtParymyYh3I5DwyHWDIyMWvlitmB5RByZvbQxsddO5kOtjnMNnPUYoIe9uGqLnLFx1GiEoE
d4hGCZOZvAfStCTZ5FvTairrAYcC1v89cuhIQSEwURyDEyoxZ5FFm863OZNQ9BtW7l3CKMMkL6I9
KvFqZ0b9K+LWl+e2Zk6XuzNYsOJv8JRToVpQ3oGut+aIIbHLij2nru/vA7RVjF/DBrh/R80XD9UV
NorYENTCNVXjFjWSykjnNCgtEpNUfDfzPEl23wF5BxGU+VO22TN0Ny4kKDIQJQJDeNns90UxXqiv
Fel/nlREJIFkrc9oGfMWsEwK00/qb3RY0WE1OTNGXzt/RhtNS6oic+6DEhRcgSfCPBufl+kmLqNE
ExtTqDpbavcb6tkr1ZKSehuYrED7riDsQdo8ApoOKR9LUXJnA8OcDOQQ9fuatjIHOrr2U/WxhNBT
Zmz26Fi55KZpXhyldGh5aAjFs+L46VYsZlp4BwSRxcgWYOHpDUND/ouJGfmStfRi5dn7193dj3NE
s5GO2ojo8Pv2MfE0TvyYjlBT4R6pVPCGybWHGisnpvNEdSxRPiS+05xAlnX+34pG/qV3QPCF2yAl
Sm/RbOLPVl1f/5pV93IgdO9KcEqaKFymUcaW+2oeLMPXs2++rJUfK2Wyjtjin6VQw2dixNq8+pGx
b9/k82wBhmulSLU5g2L+E+sZ9LYlyBtaT4C9Y50AnWSwp+ysD2IsI/7pFJDdyVFheZ8GgSYwLCXJ
sQyEQ8LWZk+9kbxBGe+OHGiJBnNtnnKJj4koxEl5IdKI3LIW8f0LbOR9b3gK8uSv4nCYJQ0Kx9p0
NM2VaC6trl7qCIesQ+mSzS7EfpSLeESEFC79UAomeGqp3fRGW19fgfvml6uOtdyK85MG77PZwz2V
wc6YM5vV9Lbjgm3NsCWjQbs+JbXhZqbF+CgrYwS0yVfamSYtBT6W+9QjQkBrZdguBPbjaBYNiwuc
/SOueVyPyF4OgUF+JVyMw/0TO27FnIVbCv8efJQ5OIy5PSissFF6fD7M0MRUfSqo2a/F989YBQY9
NjTmnj15t26wcmzrAqSth5aRSIuCAfhZHmT9uAQEUgAJIa1+HyHhF9dBrDIxhXmHeKvJbY6zQN9k
/AuUFI7trTefrGYC9O3xh0PxKjQFlhMMY2vBt4nKtiwriX0KNODkHOmcV73ByB+QzOrAjHH84q90
K6Tm4Dl5DlIlsaNdgvspZwJ/je+icgnUtbosGbY75l2kwDe+u0kbNNt+ln1SE4McHXs9i0p43WNv
xeglfaUKkkYJ1LUwxLt+l97INBP+df/dQ97SeR/dAtgNG9lCiq2gHsapL0EezpW1QEmKNsojtvHa
kH1S/fd/ozlcRhk7gKNoqKGAwv4uQUjADBNOgkI2nJQKeUUFHaWTb51LlJmpVqYiyHLkOUy82Qch
u2rbM3qzYU2uTzyToFVxlMDsC96zOemMDqAUa1FzPib0MsrwP+mZGTX+mzQtwkT/jnSTxTHK4DEV
esNaoQD1XdBxoKWbdp5Q1FvdGaXveb3G1IjksAFN57a/H1pBZCXSI511rrOE5W3PTeL9fNlJ56SN
Mdj+TRQrkUuq6+Zq52zcINiDzKBVwbhBMU75d+byxt6w2JtBkWyZrRl7OxLndC/5wppzx1nA6B3J
NSmUlCL0FykiZxoEbIOUAfjy16iPQDYSKtkEuG235K8lu38ljbXE2Q5CZ0RNBsV7kBJV+bqN++42
el6MY+JnrRGUTfmXB4+I997fhT9LVCWIKNJ7WXAI1wNLcBftwe9HC7yp+p/y9lsSnUpnolW5ZmSb
Fp+Z3Fkv8YZpznk10whrCkKTqYGLWFTmCb0s+ALikwZX/w1VQLbdAEhxS8fTNAkYULjlIsEvdzwn
tSW0r0V1Ki60g3E9jJwlMyEh+tgtVEgmwqGNqBwCIlhqKpP7veGe+2WXbSvi+SzJtW00auiDkNRz
bDlsBVhBFeHHHanKh2VrAKrndcFvUFH5AbyvhoioCysXjM3AdNa3n+BxCQKpmmUbO0eQolPagVCH
17HNf/Anm8aRWh3HYXhEzDWYL6ptl0VSnNtI8ScmXV3dIF/65f4w09SXZAFHAsBaJOOqB8e9I/zW
6AFvt+EpZ2IMDSzwiOCSlQ8f89e1+WzSxWY0dETes9GRyBTgmBA+ZxJ4F1JW82qyHo1YN6SStyws
snnAnp69idUEPOcXlAtJ7WqSxeGrorZGu7MsvZfEtUrpAD4Lm4duiwfFLFvyB2vTLuk0871mxbdU
hZhJr5PKUQzsUwKMateTheH4R54h3TAu5HRzXyKhvWVmGhGAQfI5viNMN0RWB+vLnv0GxBTN+od4
xzKFJhKC/fN+HBDcdxoXVaeIlriWXfOTtgl4vUhtlbJvOr00sVwI9FfGsBxti9jjbgzrSBLUwDWu
J43KiKX83+3p0J+HBjCipmK7Uvz1eVsQt5QVjL3UUKkkzaQlfQJfsJD0amVuztqTa1VcmBynGZBK
BPMG3NvjoKPUBUAW9NFxJbkgE+EXLnvYWFoDpbS4TOMWsPHjr8qFV/efTG3ZA7YfInQjEOxNbAX1
EKD/FyDUJP25DZjIGgjL8mddCHtrlIwnnU7E/LGpDrKYSF2pGFXsOpcRRdTFcBcf8k1NqcHgtVrR
zPM8epi2cjhDitat4nXlQIcR6RF8tO2R2z44pjCqtOa/qFJVPT5TwGA21RBH4oZ4WWy/azw2wKGK
HFLPrTo1Hv69pW83Hs9I6vf4z1xvYYjW3yM2yf39PjrQO+ilfbWtPBmfL4wwC7l7T7Dr80ftErhi
w5jni0wmkMa5vT/EzzKJscfik33ifb3nKSAgkSKOIDpGYgYrLc6IL67iOSfVISzfIU7T3KplJq39
5sRoLVpDFuSmQH/yBBqW0m6ikjcRjz+bso9LDR/f/OnVstkDHkX6XZOwAfJD6uJ7Xezy3kiGMJzo
9ZEi3EFwOS5wXPimtKyt08kvgd2kcbLh+5q+GVE2uU4N++AsH8y38a84Ue2r1cwfFks4oP5ismd3
RRi5BEcSDGbD0Kw68ii3ZMrM8Z1B+oZJLBc1+hj4sb/V/VOSZV8mapJezVv5h+YPrLoD8FrzUEng
MCegDzA77vk3XER9S1xIHlJ6dSYctjM5b8vvX5zUQ3RTPr8YNgSMxsG1Qpaim+rIhpasX4KlySPM
yDiO80wxObJI7KBTTqysZoed8nORa0vT0G3TVKOZrRDTvg0gRezi6D14DdrCnKTn6sVJ96s4/E0K
tLfMDvh7fBGfGlERAhrskfT+nANP3vc+tgWbMuKeZNMP9DFh08NzOGdeeD38URdloKLDIDITB4Wg
6fJDElLZ2BRgLn8ELqgKkPscjmAV8cr3kG94aRkfrwgO/bg1Y3NkVfmLCI7JC5qMvJ2mvnOlrDGt
rATGS1eNbStGYGG60CsRnNJZLNlknqSQcsZ3PJKICZShJHtiQqEwO/K+Kb+C0UpDusqvU+fOY5Cj
7BYtw/iePaitkWcW3VHvRmsgRVX0UD4K4mxndflEVZO6Kz03mCOEVs2KpIu9KMyKtBPwHxyGr/EC
a1I9gcE8lfL8N8UTk/PK7hXAEr0IfJEp/a2keV4jSDM2JE/MrLr+iYu+7INyHTiuNtySdD6K3qWU
N12lJwWgIMMY9QHcFq3Rdr9x/n+saDULmeWjwwYdNW2S01wdOwKj/iBpD1YOHupKqrjVygUjObyr
RNkeIzKG9AQmuaI6ZKtTQ9hayixuhhAmHxD8S/SsVHQXqHT/jisgsbiTJCzNRYVrc7tEbBqSqf1i
kfqvJF2HGLUnhiXeZmmBM1UBXVFz0JExt0R8ewVezpmOs5xc4DkUO+AjbTGQ4wdlciwm/FXdbipk
y3LpNg8xCBG1SEkKAWvtNErNVwh1GFxvvO4q0HCd6XU9Vl18dBDwFYxFhBYZGAndJJm5bMXsdEBt
cOoBkT2cc2o0Dxs7wVN4Z3ImasyPZlOUTpEx4TfdreCxwt4c3+H6jwHK+EHJnRri8LbIn0spx4pd
NXOXFsEC5me0NuN2LYwMCtalb6vkEvqbPFltTEy0gEHGLLQ5Z4AUiuADy1GW99Dq/AptvpFOKCm+
BkmFtw9OijBHRL+gWZwqI1lS09mKjcE/plhBhG2CnknFqucz2qLGPHGkF2sxD/s+yD8+X3ZUVXZp
ilXgGArvUty554wo22qKdjBSLCYDFJAcvzOLkIn4GK9deuavXHWm0KTHYFeV+1UWCawNe4cc5L2O
zGi/l+v3vzLRyK6/qxOzo64inEdA3hYfphjXRB/AS4KTUDtB7XIXR0qCwPTNmKdcwtCbNCJPrknX
GNO9r+g8vTI5P2iMDI/k/mWac7aX8mGlyp/iOXAh+0pJgKOVT19LZb1vDzUb1If+pxQfYf+2LuUj
BRsDPmqIhEH3eCOkdRWgoSwS4/9UCqK0v8Upt7tPHVo119l5YBHBmlmoRslnRlqVm9bH4sicnQwY
5LC7VsmXJt9QTDFS0mxM2QEjiDwS5AXXjRyAzz+z2ckioQsMS7aPbMqZkfEfEkQzPXQAos0Mf8bD
XMKZeO17j5rffpHQlTiz/RNovOLxGg90RWQp/2jry9btrneJurwPAnokD6IuLU4tNjOO+UPdpxys
KFq8mKSxibAOQrCZoBPNTrrmrrjNsb1FvZa/9a6UrU6kUlJ7PqP27z5RnrWI7rQvgx2/JeerGKsA
JhZyO4rV3CK0jRXX8afd2I8M6DKbKNc0Lqajkv9H60c8aj0UOO80saP9zKSKwCZcA8HjW9ascTci
IPgjwIL8z3OPhfSymFRr9zCXtA/gioqvxOV24XkaBT8QGdTdPG3drm+HRGmOKaFoSnSks+tCOi05
+4LA9Sw74nx+3JeMNYtRb+DLfGvWwOydkQBa0NeIP1NYJlGfrWmN8yRIjG8YJ0Lp5yEdZGubnbMv
mCR+u4G8Cp/RWpC2o/1nSu1S6tHELjsXyp7qeQIbqO1Zkvdzusvr5W2B0yEgKDH6D0n00+Dtc1fx
pvGFyW0ZwAGM+wndXunnKw04s+JU7CEGOu4bLP+7YUrZLpkFM6M2Vd6bQ5qithel3PUMOvvTS4DG
WIpz8/x/rMXEUpVd8mEz98nZeFakXekEj+a+AWcrRLBJAE38jZjpHcOfAFLPS5G41IK/GbbEo9Il
yFYd6T+RZvxFCzIYPg3HHtIkJu2NxSuZkoIoSVPdWLWRCi5OUJzbI62RRnTadG/UFWBoVPkNCFXh
Rrqp7xrm3g8hN7RZczteSoC/rHsi3XB/+ll0ypzWDuAD479h4jrAtXOiB7kdLBgfz1iwj6Mb8gLp
3K1247at/aDj9WFgtCICAe1va9EOW62zutlB8oOKHghLd8LB4rOq8O9HJvcywdkGMU1TKlPMlLWS
hTRR/rDETfkKYKpVnns8n6XZa810oDhRyGol5bBwgP7OgsNIwgqHv9PLnWF1OLnoUMCshReeX2f5
evIV5f7bUQ7HA8jN9D4ms54TYq4m1lKzvGeg+HAny27u0rkWjDYi47pflb+0JxZiV0UaltrojFsu
TVq3l0bspBY5ZxLi1mxi9oWvlCEOREOx+g4mnHPDpqI+TIlbeyr2DYle4UGn2+s9WAeBHGdycYNk
lCtHCMRPvPhJDX80ySWGtppDvP3MdeyuMYeidoVseM7RMi7w5bzJnzHaEE+AAZ3ymvr78359mxB7
d/FqU7jQBPH/T56PgX4t0AuHOqKoMNrQ/0bPwNfbnWzjHW7916RvOGfDrtKYv7ZhHv4GgTbSkLZQ
eOtOg7AdXz1CGEFltWWg0esCncRMYRVF/FIb2LM4S1HR8nPbGD0cqUZke67Ht1eZ8oytuwT8Judu
yq2l+Sfh+81puWE/FyfbIBitGvWCyQP6cyWIj+HngGuM3f/+aGRhIiSzZhWJK77QxJkF1DjFA5Cj
V/6PYxKyiEqsQl05HrqIqJ9G7YNS0SPrhp7RgwLlfMaHE9t2ULQjHQyUY+KCaI16e0prjxVZHwNY
F+S3tk9cN1WpO5kSja9Z22NGgNtr/Fe2+CN4Pwd6/VLSh7UDN9fZJeC//8mdkAveJXvIazp5SusH
lo68Rw0KS53I1/8M6NuVjDAyZ0THdg5UcIEjswlEBZeAMdLi+3njwYjZcivkIgfbDD2NHEaeEFSI
9pLL3ljTxE2vbawJDKxWDn9iTKtu3MzTbjBZTEWFCY2ewHX5HGwuDzuQcqicTUOw21VswFOAYMUt
xnWPsw16bDyFoM7fJkgvXgBIUEn1g8gHYZ1pmE1NvguPA8M6+O8c5HNFk5fXg0EXj2HRzdPOvncX
AQ9sqGjPjnPNJsFbciARiTfoyOmUrR7IskHPZ8u18RT5F0JSFeSJuhFHPDWjwWKztBHC1+W9/MXq
imSQ6eQarJJaPaSaQycXoey/hKsBZVrnZoCFFvLr02lUgd3HHjA3B9w9TVtufeqbVl5cRhBPIxjy
uE14OP+wuWlLwU3fl0kzyT680m3lT19aY+dqSRbNe5wtLskmlk9URDBuixIGx3I7FMeOzGdrVLcW
YfZJ41alntzDkFLJ8ATdKA+UoNGR+L424GC/518dulg3NPgF/AbM7PwkpJRLTb8Hegq5Siftomo0
WHlefxNbU0YPL3mOys5Q3wNlkdrY7KVPCZvmlaK24gRg1Dd1DoAArfO9PeUQw1pjwMPCXEJqPyOX
qkd+evgNQIQAF1CNjeSulRieD6Aq71+KvvZwb0gy8K8gkuVZ+uW5FXtWOp5WBXLXW5tNdTIPgSzc
Pgbh6oiJsZPpyvL4klSDeN9LWb0lZ9FIAxbxCbElK09aDnnBxZ6G+SfrkKZ7YknAblSa2PFSooH5
oSQKsaESO/b1cOtHTW/H+DhmQgO9KthQRu+8D+NOdGH+ZZbK/fWovvQVKi/bng67JMCfqteIfFwu
UugfNuzuhmEs81xQRoGUclfo7/R6ym/fnhf+bDJNLWJ+NkLvhzj12uvuuUJB7qSABK/gBD+x1pYN
L6SAzaIbjihCdxmHTRftbc+ZIov9a9EfB0FSaD7aTxJewwYigwQLGKf22rTwX+c10NziCS0kfWEr
T54UMsWe/X+RKMeRFJejIu0O18Y8p5cnptETylxX68Jus8BDlYRCRZT0krmpaTK5M9zJ5w1igKxu
Rhx2t2lxf46NVMnkPsMdmAvpnK5OkB/f4CaK8vxIGA+5vdMD7r6icZSFKlf9TYDmH+doz/QIjckJ
+ScXijwj60LsO0woa7PiO+w5jW1PCawoxX6QmaHT6Fj+gNxj73hQg+XcnqV8NNF2Rqk/ZjFY74DI
ufjtdb3xDRSrb1Eg/EVFq/gN3Ch/F0oEDCojppktw2DW7pRjhHB3XGPp5gpJ3rzj41OFER9OM8sw
okWD3hl1w4mCZkOmQqp/6UYdWbpViQIejUKwpcq7faaqwu/BW5JQZGLdGo+C7dbRb1DCdPDfq/DW
G92/NrYzpGyWz97BwaOu+Me6BEQuVHKa8Z9zTVJqigFw8+/u6WOc7Mg4FBYb3R6x3Xt6vXpxgAtI
TPPM/us/MwW5eDQ2SNw7CqlxFQgM/Syhn2Zq5wUSQntgtyf2FvJYLp5T2qU9a2Gs+o2/5GbRuk58
DH17wRLaXpJmqYyXVkNWKGaO7fPi6CdJhiXLK0cOdvU8UZHI0ev6ODO/W5vusGykGOexcBvIH4j/
0snPp16ooEOhUnzIw0qgpBQMAI8JKjBLO58evZSo9NXN8GZV0JA2+Rw+vrfaf8vPSj/4oiNmJ0pn
snADBbpT34GWvMqDahwOSdqtR74DbBbFAY41D5tRFx70n1apbI2laoHnlYH13qQyKublF17EO5A2
WC7yFUbHuopl+b8ySuz/LjSbGJYD+iavZc5y+/DePE4vM0GTi6gnLiwj0cW/zeGc33FQITWCUnO0
ENC31tS6uXA2PfLC/e66q28JaLBNa+NptLKpc8JxAjWnu3hy7VNi49m3LzrU19F89hNQSr7lFWX6
meAl8nbfRSbpVFtawE0vTEOoAHFAjCVyQ1NNVkG1bldjr8VyjnvC9W9vorbl4ubCTIzg6NeZoBVy
h9p7I82IDcN6jBkjliT+5/FZNJ3DVlBznMWY7JGNgV4MONqkStbNdBLP5BWYpRhzu8oRT1PX0rfo
3JiALg34En8dWIDiCZSBNxv6A+IXgCy6iwdUnYUgs7iwW+b6encE9uKBsW8W8H98FzXbxcAZRCnZ
ZQpPJQQaISp/4ZzK+/AE5vM8+In2Qqjxx0CxMC4qcKFXnXbHCQ9tLG59+EM2141Q2b1K+ZG7z6/Q
qU2c297wQW6Jwf/WgKJpf2uxnQL4WFGdjFQJx3hhqvWk5YA8pvupUAqAb+o559RKsxrN7mrhoT53
zw+3apF8zeRKp9hzk9vT1lxidl2PxRm+axWDQ0h29SQITmsE6EewYsV4QCMwJ/bOrbgVCB8gIj5n
fznVFM3Nni7mJNGEJuun2PHgotyayIM1xpK3dceqMqC2ShZdX5V3pLAg/g1vejBo+dMNnLh3psEM
X/ZmCvtdPgi7iKHbeBntKZ7M1K2q1GMTuOiUG7KVCCyMeDZ2J6T3AeA3V48tbUJqzO3V/ctFQObG
2p0WmEdNEZB+7T/afoyE3PcoH6vjeNQninkWcIZ4lVZo0IY2LLVsTWbrsQ1j8SxtWg9BzjJqDAyb
1I+9dT9+1BdEObeGWimsEJn1mr3WdOILMJixGS45JckFKK+T91RrE6bjqw0g4d4SID7S+1UAqKGZ
VCVKW47ULoC5I/IQ06l/zcbq8v8CDMKk8WtYhLh5vXLeSWRlnfryTuRGkCRgGKomVXuFTQtBPP3T
Va6/aFzB+/kKoUlfUqY/ds4EZmeVPvdNLlEPX/+Dsa9tNWUmU1bLjVdEqMwbFZ7J4XXWrYN78NpJ
USdgtbTS1VJuuxK4R4tLMwU+uuE6C4rz2skpHFJYzVTlGkpPpiXIO04hrrajxeGZVHB20cpepqLT
0cV589PquRcPjB1q17BmxJeXOW6G12AhyM9GoqfAmuvQYm05BPFp/8/oRRtYzTuKwLja6ymXL/8j
VZnCncwjqMq6v0YqSyw0Z8Gl5ztd+Aj1p1mtXaZ3cEUmtg0bFW6qNiAba8vQFqhdW1ig3gFbi7Ps
RUT1ncV4oiBDRMVSg+Er4kG4gKaektQUBXZiaagkzURlqOj+0vfOzFZnrHVV3yUjUCegDlIXEkOe
hoJhIQ4yO4NUeQnnJlQI755UxtI4k869WSmuotT4ScxhXyNYqJj+s0KS5q3YX5Nh+bW1J4rJdjq6
VexRBgUzcOllRl4zgheiw4ae6ByzMhnBaxjDRsWyMzgz9DojL2rZnJSPjc3DkNvBokmEtgZyy2O7
COH6kKKQwufwtFeNGhtFAmneOrrhGWMh2j/pUIpw3OeC0ievG835rVX0cr0DgHpdkiWBcIw2pZJA
RzeywkEbBPUE0K616NgMJCyZF4IyvCZZP9XNjyNwm/o6i4bnlGJLyHaqTcMC/ys3F6jrdAlKtqY/
YSBijKC3Z5oAK5A2E7vFCTW5uVqDlnBf9uoCv08wDUXfbJic2Dx43hQhjUrlcu3GLKh8PDYp5lG1
+9pz4YXp6GS+JhvF5MKAXQb6OeQVUra6n0CZ9WoPCzQQWv2KYPlzcST+pNT8hGoyyRS/uxktu8RS
4sg2kjw0WPzZySLtd1qyIvyO6sX4qoXuDfmyNdfF36iZREo3UKNa+UbnWMzX7HUjbLvddgWX6GEh
t5ob7+xPU6qc7Y6u+BJkVlT5us7tuyc68ELjL41SVFi5WOGGul3FkTY/INV8dQSEuuVLS8YM/PJa
SGKKTZTYOrXHehdG0PspBJSyDCDuxWsjiP5hi2uWUA1g61XySkE73PRxzDxcNvzMbYKIO2uMLmih
W3KH8yy901ysQ3acOBbTzSttO2LmFwZe7MKZ/uK/ihU9Z3gSqoQYREPMEXruMJApyu+Is2d/dwsa
fl8WUUClKy9VyYE1drdkGOq51PR2hMfrTzYKdAnDZCh28zIpFFVCb5DxXoPKQckJ6sW8YHG/ArDo
8J1qwUmoJAlNNw+3rAOucC6yrCoMIaWUHO9fGYZjYBm2/scOPeaPboMyt3E9Hy392y450cOc/SNa
+zctFvKt1eD9tknNjeOOOwyuuoFsjMTKV/jWXuxJGeH5RSeHVsupMHJVZ5YfS/rlocjs7DOP1SWT
Ct+ZtHT/I88DhBNz0LYl+SKKBu6MtDvrZvhuVMnuPR0Si8SKmbmme+LzyyNa3m9VSgRcWiv0riLe
oyp8sg0Zwqpv3fIK3oNVM77sZyMqFdq7elQxVy10CcZm5Ms6OpJ3RGVb2I7aNEejXbS8qNHYmsKP
+6ZTDOsfiXfI58difwMW8YNPgYeEIxr7Llu8YvwVAs8L9ALr0RB3w2Q4ntFTM9BoEST/Iu0n/gwf
je6Na0m3YUB4vpZ/j1uMN/zBXDN3OCQ6H32wGuGKTSOv2Nnaf6UiT7aLMo38L94BHuZ2eeFjLanh
YhkY47yB77kb94rTyH+icAUAnEi6gOcYxbrfJKu5FxXleZqRDoTF1qyPMNT5y9On0qK+ix16vBMZ
uqfRWdk8b+9xRfIbB7XGvhyGtJabBlnNN1+WImHP+umBqDpA3W5DEq+vVsYqSnWElm9OKMOzu3Hd
3jCiuM1M/CLpzfQXvvkdEb/9AqqfB7o+ZLZBkMdbUjl8U79cXkkfSoreClTIj7TtPXliSLkLpJCp
W2a0gs9Y2uNcv6YeiEMXFhEQQlpEGJMHXCsKI+H1hZ6Az2NMNYIL8KLw4ROx/F229swBaF9oSxHM
x6xIbWU+tBxVB/pqmOuk8e5F6/zYTireWkPlK0zD7ArTVWRV4pPBV5MUD01McFtt7DC2nJ39yKaC
Ud7zaD+DVQ9crfzna55PAOHYYLeUp3Mut3r+0nAuogeT9esonLnL9V9mQaEVVi9Jtchmvfo6KPMf
VwC8P4OGTY2hoQKG4nOmiX/kOGuUb3IGbn/jHZoio2F0DiyXZnvvzh4i1OvwsH87JXfy6EkWQjLK
LI64Q4E+XAsAuIcmkcnazUkeC6VHjkd7DnMoJczB3Y0lb3/SqwWPaQ5pQngYNq7j+DJzMuJRbhlF
HDkLLSKtxOXFyz9pusaPqdafmwwe7GZTrt+TPNKXmWxsLz1pd7FD5SWhlRbjZNo/zmrzflUeJO/u
qQakVB6CZegRLq0L7Sr3Mfosly8BJF1v2u4mFFtFRbEPFT+flgVa7+ifj0zvGJY8HnmjnKv2WiQM
3YFrnxuyM27jHCbLLK/SEGPx+5Bb/hZGsgl8Svpf2sZOlOBGRMJ4EyQbf9z0oqPOjg+Q5JzDIOex
h2wA6HqJ1Mo477xlDtpS3XOO24ZFEdV9hUf4u18OfELWfY/iBEzvNjQ+QystTJQwN7PDLrwSj3PC
JrrYfHjQ7UF6IotH+2jquYOLhiOjfCAM4o1e0/GPh/wjefT0YrJn57QHfIGCaFYkthkYfPg8u+u7
6ywap5pLQ5bhNfRdDU8cI7Xijodv33w7TXUT0gJTAho7x/MJrPtuFjopRWUBvlbOXMGnAaxv/nlY
kOc+mkJVlGR5f5HXEV+S63B/K0RB21bsezoLu+tBzyWkdlxpbOSy9Pjt9FPlsGomG5knDyugBJw2
I/UuZPXeBhabi3Z5rLZnmFGwf84s95FB+6zMDCUBwHeSGdaXpRW/KXU0fpqS5KjzWfqellsDgRUm
GpwqXwz5v0x3N2rFyRnwJNB93NeV+ERZlQGc7RkT8Q1c/hkUaJCle5wx3DPPfQMhqAy96r8wFene
Ac8ze8bj9vB3N9oiuTK54rQuLthrgfuh+GAMfB5UrxGADzAdOqnSb1yu3LuXm1g7ld52D+J5bEYH
4QIdSXRgpU1bHG69fFRxGhdb+llnIx8j8XRtmr8muUCG06AoQ3IRfs4wiPX7l8mEFEuhOaLOpzs1
I1bWWg3ivDTq2J+yhcZIsVXJPLPeNIHBJFJKDYsWTNfGP25H5Z8VKjS0AEvkq16kYzQYZMdzNH2e
/YU/azN/KEuQw3SJZDmk44sgZVCWC+6ZmrLmRzhjTjmmDNw79hLlrUVDcMN6lNEshxhhxEhahwak
EgjB+HlCIuxomWHktt+K8k9wN/fJ4WexKY0C4Em/jZRxCtQ4/TJaiRD+Jl+5ax2sCYFcOvpgG1U0
lyAevnDGvnhiJe5beRLFqMsVElK9eviZCJbJL3vIVGPcXWAE6WVgS/teGQDY7QyBYUnD5DBNzU5d
x0COePVPujlAE9z1W19ywXtE0F1VqJ7QYN9SYaRcUlW2vpOZuT8hQggjIO0Jk3dZGh3BP6CghMdj
H28Wwp4AOBReGC8LABzP1K5bpoxSFhPd89xJgLpGkZpFcdw/UvmxVA0VheiI3iUMufFz9xU3S03F
QVehuroA2zAp/VE8dKjNfgZGmartZiWlFOEJenSlpM/OVcYbsrAC/Oq0rp8TcP/R+iZHkNCaVWuW
DMR3O84IgCzywUa9kf0t34qKWPFqoFkOFqtuGXDqUO5K0w42X2iXtoYOc8jru1sRfy4FJCWs4Z01
JJvV8xOMzTrdB1b8fPO6nE68CuWaOtAAGmDtQVHWzRCafy0mlUz3BsQny3k2qU70ZMUgROlVuoqC
SO+z9BO+pG7O1fnzqyU9laW9CcyGNI8aF5VLQeZO/zR9EjsLohb8mxIMEQkNgXjUiKMT8z62eUl4
eEV7mrhGDfATA2y7Nbu9Y69SRKZMoM0eilWlC6NvF8Nhn3V8wH85eZ6fwuLzgdkEJCoSaZyq64UC
eipmBCxoda//hVKWbbIfR0l76hlAk5X8ChL6pUcOdPWDdu+p0zj0fZH+L76wWb5YJeTDL1Hkqa0o
7YuQTHQpTx13MhsYBhekKyjcfBdFGSct0UBrfNBsJ+U2jbiiZFIGprlPmG30ESmvx68MGqGax8Tu
38j12PbSr0v4UKfm9l84PFsdwNI8kj/yGHfD4Z+7RmRNCgEPAtVYxpuFdN3B85wYZl7LForjAH2O
zZfiVTejAoHwDO56aQvPuFmBMrcMWY4dRQT7d7yk19N6VZGOzGtdHtB2oomzGu3cx8PrlArSMEiy
bEGzfJpfUmkAtgQeYLBAjFArO+YJ0cZoNq3E8Z+ZnntYmiioIV+lH1PxCSliCNceama5Lgr39xrl
1lmMGTHzKLpLEgzOk7VTIGs23IOqbLFXlHPjj7RghsMW1L7et0QDRi2QnzfS9DF2vhER2apeDZHl
v1SRc8D6qNohGGBU3cZ1Cfww8WFbeonoyDXWkpGZmS0dx0hi2ut/ITAhWf6hgbZsfnbF3RtW7X/D
K8PXmS3x73KRWRIML4aUlHH4VA7d3me+hj1agZ9d3ajiPlKpiclr4vLq4tBUEEqDLsLmLzVfMO5A
Z/FTdsBUmmzNDtozIxlocCkQn+CjmSHtKZpPzYwZr7J5kI59vlCQQA3uNyRMrND3ECLFdmJxatII
BB6csbpS9s/WVMlTU4046voWq+7W6u5qGdquXtOdIi+tjrQqFB2Fr4VdUE2+bGGD/Ag20qMwvdL3
py4E1FqV0UYUWgpuEIltVv72CvbrS1fWjYzoknTv221U8TLrwFZgBnZdZx688jDZl1vBUXqH7tDF
CTnZP9kZfOQHimE2ZAAd4Wto2wu+3Q0SS0jCXotXdco36suemyt2wW7FSN/r2Q4XQQRnk31vTgsD
k7iEq0Vd3qWlIyCAeSYDCSwIWGEiS1u6efve+0WlsGoboWi0l6UARklLc6ErXj4b+pbkUvMnUjBt
lWyNPoXyoFL79AJU+O3jnqkDgQ8WZN8eXFwBt6umpwEh71xQEv40FE+8nvZZwVU0EVm7GZ20YYrP
AKsrbBoRlJ30jiMkz5DkG1PiRhG+IUJ26JsDWoWhXJX/iyLMSD+bqgWVVuzTU1xUK1IjVb7dTgpp
URqd3TH51UsQB+UFpL5OnPb32hC3h6aSSS2spNENQF6KUcMdUHiRD0SaXLRDiOucZXfPDOOUYaoC
69eUEGqsnOU1E0H7gqNR7o08b1PjoLolgB2iZwdfJz1zONNnrXn/Iah9CPrHo1/W71vY6uhd/UDJ
VjwZwYbE8WaYs306j0IDIaE+2/OR1pwia4FarXEV2ea5ZQ5EIrzaFq2g5UokAVw+GrVnaqm3oLHM
R4oUz0fUuCJBxgTRJSxl4/SpbLuy3MyJD0P1PWoCF+qwEvlHC3yfMaesOUqVJznOFWsKJJ+N2x6t
7duz+VCW1Bo+86ssOOVZZ+QzeNGAQC9ClTqGxiqFfS9E+/9cev6sWCPTfmHC8zYRPqK3xKOqONjb
w+R0eGHia0jTj5UJ6JUqgKlgE6pD2NblaDIXlB2Q1g0j8I+Ku+qjel4L244BqKXbjh8gT7RYFHW3
gCoAB+THeq6rj1C5Mg7uBPJJ43tWF8Syv/WC9nVloTmx9LbiYpa+a1PgJxpj/wX5jwzi3nwKumQ6
MrZBILI3rpjQ9VOeDjz8vDcQK3d56mSxsMSjPV3C9bB83BEMgpmljqxoEv2mYwQNJ7ly5u3n0RL+
QRS+yJcn49zsegS15DIWxYIZX7Su8EgZorjg0jmYvSHqRlMcGHtP0zcy/u1ZWhFDIu6DXp4VkEAk
54+jTtojN5DwDTbL4J5InpxfqNqXqZXgYmJNvGxsUeP1pg8GR/Yz5jhQzhuBySmUCe/JqS6Y5c9l
ePZ66kRoMVYTeKYsRdbU21FusqnjltCRLzHqsaihpzAfawRsC961jOAm4aIfs0srN4Xho4W2Pi3j
sbbrFmhvZcmCCrkXZM16cQiJPj1iGBMt12y/mOLT7Po4KV4NqaQmzZSw60KqJwz2j0O8qy3jPKGH
V6b+cw1laPmra4m9TC1wqR7plvpUwnLDIgj1JpjT4aTH8EaGGH/u/y6FYaQWE82yIiDGARlBBtEI
FCoxJIRESu+pmZ/riJeqHL1rZMdyiEDgl5ReRTD+fLwL/v0R+hXHUphUUwhCKuCWtL/V2DvjfTfE
q8w1Zy+SZ9cdy1izPKgNO2iKMU0Z/PqC7iiYCnP8K2lAR/Oh2a0NF9OGs2qj8SxKftf1FPiH+TTm
i2aAnVHEy+eFskLiwehPd8CCd8rGsVBhdOZrhBtXiCtA/utgmlRBu1uh5cxhnUPVqj5JGQpwKGjJ
CHOlb9ggCJO6biWj0jnQRDSIUnpxqimWPK0/AnwbvOXrrJPPgnrRlcuvkiSVwvrlwvyopAwHJhoC
a0/lIj2gilN24UH0XpYx7hHiVB2vzJPybazj2Z6naEGxmb+j4BkWRxy8P+LMz/Isaaz5W0FR76p8
jHZc53qoFiyXYWeCazgBl8ynb55WrIdm5vu+qgkVqfLx7N+B6R1NeF2kwNQxy7lgdPgucVjm67yT
YD1lJDJQkOEebWrDkn5uC1mAgJ2eRfOMKVhV7c1MVHy+8pacterjYnJL/SX2qDy/8iF2i3GgHqIs
l+ZFfryyKW659Sl6uU8oa0yzhRS4MGjQCHd6yu9WfK1UM6RlK5BAURh9wsfn/fE3iMFhJ1vcb/gZ
VIpsIFEgc24jhS1usqn2ybxeUIrLONKtClBVwiSXm6Z32TQuBNoG1xkNqiGWNfVHbQLvZ190TdiG
PcOnQHrA4fmAnW9HJ9fQac+lVZ1Ja2lQQnnEJrkUN1nu68JfWs/6dMYQ0vgVaLNDSY8yviSHCmmH
Pcb/3Qt7p8TrIxydNJs3s4p45VVcVKbaHZE+9CAboGDucPJW0F4eKMTLjOd/9Eowdw9MtFkhGcNA
kEJLX6IhNLizseWfq3chTBhpVoJaq4sHvKPC4jGsSdVQfXaRVSyOB33EGqqovg8q2SMAVkyxS0RV
FFBVKq63Nu8sa+8+T29scsTj+2UGyI+Mv0SLC/FIz/NkLD4NItfqtR0pHmniCUjYi16BykzMmORC
y7DZwkbbaDQJSYY9FTNqcb0WghLWL6Jec76u8xk7Ir8lg2iU8Em/6WBn8TU/1pQ5FseWheNjsL1J
tEstTvw18CCxY6Q4fFBX5gf1FGBYGFsdmVY93PQwFcfMWjIAKGRUFQ4oYD2O1ylqrJEB7GHUfsdA
a/yPdhAToWW+WwRIDCL3IYXgQfZOqqz/myxuhHZM12XZEmMOETGwa3ZcY+oz+ceVWib1hTGVe6ud
JKzQDzYkqyPF7NS01FtgImA1VeQV7V3FjLl4ga2c4CitJwhuOTGZ8oEHo6V52ivWWkRyujRPpNQ4
dV64krzgh0hVVBoXfmpe3/25ZALl16v5FvYzSMhHunBesa4x5l6B9KDzZ9FVNYcm/xhuHTz2wuz6
KGZ22IN+GhUBRwplEX5fznGRMSgEoSxRaSQQ1laMNrwaIcktWjTjTSf+GOBqIIqQKASoa63HEZa1
JcJemVD1Yl4RUYslZZ3MsSuuZyiBIrthLsJ1+fDBdH8jePftQ/80hPeNrtQgHnBk+WIBNCYBLswO
DxI5s6im8xkTpZWmZuZQuoYtw3Cpe8MEsp1bnswvWPm9bgHN4sIy/sp4PLWZATNK6HJF4rYO6S5g
JD3d510Aya7gCowJkaBimLx0CYZOjaNMki4Mu+KW2dfxigcHuI3FzwntHSFIazJqnoykYDQNuTOV
jABmJmFOs+P9scmLZ5eDMp9q8COmArUNmZJ4RaiDqFqeG/WI0VsD2vHgU+H/N6KMk0DgubpDP9bB
IUxuQeLt7G6xY/lDlLZCVaNjkHDm5drYJJRGWPHjebmeqZCldl6wMhl4aNB/1Hs9LnUGfkUGqD4F
+WpEqKrZF2mDWHhm7YU3btF/HeJyHJnYoGz8xighWCeDo/u6GVhnzQMyb81dy8UYTulmYarLEHH5
QRKQeQUSoDCrOyBrBkdBY2h9TlJ+q3K0zy87K+rkY+ZPPrFEfVKOI7r7mWg7HjGZaVJednZbCAgP
GjPJKzCQ+BuTm7DF2PoldcOO3CPNJw0taJ5RGa7dOtcm+s0A+zFvu6vt0I94LZSRBrRNV2MnDW3P
T5owGBULFnA8R8Xk9dGujz3DE59R06ncxbM5R57EuBjnTkCcl7JOtT8JquoC8j/td0+nCZRs3Oby
OBumPWYdpGYFbGS4mhzy++pX/bLpYa8W2/A0F9Z04/A5y7paV2YB5nyZDpP3OhVYCrtlYixGNX9v
C/MpnYCy/GBvcT6d8Lip0WrFb8OkeIMrxjbVX+cBrIqem5FIcMCxb6jik1v6Lt/ATq9haJqcJYCM
vS6u2raEOFlaTgqE5P7GVQNAkOcFY8WWClyOa4EEaaIiv3B/tQJaXdVlpF/9od44hgY18KIT2uRV
SjZjod3GxQc/5wm9FF5GMlNUL3pdS3i1vkGYcrobtpCN1DltDu2JbZATCo2mM6/nR3qroamYcNAZ
vqTYBdJitZDo0yfJOd1KciUEQp664X4kZNoa4+xzf5VCrumZMYeLwVkISnDu1lViM5MpSzHyJl1u
8AnOnXs/J6fSxTo1Uhf17bjrggLmZNlQL6cebjqH9aDBVTv2eUmk6kCG0PYX7yfD0xEdDq/1Vx8C
EsLOfIGp2dA0KaRXluN3S22xFizCQE3o0bRBdF3g3u2GukUYXLG4hhJPe8p19vUwIHbeZK7cSgdT
/P6R7bqNKrA0E+lK4wVncxfdrXAal8abJY3jT8cMzp/IGQrb8Nv52sF/uTvGzOiOfO3NNujm5hgB
LuEbxYapaTZEilCYcTQ7bw6PZtLVzD8haei1aRl3+ywRSAF8TgBb9ORA2uiXH245Cz4kgWb0rFkc
maUIHHa9wj9v7GapTKpZkqnZiQVPkTgrlUW+TqU01R3P70M0rlL1DXj5UBd4PRUSSxdrTQsAUZN4
5qtQIkk04F/oVUGO/o1NvlAy1wQ9Hdfpkxe+IkUlhikPjM+Hs7XuQHR2xEDSWa+WlFyrw9rKJtC/
JGJeDngux6cEp0rFTTISbm39dvMnjU6D21grHjOEJ3dEgQE0ajyfFNpSw4rc7pkfG638klYZ50O1
eMtwgIdKRQLXHPOCFVoyACu/a6zIijt+ZbgHS6yvOSN/9VouzvmNPPBy57xpgZ05Sz3syiaHBsak
iptmNzTtpa3S1VB0fZvh/MchgmyqhyYyUv+05eEycYAHjcfiwR0e8lfT6qIuMZ4X3iJFWiKZ05yB
hDQdY46VLZ/eW46MP63S80FfVm4Alxk/u+3HXtRT1M55kWJJGwhGtxLrQNZzY38cp6ivyDbMpAZS
MAERpDg+rIckJveZKuTt8gqcDSkfcD/9SbjLkmaqRS/NjETmNsZdNS79Wgxe0mHC9iLO5i97uQeZ
b8vjldiG1zMqmy1JtceIjig5ZCyc64S08CdKc4vOynbuHT2eRu4Pz3BN0CbWYZzcwU3eYHfE56qO
0FN7K7B9ia9HhH/YC88pB0/gEzoWGngG06Z0wXah/4mhJ6qskvEB/fzulxQYg6Vircxengz+MViY
unFHsPjqlEiD3jHRCto/Z34GKjKcMu8QLA9IQM70jcifwR8dXvhgoGUH6AEL4rZmc9YPeP1wz1cY
avgwS7WH4ktwtgH5ruOm89peZ0zJ/7UzJPmJD6yxZ/yFMPViOnV/vmW9MO+511KKkpjeDHFwS8XX
IHPztoVXYQCK043bcM/gKktFzIEwRhKfT5gu8Cd0O4LLtpQ8ujIqwP7ccvMfeIFcwNuxAfrFYc2l
iWw89QG1YU2uPttp8oE70mJSD6RyZk5K9nH7sfQ2LwC/AUsrnA6se2jncoLwRWeL7JBgFVeK9GL+
RAVjzPz1ixl6Z4yV8aEIbzl0iD29/3xLdr9AOifeqXB54H1my71zDFk04Q8AqVC01HCpclvXcW68
w36HaSOKX6QeN2Jpjdwg3aJniF5LGGRwOkuvVHrd+nMumHKp27cTJUMMYU9CDla2U3KDjkjSXT+O
gcJOQyjKH1w2ix1K12AaZ3X/zH4bOPgE9of967Pt6V7LkyYFnmPEOdGXEsbvIcRl+ir5n9xka03W
Sy6KQpWOoGJAgcjfHfdRDpc8JdijJcSZh5NYR9tvaJLmNz58c9HQdN7MNJl13C6/nOH2pnD0H5Ft
bOwiuIgmNQztdyq+3pjwobDireQQ42dClkTYdYQXitSeXsymnqV4O0LsVI7gpdoYpnQMPliPfosT
4SNzrmvVcW72BLuobqLgMxxB7a4u0Ht9xei0kcmgNw3Wl2+Om+GL38ZSoiv8wsmEly6+5PSCk1cs
+sVgBw758z98WRCrv+9vvrz+TzKvgevydija4mYfP/PHiWKy1TadjiPc2gdX0jRIBvpr29uvg/1z
bKz0Jyo/HlAR2cEisUqWYYWrUXSYsm4+r0gFU5TozHjpKN//pLYcpzHFz6mCOxqos1f4WR1beXpU
WHsrP9AiKjRO0oyjnaYXke6jE6eXxA2y5W2azymvfCJl4wXfEKhwzMskqQFcTve/PQ0Psb+UN/9+
PnRJN49eDA0GWmnvehsbpk/83hcUOkokoel0AJCCc8XjscZ92QfRRitDWJ8syARkv4i9pXdMAnhC
zrPa7DC7nwlIc6KEQkmqsRMg3RtWfoHYAlcZTbfnSOWmiBQ6E58Pr/HpQufuIiKAEyM0XmOWQBEu
/dQRfJSry/3BhrtvZVjEtVtiPR6lPe8rvU6w/lw1un0wQZJCEIMN0xk8ZvSYgG5daHl1rv/Lwxzs
D1+Inkcezl7qBujGoZHgGdh1uUedJGXcaUYWwT3kQQfPWEt6FDz99KPCuZnCJtDVTiCMNPmwcoJ9
MUYTj5hbjVoqORM+w0iPaKGUR7Yy8xg1Hig0xiJE9xWzFfNJlwviHZ2xcWi9isz0GC1NLGlT4Xml
IwaiVfPH2ayX+CmLv7oeXtzodYykFTp53xEnzlh/vZkSnW4doCanCZdkei2UaiarN8SN73RwQKX6
Xz7HGRVx7az3W6wCm1e3i6jnIJf+oEPtCeKAnTBnAN0IZY0/V4T2fuZ5ucegMRB4MFilTPcL339M
6aAZB2euxHSJvnT33tYdtvlnZhT9Wz6cBudUtNoDfi0eLFwJIL6IzvvkBcDNVGbDedYVHoAEMTYT
jT1B+51YSTf3yJ3d8iAbwQptgdl4KPxQfasKo/Zcq/6J8D5PrVxV33HhZdOoj6AGseCcteBwuXIT
NY/swczVdf+ngQfTg5M/Wtn1/p7CiJr/7W+od/HMZCc6yYVn9W6519FA49jBH7+l19RNLu2rr9nL
DBMDq3lpqjbJ2sgpoSkTTcJzmOLK9KTPHhVBA0iTaQX69DSMdvT84m1huvHhC6bsmOUUkdr4BZNh
/7xjTd6qO+d5dxDOMR5/kFw0IZ27fNCmKHLLDH8L68wI8KHrAehf+lqGN/NfAkxPMKfqsPuYMmtb
FQ1DkFnB9LaMY02BCVtHEOR8NAcmuNZA9ORseAcbJV3SDfJEENkZeVPuIz4zIpf+AfnAq9G/HbcY
CGGthY9np12PKjGhXx72d5LHzjFPAPQ1RaBRBKOgR5/YJItkDWEVXHhQoCECU9/RHiBDHTEybK51
dz8nF8f8Fij8hJwwqFxddU6FQ74lqkTO/xxWKwfVqSqad5x0+yI23XN6t1r1kSqJmuogc7xgpvje
ZiSCFsnSSAGqSDh9edC/qvlHj5xDTfWvGem9W5DJhHU9vgbI/APAb03EaVOB+IKKcJBdZ4rHJsul
NWdMfLent0Zry7VMfYsQxrxKHQjTu8sqJGGQjA+Mz6MpDvlDoNpUcCXb/RJeXAjU35uKfc9UMBDo
WOEkk2XpbLWJCUYnyGtItJ6k9b3dtHTNMgaW7MdespgIlGQeVcA/agS2/7ERLBKjU+OzxjG5drVT
b1gqa8xoxsND3HkGIddHo7o1mSwVuT6CPDIr+xVQSQhSFVSfEBPnZL4e1c+NGBVNcKR0zNnr6Hl1
tuNXA6n6FvZynwtQplXQkUvKgba7tGRYzfippQOVppJf5bOhY7/cKQ/BFy/14zqZ+iT3KuihyG4Z
GoR8LRYuHujKSmHoU6ckILvlHSRm+tuPVxb6UrB+233QWi7ubQKwQ/uG+yj2t6QaEccGde3SeXUW
NpxzPE6s/k3dwnueWn9rq+U3/zhBsS3SRciSK5yzPL76nfoYxKDx+Iv6fBCgMA/E/QGWN0btAuOR
2aD7biwE2OeYlmVxJqpC+GrV6bKb7B5ixzEWqN5UJXhUUVvDhVWkPvUmB2/0uqhogiiVoaft1LL3
LuzZFvx5hyZrxdvKYSDRo7HtFsBQRGzDQIr5Mq2St88ZvsPAfsI0VDY2qm0WAMDD1T0xYShutxuN
Sjx4lLqlM8stGDQp7HASdY+lZ/5zT9wbLpvVnZMdYl8ttlR4k8m6VkW41TmKUt/KE+vMVAm/oGiX
aFFEUlv7DxbY8M5tQGaNn0sv25H1521AUHn+4AqbEoXP28Ysv75s28U4bcbYAxTDywoh9AkCXfE7
DjTENot/U+gGsZFBwzjDCDUfqRqRtBYhen5m/UU4fJ6phozd3aIujOuEGN0+CK3sldP30VDXyX7P
xpgvOOXKp2hSBGhx3opfR7DbK9DPDyGmb3OuNGcpHczKHxaheAoZJy/uwi60s5Ey+1yGoANArtX/
bw85o+yl0O3LpR4CqQGMKKnJYOXQRbf8vdZxRks8qvN9Xzcb/0QdGYqMjal1gl3F/C8MCxcYqapQ
tqwC7WsnKKjwKygw5pi8PEky71SavfwqqNKPrJmkNL/vTemh2VXOxOCqUZ4Z2GADvFVBzIyO9Ugm
Yu5PINmnVQIh54ITxyqAnks/k1jANm5+Y2BcbNtdYrbY9gIPR5Cbag19BIjueW2laKv7xl7j8S6G
3ZD0RXRs9AxOqLIxwEZJPGTtPJkC1xV3HSKe/moTj3kcV/kYrS7sXkvrCB3KfrUdZdpZ0/5ANPC8
V7f2MATatyb8T9DTK+Z2HotPJ5/UcVqGej+RMPmUaVcYTOnE5+SDCwes8N+idvsm2vFLpKUPilkR
026DCnfMzO+sbCsfFsG3BeFFVH7t/Q1RgWKxvzFiL8IYTsPXT5VqHskKMwYeXKwJ52JH5JMVma+U
JbDsKsyfTwYgR8k1kCbHqbirTkdIIJCGng/R/pFqEIvBceJj/OvZgOe94XfPg+KjAsTeIo0RPuVp
6Ki+rMx6GFRmDcrMOSs5W2Xc0wNCjCY8DzhagWd4MdlKBRr2WRCtiA1hrLbiApXEV4h6DQqsmtV2
I3MhtBdalnUxsTAeoA8wgZHdH+9LRWHmD0r8Fx0eGyF/x5Mqs/OH2x3CccpjOEVaFPZJkNUTu4xH
t9uvCTyEXpzoGuVC1hISUPvs8aI6v39zF55lnKubflHQEQD63iuvrEBzvgRbSRAAxxmnCRUv0Iv8
OhvTa3mNAKm+Z2j7k3qvhifllkEC/iJkqnvBpb2vYcYNxIIET1GtMAmhwIu2QRe/tRxUVf54UfoT
HEnhV8mzliBRYfuVL4JlwpSPA/5bH+25Io/LQ12afkROo3whXx3Q1ufUEhyj0G0CX8iFbUut7ucp
Tn43T59spbXQ4vN84+7F+uQq6ApjxBXju7BFNAlD33W/GbWwUuSDUa7edQqr9P6nl+1Lr3KOjzWc
9PnpdUWb5QObFmY7UDKKIoY+pyqN4LguvIiDCG0PQG28swNaYF2d25hhdALhhGVh3nbIALsHZFe/
3TNdtIUiX9ut13WeFDcJFu+jBRnYzXBXpYayqibYddQQfsyvx0JAWBzjFct6/TYAFhuRwWE8ZfsE
coiU0IZWlUMy3EPE/14RB3Fr+ozsWuCU4LwXhwPReJMUchIV+7txxlg47D+3Tx5XS09q+CTLWa/o
Ihep5HHPd2SO7Gjtm4G/txxDo0dg1HKvuhbKztzJzY56ki7wWTAOG0Jn4PA7xgGKwzx96hxIoEe5
Jk7D+1L2S4kyvpUC+zcD3sNb79bCVkTqIdNoMqdTndEqKU6wF21U969s3zY+g4jgGCbmJ37LG/LB
Tym9/MXHSd28XOAn6e6RDqeHHtRlLGP1W/9oA7nt+ZCLOkh+hm3o3kFgbMDJBfOfIRvjhDEK7GcS
ehR5xc0VjTNaCWCas1ulPxmSZW8AtP/A2eVywtWBossUna6UJPsGn0mDqYVUuTuWMEJGeepFBowT
U2KO0dKCxoUcMevZoJqhUhuZdzP+6Mm4PCHTFq9r7pWG2fRL/0oHsl9us5ub64UX0VazYqC8PCHY
yyubw3s3+j6g75ynT6SXVMxyZlX3sgM9jj5stwFfOfBcvJn6oZlLrZWdxv+Seb/ma6fW4gaO5j8m
DkQxfdhPKQZMKYAM1kn4Xx1U/ntRczRoljgK7A9BpqBFYw2B+/384hur3nMCJh4ENaj+w8h/DyK/
1PGUBktk0+kxZF5O5+B9xQhkVDzzMyxXrspXdSghzz6Zy+I7DhVE8ghAuHflXaeTGzHYSVCfN0Ue
yi/Uu07jKW0B4ezDGZNSIX4EX7DHEg9OIMHEtZlTEq+9UMEDWVL3b/akdYdBbi/BqawTUydM9QEu
Xmy33xGvRy2tet0cLTxicWeSTyr0JjB1DkKH5NsCj6zxwzVb2rfNYF4NOp/QVlFJTQG3QFzg67rt
p7zTSNzIUpKaP76KqvW8AKqhcBNXSl2JA6S7tZ0MRYgaana1BorOkclU2cwuhnjEyjy2+Esi5AtC
I21tcAPiTOhx3N7v+0Dwrn/wOJiAcna1BAeFmddvhSdadISirYu8/nvv7xV3qgTCz05mDVZEI1XK
Fa2ufrj1STgIJTkZuSEUgxTvXZZsmHfQefHooMOizqT0zKo19I66oxWkD+fWYqTil3pO2hFrxUgX
NNXuUpKyogalCs1T8TBvjYCjeeOOJJqWVSiDGN+AUlPh8mIIeWIPiS5eX75qQQSCttvmFXp2czOS
+ZW0xIaTPPOTV1nlvPtn7ZEIE+bXcIuMtp4OxelYOGGkDBwf7ysSeKLH8GGRpKuyFTGSdC8mPgcn
wQxVmpz0OMafeKiIuy1TR6Ws6727ysfBKj+VP/ba+J4Hplbsmsr/DykOB1ll3ivoT9259JkNStSq
LpFnk9M/95mAiIxiKzYXCkYk+GKKbLe4OkB4Swf3krYphroQ3J7FDRNPFFqEz8kVXBnf4HB5Yknd
3I7Ql2IsSP9XzyeFhpwV7yF+xPOSPv04QVaooV44l7RtO7d9RShcZq/erFiQqCPsq8OlQiIpFzgS
EzpQJmw0v6nsQ4dyhuNXURKHplLXGy5KMD1QBpR9DgUyvT4bhkPWml76IXijB2A3/rm5VDn9E3Vp
U4/pPHeqJ/083i+gFZRdAnlwypTn5TEzL8EupCjsBJPWfZos9YBG3IsHIZsQFVFkWRhMgOzOjWaV
x9ZhuYyzPb5iyllYyCRaxYJQOWv1miZ6+wd0/M1neTdkUnWuQPmpxGtmGNYqkvxzeki6hATmvqsW
cpkkAAjG0dPd4w49aS9/yIaZSl2BaHhc528dcG/ziWg9wakJdqLdBL6LKUR57Oq0SDX1G1ST+JnX
BXx/VAaU+Y//dtT1dMWXyxMh/JytXRtJgLTF4ugqY8/xo/wLWXpq82LD/y97Wi3WnVXBS55DmQ7J
gEfHZoLNXy0k8fqwq66V4Qu3YH87hn82LHQPyRLSiuC8TqA+QhCa9YJ+aQuTgzW/qAdfM2YXzWcd
7BhTPZNuVOdprC2s0wCfBJH1XkaUmLYshNaAZCnVj6eC3SrtNw9X1EoNaZ1SEUsbgZXNJ8syZEcm
fTAZUzx34U41MsupD6KfUBdf904Y9zSQtSEdpxOCRQsFmT/ulrQp2aak69maiLPa2BC6Tu3h7Ahf
ZDR5LAlcS7WtW5lB+4pl4gwajq2/c7hPeYov+7BUN4MbvaxRl9OFy9ABdjFs2R37FK7DMJmCggoA
ACS+8Tu3YKQvCcQo+cJKhsI3lxFcTPp7XHapn8AWWKOvvifsUQposSKGysp+CNyd555YkYjP+oo9
98mMX+VPP7YzqFDb9UKD19uiKPH+iVnRE3g4yYesyQy68nc+NPPZpaB/USkyaj+Um1+vzESeWu6v
fbUDlB1nCwllP0JUmnTiL2jmk6eIRb9Q99z8vhUk8/cM738NNt9EDr1Z+UWcoHQ8NHpbZ5g3DKmn
2+9qUIGkRdSSXw4e8EcZ9pop5rPRzcT9xdKB80VE4mFUlN/jCt/vHjGlbnEJCIe+eRpXd6mzr+J+
dJlS5rHkS9V6jBXus1Gv8mRu1z5Vq8+51XCx+IrHLtTAk1sG5AlqyU5Vwb3nDkgzGkTB/5xz26+N
YjCb6LxKcDq/mMG8FwNG/YUrWaW36H5rbI+gtbCD3a6M4BCNaLwa7QaZMKCMgEWYYsqu5tLWtwCw
aChejlzSctgPiDA60EdC7R5UMlUPw8W/9nS9SXzlGRixPMfjXwHQVoHvmbUsdnD8SB7YObhVBFYR
kU25fu33cHhRgu3sn9vZ/QAFpwnCI779uCWDrV39Has93A5OlMuNN8gJMz1/OCcyrBuLEtaThGJ+
ckOhZ22Sh1cQgUImiPucYWRq0tkJFFsZvsK04vu5iAIw1iteeEYM2Ge0LnyzHjqQIC+wXn5/Ob4b
O38d+lx/DlGRoZsZSpZ6YM2RnY3iC7cOUtkXMeg3pdJXBTJnylb8xPUUNPqjWbrlu4lWmewXOBl8
9YoTGVPUlJ6kSs1Pw3sp5Wd2ue8Bv7qOo3hMJaBRs/FjXGG2fLcU/0j7wTXASoVV/MBs9Y76GX2S
NJrt5UsWDhORe3h4XHaO0UbQA+R3swiCikgi9VHtCxe6RywwesVDSG1WxXqjtqtbydjlHGZEKo/q
ebVmBgy6HqoP2MI5Fe6Ms0giD7K3y6dms7EQPAMSVX0k/mjPDADdstugyxMrkHA6jDFIcNLMWrOD
h1ffhKMRY3qdITeENM69NeJbwx03PKiaa+TKcOqd6C2lNXfo3kxdYFESmPsi2BR/1giu3NqQm5g9
ChBD1h5i6WnnG2HDj2vQ57coF6W2gqnj0fy8Pq+GPJMnzbJr67MQ/VaCVhYaqYCBZPhmWEq1c6Sf
pppgtKNYagHzYiZHMeFr/tCpQV+TaaJYIzv6iDKc7zLliVK1wnbi+Rk3mDRx610ECwlNwG4RtSeC
USM5RbRVXX6JMecBq8U/12mmAAhRBQPZuyx4+bPjSBxCFScm3617mhrHMO7IwfcQVfl3USQF5TJT
poePkGReCuINBQwz6RX54fhUb8j0HmMOHCJCnEQfAi94v0WTlz5UvZaC842abtbIu1nBEzJYCDLw
xkE/Wze3/huu+PaYaKWkhY4bPE2xZQHIwasfIxfWqVWKM+gMdyb0dNtlgGquGT3NNCLB2VrjAbDX
nfJDDWTYxUt/nv4fSAqjHe7hDP/jAekFcGSps2R9hphR7+pPtPkDaAuoiB8hAyFdfIaumEB7YxZF
SnuQVCE2dbGhJi3pdwpnWy2Q/+ndnJSkfsEATW63DbKRPYt1wKkEtR00erWevebeS5VBWLX76O62
LOEW4ivHn6AIRWrCrywSlVj4RusHJZHUKXrSuwFgzBGhgthCQ+21zUCfiyD5YsmTZB6tY7Ck9X01
cic49Nl2SZ/yNOXRhqVZelMjUGNggCwI7fVIL56Dhk57x0LKz25nWqOgqHlGRuZrZKtg6Dg3jE4P
Z54aBiN/v4JD5bl/G/5AnR59Mdxy0qPozOy2/g6gZ3/rD08mY9byMG1y5y9meL0h7vSFfAjGGqZd
UPxmAFoXKGAHvnJAJTdqOTIAXnXld9QtrmhERO7b+3nXLmBtrnARhp8HwpVduy4nbUw4ZI/Xsn1G
25vn027Tm/ONZP8xaXj+GQgnnIVIVgZWFBcBn9+a1LCdoKUZnYJ3UFUS0Kcpi8gmZV/D91IeRM5u
qnswhEbv95NAQ09QWJtxe3JmlgaH34pkGskBCzhGgZ9OJcn/i5efcke/6ad0VXBgSo5pDR+9WgKF
2SYMdBNdwSyyLD0CG1tAoCCNlUeKa06ezCcoKhbhofWBZUAt8AXEGdYK1v8mLKdPXK0+NKEmTDne
bavzrMMRcTnj3Kad68HwSt4VFIdcpfOvTFk5DniHyhSXhaHsdWTFvlt73MLum/U4Yn4c3CgUgaf3
qvCWXpLZAB99bZXbyZtIX1YcBvbibqFMuGNxwDJLw6iFQfGWCDDSKC08/0G+K5MqfHrzEowO9TOJ
b6y/RuwIc4pqMmLa/wFs8u20y2WuK3G5PX3ME9xSB7E96OW+hhmaDCbqMz8RiGYRsjf/ux2X7c4H
dYgd9Q6SnlHV1/bAZGTSBIrSfvSKp1J5BYLzdxXD8AVr8gg8qXT4rXSB5lfWBRQ3PgrUAIH5gIv+
/NU08HxTNb+bDUP8F/x6IUZCYcGuglgq+dnrN64fQk0/5q0MCFZwVuZyQ2RsJQGelgnluQ7Wt89v
ySVAAmQGdxJke/GSZHiUPmTC+Y2bD42YvTAB9UTGb4PpnyyEphgMcqBip0ySHoHZAPot8BlTWxC3
WdyR8gl5EngtVR9vizwzg4nAZ89lFPuF7GqOCWqWtYSnyM70TFRmOWQR4/dRrAhDekTapyL4PuOF
+wdeucCMQIPgCYzlHUqjyUZFbAgcgU2v1cq8X2zbI5OKVqrjogx6NhBwEGv78CrwgoahqcP+XE70
o53QNf+0NXJMgyLjWVBre3JdAWC4qyraqukoeguMqEtEm2b5+DwuTvHg+qnz6nCn34ZPLIxEdYhh
ur17BD8+js9eXUHzaXijq8HCRfkPk0HTV+Zz2jv9/K2p3TRO8/t3H/xGAj0ySNpyKv9P2XbK6Vzm
AW3jKiscqLPDA9vrP+1VYccxSYt5BYc1YCKAWMuKC76qm/OzUo4CHtXKe5QlmXHbA52m37sSRjht
5GiqS999JGWs+wNfFw+Uvmmt+xuU3XQ5cHpqPnDBnTRCzFozfZ7SDKCr4PLPQHxdZ0aUnopAMNFQ
mD3FcoIqK5qxDNlqd9+mT08widiAKtVZzCLWAXgrfDB47jDQ/wjJ83GUEceZq1yc3eplQmIdivdK
7wn3sb+pbgJf71yoXsUmHfg/BcACjRsjgwQovrRwP+j1xMpUsQQJHVOVbxs/jvqUwern3WSmeRpZ
OXuz8M78UA5nwyZIhE1ctsj87Y8U5L6RCBSt1C2aiwJoZcnthL+KbZh5sDAs9aWgEy42sDufuwwY
8caWYQ8bkolgu+Q/5aaMf+glnxlUZ+8z8SGl+JD5D3dsX4ijcnuvMxQ1qCL+plN1UJgZcLAUO8wM
htGKurj2CkqmSAdKS6ghOnp2nSsfpyuc0dRLoWklfxuEpUyq1M4mmUZU76Xb/Q1j6tjXGObthA3c
8xodBRaCFBanlCmA2a4+Hoqo4lB51n/a2RVfZ1Hs2n64t5KHSc2BauAlwTl2R/0UqpFL9e+YkNiE
mRLY4dXgsjjSZCmTEKUMq1UR9vZVkIOpqv1YM/HfVVQtroVQI1bxGWZqGiH5+7LGhhcnuULxa9MV
UAP8Uo57UC3+IyouCxiUbfsOALEN+ZhvN/vk8+yxl1v2ES+7wTVPn7I0D+gfLWPPB+J26U1qIyPL
nPBSbR8oPQBNmfyMEcQilgG5g2/UxGwKzpLtRyU5C6LZ9LwM9OeShx4zBszmjVuIdU89irvTq9E0
cfYBcTuBtaj8DHqiu8YrhUbizMaGWsd+c33tteJFxynvTtBHJ58uk6og+S2xNBttUiawngn7XI5N
ANn1QgXjxswuOTez+07nfaHPT/KvMVGxlzwWgWJ34MtCUIxzRC92wkMLOgnJzZnVtE3w7mE1O8cM
qLAUn7A8quLyRacIFNAr1ZRYj9ojvqAclUxbIYBqIMaYhNjv74SpHa8GbJjTfAcBzgFEdXuhx5DK
K0KCl9JBcGLw6+N4f1e/2ysF9F+CJBFffwVDTIjZmyIrJ9KIzjw3px1/a5t0iCtjaRi7zGf1riqD
pfEMTydFhiuZ7VwyttmDGHYeyjev6tgwC9MJk+YDMj0PlIuDTT/ysGfJBMkjDPvQrEZ/9zHcW6Lg
vqUEJIqgAV9a4eZtKBSPNyBwfLeMIc4/sC85l78HZKYLpDqaCQZGwT2Uj7QuaNZOLbG1BoqJCeEY
0PcamC/PrVFzJYrBWkchSDlTFkcZqNkpvUFNlNbKg9nj9q7vCmBF5UXigj+i8oIa1GfIwm7hTMiu
8Mitk9Gdf+yQ+0cxRXAGtGA8iDuByqnHqcjpcHZRl/11fCcfFAESAmCl6eFz8gW+u78DwZd9gItG
f4GSegTPARwADWV7cqFU0FO9TNhiwv55vlcIqTokIq1zlDY8RSCoD/VGmV7DoAOGIn6wyyX49WRo
cVcM/RMts3eWdR+ARzyTcelWBdBt4jlebV0oNkQvWr0vMif3b1xWR0cBeG1Do8x+Tc/3wcJN54Kd
raCHLWyznegdlH/Az21+TyUgDO2RUXL1d06vrjXtYrmSJBmT/gbtmJ1mYE7adILDvVAynvYMx8uy
5LeLV3emQp0MY+0vpOWeEerBXjDA9+9RVL6aEPXmt9gRe62ZjxKSqRuy+djsapLpA/m8KtTngD4u
ln1k4Kq+EhuSVMTdyWbEZ+CdxvH/w6F+0ua3d0dvcNNseyd6Cr2AZcOl88gFKJWJeNNAxpCX371p
CC049XlLKMVOLYzQ2uvv35iqeXa4u+Wv07WJ4xmBnuGInlKVc9XYhtRCamHxwiy189Q6jRK/HWY2
ePUB4RkSVm+YEa9emZaFGE3qMpIzCZqXx1M7aPmrHAXG6eX+PEgK/zENI3EKtA3YZcD7tV9IEysb
xIE2rdKBmz7LAClgz+lWYeCwHv3Dx7T33HUO+Iv0FbptI0tlYcXAiRxsgHlaqHrRO6h2qMW+ewUp
Yylu4DnAGzVWVY2DF0ccgje6w9H1LTmSRQuQecgNPPqkPqPeprW1s5vJB15XCqnZCuhuBeSMKuaj
7xaYEWzsRzPBs88qe6JuqIE8+PdNYyhi9u3LO6ak4J7P9gzfpWLXl7kkpAjkWy3p6Jg2vouRrcxI
7pWicMU2Moc8yJ5uLG33QL+vM0XeNvKXm/bB7oh7LxP2aknqEePB/P5mu65GTbnkmnl2RjnPEI8h
3gxLnC9ROA4RqMu69e+h0V9NruEQiMmnNh3MeRKL1uhXn5sTe49SyjbnZpi6/DX9xMPJadwYjnX7
y70Yq6Atyfm9Nx4QK9QkkXQv8SUJmBABNr2T83kss9PDAw0UI68S67t4NFjSiRR2P69qqxvjdJDb
LBgoeMBoOyWzKjjOcUPGrBFwdD5nEnuxb+GMnNJsBuH3clL+TZWXjxiXyRFvZvv8dcwFHh+q12f3
G/nWjdR9DE8OPlOHkhQfTm4hrbWgr6jFL2CKTDPTS18k02Qi1XcSlzR3zo0uWwKpfYW+Tggf4WE5
WQ21gMK5qScY6Gr7PVNo9xwxcLV1sBfC7d9ooXKHmOTuTTCz0Xy5MOG7AUAekR3cnWW5JAaDKKZB
AqOaYXyekgfJS8CS+EzA0yTWMcR21ZL6uFnIcje+x3nYk4DZwCtZveUw6d8zVVNUtY7/lMB5nRu+
vI3ESxV7HtBlQAWQ2cZAoGuVI2tvKlVkw5n6l64RyenoiuBl1Z82PbPCIBgRBFmkx4UZd5EXkozd
8+Rla2ZDIcGXT5hbt/ELG1oGTupbdwD7scit0Z5tOn5wO13usUyuLWL73veDtzNJdSDZRhtolpGs
l7SLgR9rfZ6ywmdtTp4otBDVpwGTnT5EP6ZJeneBH5nAhaphghi37AAKG5gQHui+Aogq4YiAgSe8
o7tdNjvkDjr6adni5Itn7UZxQtL01vW+SnlTAt6jjaNcAET7yunsgoMQlMc+gKt7ue7bIZuF+Dk+
qFeCGNgtUdgj8EL0lMBBEeGEuhsKiYFyFJWo8otoBlDZei/7Px4l4t+1xhscPER9FNL8rbsUqPeC
8i7D4JIo/d2pNOiGWdT3tsLpI34HnhB7JoKvJ97ENWhdBtlOIsBNB9hx71WauikdR+u+ynjzNDAo
kF8v1pbV1bY3p0gjUgViY0tEPIyGi4WKTglk0LB+o4EJKNGGMkSPwvLRIVCI90XRiyhqKXSejiMH
6Tg9nz9GAjZZ2BjEAoGaWRrT1CpL0PeIc6u8MU3dfphgxH05Fo938qjGU1nQJy/9cGswoFVW3eQY
580yCR6cDihEWReAOrEPuep4TkiWWuaGSqEzTBVtbDvKOTXC656TSrnK+kEDAS3rkCqZ98K37w2J
K5KKe+hN0fNwqryojJFYZfYnpT94eSpskdLXW90c3r/dRVtpusbo6mOFRmSCPuG+uwho206F9h94
+3v5hwLkOEyhhsezohR9w9J3S6p+rI0B83847x4LJ/HASxJGu1YHrwULNlMph0nRBvscvhetlRO/
4d+HRjKzsSp/x501H7Q6yg9q9/X7kxJ9ZJEY+7X8msufngI0ZaC9OBsnFxhrKJUOcJEe67xwjMGn
vtCD83A5SjX0gXPn3cHZwyP0ggtijAito2YKh/NOVCnU3wRf55FfOCV5DuOzd5t/Loc0H+o/j+AC
5j5l40i6TQ8dsGRfw/XS4/3EtxLeDlzlafujieGIYNBtVaZsg0oiHvmEADE1H+/2O3PxdA5KwMJ7
aJS3dSMAfczjdfiIg+ZeIjevbNmS/e+A//sw9llCs0qpfpYN0Kso5FQulEN9xUwRfkKzmd71S0Bc
R89zyz/VwVpVb25k57cpbxshS8oBkmsRAtR0tWb0QhQkJqisADNKwBVN4swxguHuaR6u8gN02nPG
wpVZMiy5DTQyfVlW+5ajOZcZuG6dE8ArSlfwikfNJ+r6o0eORWT+fp2xmyOB76DBDrYe4wc0msAH
bCVxUuSuiqNuRxWCpzUCyabnzGausrOVFK5Jtf5fcZcCBKbt6N7AvLlxG72KmC29fBlDZs/N1zYw
qHszmVFXyr2kM+HAEEewOHeie+VJdq75HVXiyGP59sYeKLI5tGrRrQJZ1QiUohjYkPD00w0fn2R9
QRJX9yB4HyT3oxOYNuDT8pl2QrM/eaLK1St+/9PWfGbtS0TYaVwu2cP532KTVPv6uPAkucj/7Qn+
A+AQiV6NckRw+3Cvnij5xuzWziDnX1qhcWwRbLyR4nbCVQqMKyhsfmby8RoSA401ti1Q9nqBDfKM
IRYvbMHrVkgnH2lWbzqeGAj0nYo0kY/DctN2XnLHVoLECoSaxk0OL6H34ZJvRPhx13i7rE5aIzJF
xfzK3lPKBT5Wp9+h3J9W7Ak8ub7dMBPGkarLV995A1GMCqJ8iCIAB7CfzXIMaIEecEiLGbFDNFYC
kG6cDm1tk0zFC2yXYvQcY4lltz+vgvELpLtdmPKSUnrSCPn1IokAIFXqai7YUqwtAukG3JnxrLM3
9dFyC3wnFJgMCxTSfz+/cPLKhKBMsCL/0Y31eytMkbcr9LvmUK2OK6ifB6eEcVsJWx/aT2hN+/hS
WOYPRYeThJBls5yk2Ht2YzVtxnUCPxy6D8UWz7zlziHFilx4bOEwq5GL0PGlaFvEIdb48ws+gPkQ
EJJj7LkqT6v4UFCAk/zFhHWqRKiEPJI14SP8/gtgiwTZh1zlDBIdXqD/WlKt4PKuUFs5G7lLgGJ7
iXirQ1oaoYJTmcKRbJGsWRu4acOSbtvHa2O3+cqO4xLSsVlvOHU1L+oXKokE9i0tPOGYoYvH7GCs
GX5c9Vm5q2+LZQIk4wTjmYHk6hFloZ9IfFDuQ3HoePO0H/cfEqGYOPKcdZEHGs3q8JEqxmGKEk+f
o0M/Id6l8eqlpK/pp4J5NB9OBoQNw0Dtaxzx5vh6jQPCMWqwohfoJJGjYgj2hkNOLoImtwfHOmWn
mgDT5CKXWSFYctZDrWbsbjyVR3neBeJ9t5PKdbgFUKFeigy69z4qZXDooS0ehc9aitsL6o4VshXw
CvW2rvZ484DmVDlijhurzjtgDYE8kfnePrCzMVsii3ue07U9o0v0TLu4ad0yq3QlBUicYNKV4AVl
qExSEoKkKQNd0e+Ch/DU10wBArvUn9HATlDlyMvIkD+zRU2jYXaEFmmGTyLEmAaEr2fDIQ09sRcq
tgNnsh5NLNaK/9VgQua1DD28m8yfYUQM6hRsf/QBi3+3I2+F1Qo4uplpM4WZXam7McwdiY/a63rS
HZ4JFU7hI5QoWMbjw+L2ATdUpSXlPhekcwQP/sW7y3FA0TyeNHSF/0DpHGdFP8xJu8gQzyN4nfHM
Us070GxL2w2xfsrFqDGU55PLvAgrMuRramYdKInVSoPfGTUswpd8sZlcthr3pndtAN3A1gk+wErx
3Naomtf3gPErU3rr3B9ZeZBa2DHZKatsFi9fuM7FcPfReyaUbWFBklvfFOMtvzUP+DdX4ovAeVco
DT9uzOGzZkh/qKr6O25m+TWRoT9KQkDTPeDmAAvg6WeJX3KGaDMbof5gK6c2mj4dFbsntUweEoQN
NY4qWynBHv3EpFc9FIGnV4rOP1pttNZgz7Y5h5HyPPU9YEpt1kMRBF35CLslW998YLYukr+NIVDy
spxgfP2KGLl0ib+wTipE/ZOxJDd6w2l6PauvODYAaTR7Ian3gb49ZQmsEg0/Ww9+gSSfzuYsGDa2
E+fmC5a17mTkjObX6VLGJgvUTDErC3boLQYsOBkrs0c1jrUSukESW6HqZgI3xyBbHa92Ld0F/hb9
HsufmREt80N9yJF1GiFBzZq7rWdAd2l8XiYn/zXEXrCiTocSyA0lhI+qxmWpaxFGPXcu61yi+55+
vtqnk4woTEGdLrhFngC/oLJQdqGPv/Gxx54QLezQg3iXP5/wV3LBZc7A/MPuMzYyFN/aeZ0k57w6
/GILO0HDJaJhO4sF9/kVeJL0GoW87zWMPM10MEvSwVVhtgwtH5+u9IlXPuEnhKE2Y0qOc+OzDpbt
bUcEjc5qJewZnKgf3cLom6XAnvh4zlXUR5V4owgOMRMRwrX/x9xMdqNRojnv5TFHqo5ehF4c8XG/
ksKqZg7a0rn/pM0QIX+KdnEynWEKLTOpiHfwrcGARtF7AVF4J6qX9A3BMtuUcKmbanPQdB35Pcb/
WHV6r+nzcmPQE/dWPEozLBrLBqj87JpTyQlE3wUiaURum+9m4PGf/PUGGzadH4qv5L80l/G1yQ+7
d+3we51hzKpB0G9ofYowgGFBBUWsgVceikoRKjOhFwtt39B22m4GIJ9WVSrk9NpNdkzmbRmiSDtg
UL1R7r+NymqG8XhnOB6nPinjmgramqg1/VS7/QGEogMlqiTHI+OhJj1VAi8JVoAwR1zzAFwN6s6W
nz/ygHYhVUcZsUVuEwvHv7kyMDAXoLUQq0PgPdh4YDINPi78A8K0L0jGJu1bB9ETX11ZDg+pxI+g
729Z6EUUNVHMKAk69BkGFG3gqUcRVV2K+x8Kx3DToSSo2UzGdEzFP9yy3ixc/EgjhrkCKbX6HHrA
4zI8jcCID5MGK8lvL/5oaWRtkSY8QS+y4VaPYv0TXefhn5EI2Yig+5apO5UH5bnAh38c979dYbU3
MZHoECpsFj4DIlG+RJq81hTuA1Y7ZFLaww4FRAz/NXnWLWkOxunowRYNy0JnmNietfhNReJWTRfO
SyA69k8wW9/u/gH+qAVUeC/YE6Fb/8QaulXKKEiV7M7HGDoYdysmhyexNhRE+18gn5e22y0L8Ag2
jQFnChaCDABiAC70pzNKGg63lscyD8Dx2JJhGd5NN9WHogNop7uvUkeVC6nUnIjTwEREt2ZxDhY6
Hi77+Gvirv63M4jpr5ZHyQpfDabPfP2HZpmHfzEZvtzCKu1qbZad0uWCXA4++dHF8UEYADE8NXJ1
XXkjyZAacomd/FJIbOf0sY7iRu6v+oK2iEjEfaUcqW3PVP6I/3V0lRtLs3k3Qxi7y6mn6Q7WRcTH
8EGrkLADcWZfFaXSLqdJchCJ9SEfnnjkseLRPdl0fNhPhLXM/Iq8MKTSuQ7dWQWWy9Wt45MAvujv
YTjKo8tVVL2B7MohezCWHmynZZWML+ZaPSEUXkfBe2zysaevsKFG+tcAEzdxveZ2eT4EgsAqeOwV
uhGCz4c75PUuXo6TGb291tSTc89wPaCPVYBgw/1D1GcbnErbOkg0eNkZANT4SY+f87XrpBIvmkP6
kgzLPJo8SrM3A8JwIDiiGj8Tip6oVUg9MoQU7FqxQZVXUIubQQLGi5FW/5Fw6pjRKmR67J58DjIC
imGdb8T1rt7arD2KTOQkgjF3/opwe08qsGl0otRhIzoKh7TZGiw8vJ47VSxkJI5dvEVY0XKY1rbB
OxdWlSJ9wFgw01lnT5SIosdfpjWhu5n2rC/VSk1EproSlx+CJslqLQFk+GQZepomtovKt8xXzrXL
JxD0Zj+02C8WU5i9VWZO/ssabGiNKUlLNdRDw9SrL0oGiqg0WhijzOqAnsGaOHgl6nyHNbaMX8hC
yEIvn+tzEsVQ2TWu6ifBgqxgx9vlLCaB/zOrYKHGZm+pWLCgn8BSbPLm6AgNyTwVETnGenDXPnWg
dRxcmd7K5EumB6Nj8Ad0wtYEkwvIQoED6TMIDaV1ORR/8HBC8nSOgEAmfaaf3R1KD7X/8o65u/J4
JYDmIGEnxrupPN2Sulfin9+6iBmsa9di38lBD2S1bYclSuRpdkhM7Nkyyb04Lzfi1IqhMYmFLurY
Zii57CP8vbW7dA869ewuNNuTkqnasEvAOTvkOgMYA2oQV2fhztENG/hILaBI1gg/Pa6AoW1CwzL5
hGf0KOS3UnPNgvZHkbqX2KdU2qN/54Qru8Kh/mXhJ4kIL0Kis6VZQ41etGVemvIt9VGBqTYbeI0r
p0LckKTtCnG0/g7n06719GMzxpMdl/Vr4t3rManUWxJ+aAu2VX7hOOqMKhPacYazHP1MA4B8rHNE
uNY9oPNLS0lsmPi5MNfzsCesZa/CMnBPVlYJ5wuuNPbyQQGL78GuK91AQ3HlTETCdHRoznhMwR0Q
4UmbzfpSTk97YnQJqgqOqCAOygRnWpuGMsOfCR5DIT8h1kQtsMjBeBhwLWUxqLlKOTZ+j+y3RSF2
jFeop1ISI0kX/INZmRj0MbywS+qklNwq7TO27MUCS67+NyCtWvcImg4xArlX9r5PkOIB2hs9z3iq
x9QaAsEkNEVfiPRVCuPZ/3YppzlR6TRNh5aX9rK32pjuPLXSwPHzXA/0B6Ktt0wGy1JXmKZZ1WpZ
VRIARE5dknMknFAqQI6K2STdMO90HSHLilumdgp7lg3gaZ1oLvhaxQmfziLS4W1OwTnxvqMlfsfB
hTNyci2Pa/MKslLpyLd5PXnto8+UKz3VBWOS8+te21pbhw0e7ixSk92xIosRoT4VESdduhAIcKGQ
SvO7WIWKxWA6Nr42A2OiynWaj+yTI/BQaCasssoLTjgANcKRD9t+mVVdW0t7N8AlR5/IKrnCZDnB
k2X5EbsJQTMD2bVL3/UYL6QcJrMAHJcVcP4QEdl0DMW0M2BOqa69QgNM8GYsrFdoZBxQqemU3UZl
4qoWG4skAbYz7NjFQZ2/reSfdM+k+Wzw+MwLEZKhfYqlWqWpOU598eKbOYrsfNTQ6EeLBt+UxxDv
qEXaCmQtAefyXQkm/sMgoMCgTv1y82TN48TMSR7yqtZIY3i5GgNpjzYJS4Kx/QXVUWzLpofRrAP9
EhqM18pcQj/EfgalAlSOvGBg2UFRz510WLSfcYDYccOtWMbPv8+qwjystHSYg2fZUGwjhU1o/4RN
GNBjITMOPc5p6Bky4z5tp/DicE0jX4eJbtVDI2zHJw84zxkqAg5FQOkxMVQHhXEP79BLuiSx4Fbf
CXJhJG6gT+cREpMWV6TEs7wW/Zk6WOUA1ArRvHctXt2P+iQTohj9VdHJGKFrgXeVqWbe5nT2510i
JQBCT0N1GgHhNgBdXpTBasJdWRQS7z49QMQbpI2DzivrDVsxt3k52t0xytjaIJPr3r/w5Lgw1MhO
M8KY0b3Y/o41g9tSa3+OCrSPB+kAMz89yXMskDDnpWz8IRQV237Gi3O20bsf0qjE+SWCopfsJR6u
oI4JnLXoVf2mTrabBr7POTmS91ncm3P4R92/RNjZaSfvEdZO71EEaGqQpz0Up9rJ7w/U8yVlqk9J
QFxvYv1BF8u8cyIpfvMyyIGuA31jafnABDDEtgt7KsXHh3+/FDiKW6cy64TDJpfeYjCFzh8XTKLC
0Qb01+n3CGoR4VwgpkOJ9u4Cn6ABlOzjKOJ4jA4kC2GVbUPRAJbeJIW4qLxlbQRwg2qU7aLCPYDf
PbKn6Ui+suEohfBT8AowNnYMy+PEFzwhO69Z9Y0nJXCZUNm/7uNPBXU3VOG3viOJ/bjjbb6je5ir
4l7RbRNFewR2FFOoILw7rLr/sx1gcSAsL9qF5+nSZ3dPGzeFc5hq9sfNuvJC1p2DQwX2RoOgNvyc
EX/QbG5SasBcx7WqPN9799A/qzKqPEcpIbWaLlN9eoE3EbdzRJXEoRUwEIE7igVgowVgQs5OwYB+
gm7u53J6KFOnK+f2uRzbFESKiMJsxignvAuMcQPYQfntqjrg4TQr7E8CiO2gUBkcJlgxfFWlOaRo
Tj2rbnrV8Kt2lI7+dlhYmZ/WDMiaZU41RjNCinbFAH7zRV8q3Kwdn/NA10wNQ9ZF/fX+1TYy0Z2W
Gb9xa8hvNYXkCYDhbJE+hM9uTu+iqZgFKwxa5gYKnVZWsk3WRlKhyqPrnPXPDM3jm4OQ08n1ht6u
EpCdzr+k3UcgNPYuyLIUR1bGLzjNwbEZVK0XPj0md0LvwmUH6fngJM6ECdxLPDcR4CbHGgOEA373
J3eBoVkvyIHwftzq4F2xhLwpggUe9GoOR/rPW2YBzhTxL/IO3V9qZS36SmPgR8H5rk/T6MlES0dc
3c2KtaR1KuEYD8URxK8S1q55QKbtW2tWf7DR0CnLD9T/O92FZeqsgRpZJIHGknBTAcOfnUjIkQtd
MF2xeaYdjpemwX4Rxn+g3gNuQtXuo3L4FARvLJE4ASzC2JmTplAXWxa+MkiMuKlnCO4MB/ylUtr9
7DHWgOrh41leY8skUSi9RlIWyGpMN4gkxzx/2lxpnZbl8vpYyaP+SncZcapWvpG6fbXqxPN+Upgw
iWgOmK2365SERc/jIczksipTpZ7ZMit0ibPGf9HwRXcOejdtVRbiq5HzrBUY4AqRCsm6ELTHnePA
TIFgTYzAYsiu0HYG2LkLtFCdn30VuLAm3VtGzC3leRyQNx1m+OY9dHZKJG3Am4Vwo88MhXkoL/lV
LSwPAqOLOEs9d27v1HSZySIx0HgtwQHeCUkXSPYcTNjaUucsiYtjy50k++3tPMMvjq7opeB4ztZF
vBtOPM95vfTZfS8mb63ggXh/9kezq7oJHTBcHRyYi5YZBffg5RJxSA9/VdQ/dNB0w2Kgk2zrzYnx
aImOzBch5BhvHGr228qkJ6mBA0ub6szFVaHnp5K9psSyWxhIlIw6zSYQQ9Hw3KVKStQqV1VRA1jx
l7ZUFI8rR8kCmlMiQEWklkV0vrO31WAO2k6lYmB4DlLUs2Q1c52I8lq2RwSMKqbOy5cb2X0vcyOp
hqFb+0qPlsnD3DtzAotM7g/KjEf+SQ36cCin+jAcej7/qHKccT3Ws4TPYBfdEIJoJrtIC6MVf6JQ
PytGDR6CGjy9p2U/YLL7YV6AtPccWryf4Zn6be47074jOYJaoNaeqd+BMDkO4RhbAJkWOrn9onL9
raVtsMB7aXUBQix6nMg0NcQ6OvnjLVcdLiA94YoyhTPo1aAU+9yn1VriEJw0qQJOyE9+hfVr3HtK
DAl1t871tGCNyV7MwR46aR5h3NNpQZxrnhp6A8XKHjBbA7hh0KaY8RcmxFDtZ+4pV1y9xPClfEzB
j6Z3LwXFnCzc1SJtH+k3x3bVLFtivfMLlAPfnjijtS1TC7dvgmKuRSTDvqHEa/L8VHcd8BrQ3G0V
TYElpM5J6Mv7MAqJVFX1dAZr7svZxGZ0KeK9Q83Gzpz3iX3LkvOg0tMsFRl4m2kLQa3OaGSHDaGB
lrqu0CAYDScqZfeZ7j6tc5WAonLh4sZuljsG5txqyiLg+Waa063O5fvAyhD3+pl6/AFrj4SbAcQS
YPTUMqykg/IwJ82mV18OOyQZXvMzO6ACVdIMrd+374pG/HQRLaFB27ksqg5WrKcSR76X4+VXYDPk
QKfj+ZehG7qquFz30Lc/lOPEdvfVufqZEt0CuZhPvDKxBO5AXQdwksXLrJoSGt1jD8FSeANG0RnD
coyzZS+9BYPcQkrreCQ/1gW2hhpfwYfZsm4gWZg5EFo03hMUCjZlu4cG/7jEYf1JSVJmraq0HIqc
jG13vSmwVPKB9RnSQPe+2p/S6vrRYKm6ZW8A/TLs42M7PHmqHbPFDIsJNCrPjjQcuqFpEaLCpoMY
9k8pmHDjj1MNFknQGdNjVQD8dFz1yHj54zDZRyeJArtjMmhw1mxAQyy+RVaPOGtIbV6TWq8Khw2T
YbuKmclsKX4JLjgAiwkzvNf5PYb5gjh8vGBevwgqDioW4Q6oMPAhXLfBHn93gsmyZch5e+LfZGPY
9zZxoI3npsA4VFhWPTcU2hL1n2z17ppmm6i5tuJeGrP9ppU5VCv2UjBq4juNduEtQ0okdx47bWJR
sga+P8WQi3iaZCHlWinlYPSkeCuIIaUJcCRNuax0J4+gWwjpPl1gdcC/IhwIz7KRMYGtb6nC9oWj
nrcCGy7ntEufHHYJSUakcrDMhJyJ6BJlRNAEgR38yvDAuim8mXawtHp0F06haZTpkas/LbTGiJL5
8rwkzdTjGR4Ce/jmsQSf5Yv7o3JQ8VDr1vAJJlYbEQgbJ4ElJd6xJevfLkSvuSmusCFaGlRlDPWF
ageNi6nM/PH9WErdyKerlOzPpWETj25hp1k4/ntgyDOKrugtdDHvPwNjHE8DZyKpPTZeVEkx6xqS
xE7Ls1DxkCMMa6M+fXZHcFtk6NS+hw8mrTBxb1VT6OpEfw+/CLcaLQyEPcgiHPQ3oF65qruiUN6B
oqio/zohZfsdTnNVJ+PXaKAGpcjGth/JnEc/ey+cNuotU0omPAmw9+kjDiSAQ0TM7simpt9yErd3
aPyhgKdQJ/wDyLq+aCSLVX/YSoO1Vv/OXhxfcR6hxPBNLhL+TeDYrGJr3j5co4MDWwQxKBRF6eqL
1PaVw7L2IIC9tmab/vXG/sdb85NtCapf817AhO1Mp31Ur8K6Osq6J9Yfaq4MwD79mCTdFC14q+7T
NIXeO9mPoKny+WpnU1hgExryZ/dmNKp6VqjrWLMtOVB7n110j+K85ujVEkz0rABAVXqj6nRNVfAU
z3IxdDqNYxLYFlXqVmTNh5nSz8DbB+E59rKUE66bicg7McaXEArEpXmBgmujiGS8vZuI77CwK/8K
XUM2cXd4MbfaxCjZtq+0NDqVrrV0DY5/WO/BjJnUP9BTOejFe+Wn08Gdeq9FaB6oyzUqLFq2tNXi
uLMoYRgh2IbsYSDJaegZt/9Z6gTBYpHWmPoc956XRztPflXQRC43J6zTlB0DPDaruEmf++Epnm8Y
dwh5DP8IqfycTdjZ+xDXKd4fSlQdmNt06/bUkbJLEDRmGlUkU0hDWN8sx2zXh4wct+hiUPj7ncTv
uXZAqOuN/YIytD+2Xy6xIC8py533TkB10LgfT7IoOjbW0AoWN844lCRq71knrYTlVMPZkiFwG9cE
hqHxV33LpwPm8oESct6yPVcjEJLJSN876sS0aQHb9KO6jTtkw6nzLhJX1T3nNjX0q4B15vB5gZXD
0XSDvrK3RR1Nwu5fKlEM8i/HLbWhZkxynHCzGrb6r+1d0ksft4RElJJT6VxaFbd51RWVKWQKBvp/
4wxMPnMY1xRN3DO6M7+qKlhyA8Ak/Bqne03R5P+9okmoi94dZWk4a5gJY0FbBZq/bsbhG/6/r8li
kwydb7gDx6Pq3q6qv6BI2hLJW4j9BOM94XFKBgxBFck5Ivn8F+B31JfCqlYJpRSPmXCLcNjoQxNt
1VyThzIVGMuZriIEdVNjvZYOhz25i2luPVRPXK7XF+kfN1sK0HUf/PvoWuQjSP7Ye9GaanCKAZs2
B7cQAcCLKVeW09ZPEqstpDe7LCXinACMJ3PxOpYy2y3FMkX2/kvr2hdZNfoky67jQCCaexiMGuuO
6X9lKbTnwb90l1vzi394UjyDac5loTCcRVwManRwSU5TNZTYnobTLldu4T3+0QJ8llCoG2FHTpJI
LRIao/UU6JxCc9bJaf16XhG7A+B2brwouZoHF0SANVymYUXIZGE1dXUAlC+35YoY1XelNKGoHW0A
ey5dygkjOUMDB8ACeBhpqDxz9j5isS/meMofmxLZLXY0+hWr7lsceHx9NepwoIMTv6sGGfRfEO62
M3eUhy4XW65AE+zqLeB36njBxXNvugB7BhDdpV1qN/ZyVSQ6MoDFp/H+oRCE5Kdb3YKyRX1DCv4P
lAkrFcd0J+STZS7f3QTgD6uLAlVWpyQoXXBYGKba6ekhXH+vEtkYpdD0+5FVyETRLi4e47ddmep7
BMSU3aFz81p0EV6AltmnTjxKfJQmmq9vAQsEQEujIhFpWsckucafGUjPuLcajh6uqRDgpSmJW7Qu
aifjPa7xuHwZpQix4N+kuPo/l7/Ca1u3Hd1SG0UA924wxYbsc0PLSYt6LN+P/kuse/I+3vELNGrB
KA84DO6+2LQO5zy8XCZjgaSAoNH/F1JGZhLlda0YUplFZgkSpRqXGUJs6pBgCVDaFxd4QXogSNxW
JaoJY4LUNMvnSeMiMH8X8BugP341CC7Z3/+k3WbUHmjgqRF9f4qyJEFfQk+ld3f1GnC4quQ5/yfD
YZIOw4xAVSfBhsZATpTCIbHq1lj85C1cJjBfzZTiWf8AwDZ+M8JizR7LzQ01JmBxCwbe7mEjivh7
RvH4t0PU4zD9zR2XuqKx9ZVS3YwPo9na6cnsrcSUr2f7VsoldW1kxFQFfp+4OoU4rPMPfFhwd+m/
ORsBcRR+K2BYOk3vM6BXq2mPq98TFCQpkES+kgD1kJ1gpsxmvAviA7CwgOr8mPVrXm5K8/SMnKjK
eEBbv9imf663MeFsEBC2O1poJRB7otQ62UvPmd4/pvgXB71q/2hPPId6AY5f7c4K5tLKkj0x3m/X
abFBxhGrqsdxvM+AJcrYdk9GG2Nx6p8ldPoMHE0RNdoZEmIK7BULO0LmpfhfqLMCisD+bVgVMgob
0oGLYDiS5Pb8iR3cTVFNNn41Y81NG56ppgW9OnQ67MqM4dcYxtkyOZonyPyxkg3YR7wahjKmp8BL
+JZHDpVUcE3bDOpnGuBxQFWIszRsNfVWxvdjTO2oRqIS/uq3r2Z9GHNCl2Sw9A4sXqm0sUzeqy/e
nS04dluyjI2BlcN7pYvUqyGjVvZcBx/hooiT/G3gM4hjdBS5fliU1L65QCnyIl6tSld9aXqg+8lr
riRyb7g7pA/CO0a/Cn/IDQjy6Z7hBnxrrBztXHkvf2gfVSGW1amZd0oQYBOla1rPxU710CI5JL5G
2lFqpNJWcW/bytXOY6JytNm4JlIF8FLn3uJy8ECSRK+kY8rzgU7zxk/TlT6J7VU41R459pGHqLmd
aroXHOkqS0mxDDD5vlRGTKWlgCAWGuiP+c8ObgjzVXq8OithiY7EV4aNVWQdWycLmSz73nLHTqDk
7Dj6mSfwkI4vb0lG4cyfGRYhNZ/LnjQH3CkAnu7o3lcpwU/AndUcKv8XZQCXrlTF4aA/knJBoLtI
qleGmBHF8GOMxxUe6LvlF4/l7t+rAJoPpOV2FbFzMFzJJ1MLKhmrxUJmbb9JovnidR+VdRnfmk+Y
7ijUY4AM9D2HX4o+Pkmzt3Gw7WuM/fVez8fzNJ9RlQNlsoWNg1pmnDHzvtw/y6fcDoU4iT5eSERa
Zv9GIzFcRT/LqWFKGwfpgsn5aciH34w3E5WCqTBrhdNDRqFZcfVNmY2ZWJE/3hedUVnmhORBONDA
86mNX+62QjHzILAvouRcjXuFqF6e5sZCGMInSgjlWf0hCnPc8vn6SiAjNLGbl/zZqP+l2ezkHZss
lQ8tH4pIFpAWlsLYEBeIfrrAcabfkPTl1tZ/tfhap/1+mEjZyJt5UmHSAP7ZM6IPKi9WJUKXUTPj
BVCO5K+VhGQNAnBsG5TUYwhhoQgJ99xkII1/T8dgWLNSLMniLQkp1uJ7L0B33j5Bw32HtZ6FmM2e
K/KnZ8VJ4QlD7ygK11H74ZBFpBHGeDim1Oy8ggEUpDIFK7cKY8BL3nFGFA5ibmjUNr1gqtLPb4Yb
ZO/Gam9d7XPNbIgCYeEmTuOK7GwrxwHN2ONZ8OC7Ra3vKnVcqLKbALsdiX92qKxkAW+BVgSZrhN0
neLyH8/HoSxb1F2rx/zhoB3tYnqTBK4QcYEjKxzmZtS6hMHFmjn45m+axZMAhYDNmaVeFiVwSQ2/
06LGcPNTfhG6suoAzRMDKBEt4hgC1LBi3ZtBl5aORyOK3Wc2xe8cNkk1oqHYpVJpf5EhaZEoAlij
i6Bb+/VKK3ib8VvGvVPJax1L36y94yVpT6i8U1fLUSVb9L/flQk1fUujJipsgv0TUOLWlaB1WXkg
/tsEdhWuEx4tBpTbARFnvZppShYpS9AdgD9OBmAQ7j3oK/h/CiyNTsyvrmxCE8hi1noorHEpEOIS
ZJ9FDisj8vk2r81UA8+yW4UBKTVBquNHLZwY6htAeoP+ckRw9w3+EFGBZG47NGutGM+nrDEl1pzl
f4uGZewkPUJWHx4x3BkK5aNqw/RrDIKd4TdPdjh3O7S2SHXXdZw2xPX0cu8AfNQjyJ3rmJszGtBF
5K+oQDJdo1tzLwzNFWuKlFLUljwFKPOw1eZbEJJt667xh/fcrKEXHNdKep3gX8RLz+al3Lg12Eoy
YOKSdcTY1u5gOUi9IWJbP0B8JAQhPsa0NFZVuJHuOicYikzraJQWH3NieC2P122nsIVlr0LxeTxi
XKlHcd0BpF+G01h6LvnBAOkZuQse0Lg8mtlkP+9udIZs52+jJDV36NEz1H8/XcBkMG5JuXbDvZx4
VOXnh5ZVvxR7ddMeBwBwOwAITPA8wiTxRD0v6NZdrkow+t1CO8+pRb/1L4cWdTf68RW+koG9H/5n
/VXyM5joFZvteaANRfSKOSpJBiVFtpwSwVHFPvyB/s246xpSuaDj6o1gXK9CVFpC7PYptltk27OH
sSVdR3yPrGQqpTuYAi9zz5O4tA98vNoK5FnnQNENRNMy7hCEfYqr0vaVU+d+gxrP3kX7yc2nSfxL
ip+2habaKtA9bumSQ6+tfpp2pBnoBSbe6vtDZEjA12+3TgYBs4GLzgpneybZrDJYK5zRT459zijU
T6mragGRjnaDW5R27jChPbEQubqoI/xBpiCZq9e60+dyPJr0kOHeOStsz3DWoD4i9Foa43re+l28
g77Yg9LELRWCiORlN0S5sy/ah2oIGszuuNhkitqYf78naSIjTsHwYazf5JB30ZSZ6HAllRJzoQsT
4z5wyYUSfHlabJ8oaIu8RYFhdYwyxBtG54q7gLyDWVDbRtXg6UdeQa8NUSUprkXED+24CzxpZx2U
Uz2roi5AZouAcQLqQ9TyStXbxnD1GhKS6VGdo0wsRNSW97Zfn9mnDNHHRU/ahgAtsSSankPICCko
S2YD7qb95N+al44xwzB6kc53O9erILzhbg+I/OcDlG9x3J0lsx0+laBesSD2WLrImVY/PHtU1rax
Bsb/jM+ofJ4fJ9aD1C/o9VkMeYuy6ceCYy3JX2jJYHSDYULwl+oP/tXnfh9BM1u54fCsNC8Khkq1
hHu9E5DXW52co7mpf9DywZsuEDFNryTI4jKtVXdkyBrymiMmPwkCwNdT5btYM60fL4tsFiu2Bcop
Sgo0BfVjDOdQVjNt8mIlUS0SYIXlhjCOun6NPuONd5PmTxnbwUGrw0+EjBbtSKuGDncAOLM0dUHj
a1pIgRJTRTy0fLdyQGwcO3mYjIDig9Pp1ot5rqSeDvHmCyivisL6oQAfzlNzF5dgoBUQe2tMpfdr
vLMER4VveCd8e/mmYVU4tE2qNXpyQIWc+T4dF5MRTBEXZr2imGg1cy6hACjbQ4icPuA3aHT6CXFe
u55JgWOjYI3TfYvKghbUGIK2ACuKs7BXv3bqrEtjGWbaQezjE02AqY5koJ6WKTUTsBoEfsSAi9Bg
Eq+0uWIJuaVCKwfzVrekC0GFABEfz4WkXNZMKGv/wuxmzmiAINfpO9bg+W5fDBGWEorftTnJsjy/
z88mJWq4F7oyoRd4k3zvDBs0qfFPwNZn+7iVxhw9lOaTWRRJQ2Khl3hEiWTXkHCFDfBpMpBO5DBU
jkSzhwvVpNCxCrg2aRtYAZl4jjW60CCMKxJBGxt+TM3cbRccNmO3UU0HcXPD01NlEGfPKwbNTBqw
4zf69LOhrrM4/qUOqyShoo7oUyiVaGjFgCqZABlQllLBMd0KYGZJ8/327YF554eICtN1ErDdrlJH
QcykuJztKp5G8Bsm3683kUME5WSiPIdp73eAxfRBBo3+RezH1ov5FY73eF293H8IKNgF0dvKA98W
k/0KE6TrPfjNqIt0pVf3VnZSEvCI6e9rSMkHrywnAowJRjtft+8TkKfth+Wq67tSey+bmcQ29hkl
2jr+c6CyVMD6kpEOqdxKV2zC+sZzOetjtEE+QeedD70h8iG+sV4ThO8BkyQMBiarhgxNtoneomPt
P1q+MTjS7d8dzewCtfgmef2NZe/NSqHHOwJVK3dIpdWZl/Lq0CGRIiqGITgsa/nErKdnpo9Ey3z9
5eYf17+jSjLtl9GuStP7yyJmIGvp4x7cgRBq1ywO9pDkUhDdb8QfeAblfuxnuQdFFMabWYq9M/Ns
XKssgqTuTM9R5BKddZAH7XeDCi9BsXlEVrOyEsEcKgBpR3AnAMv1eTbHJN/0GZDxDqJE9td1wS9k
e17+q+JxpP69OVg7VKcioP9B2Zum9vDj6oektXU9exOfUCCUmUQcuLzw3kIgKfPM+fZBPTQBiN6N
Nto/hezmdeU4wyy9Bu4vBqeQbULVJ1pBxn1Vm7FhkW3tyceDrybYQ2MI7+KyS0/7OZwFbBgW2hcP
CADt9Gz4uvh/sC9hdeD674/ZFrAN1WGhunDj/jN5+pfHhMmEHNsIyZBLS3hCcpxn+7XWU59D/ADc
APbc8EM0bjoeTn5srcwiU0ORzTiM08Tlr0g50GpWdRUnKDjwFwH889z/ngGH+1tjWSR/d5raDwFg
qfKVhZeddUnNzEulEEN7u2ZcBaoWoHsSyfJCEvuXo42OubMtfQamzsOC8K9PCexxg+e41qOO1GtE
TvN0cIJxCtAwMZkq1rznzI6a9o/zBqUdD4JPBhUwx5CjemegmgWCTrNSHfxA/0B/BEUNpMwNXVca
N1Ro8MOo93rQzPP2kUmWfiwbQZcKdRxXrc90cb0E0oXkXPWn27zL6D4VegjzLPsH0e0CPGIYB4eM
RhGeJGKVRcP86LKruIutti7WXJh0WAnDvbbrqxGwrY6s6aA5Nyq1uVnDyUZGKE4lEUqxGmg0Q1z+
EAP7D7ICKAuhzi/8U1bMRjgpyast8L0BVFRSxEDmCGD0d+8A0FFKxPGIizJ6YxFYWP2c5gtpuqXk
AthAS6SaAeYNs/spstkA6Qb2NtJQ0gnBhgXcULdILQo5oekjtrZKMDBIZfYjc8W5hObyscYLwQNQ
wJ2AE2AAatE+V8193DTeJlFBfkzL9LC5JO1FDpAgHdyPxGK1KiIPcoCFgXLLfRGYcEQkxxS6r5za
J8ieBpmfG4qBIddNMf548OWLu3CpKzns/11gEDF8qYg3sDbBTbL8QfgvpDmbc1WRvmZ5IeK4PIA1
wyIkT6d9bgDvyREemFTNuGlGxa6+1jaUInwZ1H+TCvO7LDtP73zWfXaOquntYC9S1NvDfoM2sxdK
Aj7h2LErWPPh3ZTja2I2A5aS4ZcyYL6eAqaw+G28z7KUCobkX0nZiVwkhpFhnukT0r2EhGM+WMOS
hFMaltRK8gxbTTP5n+h7PhU7vBXhJ2ZGso4HS8zrv99HDUaw2/llIA3blt/Ru5uKSQBkMOrz8i39
yq6sF08yMiDYqGBeqvzsoOalurcKyw4t/WaRw94UxKEM2xLbSaQmgwlfFIHviUi9Ac9+qfqJJ+8d
gueM/ieG3Qde7bJz1bYoJtRFWULtN7sA9+Q9PEsx6o73z0X8VcFA76RybP3Dt7gKm2EqGRrWH6Rq
lB2/2ksqvtIeIZXOunMlpdwYNflWreCk/0RLT483579FCwJ81pCjnTjH8R7FlUDDXgfgt5pn/zv/
kJYckbB+Kno0cwGGyW9nlo9p8irANHrbkh7Rj9j0wasfuhbDgrRQF/1x5HGB/aVj7idpQsVXMjp8
99hbLYHSYi91A1IkjkgSJy548UnRGVJF+fMkYDviT/b9reL+o0tCR9129ZFUc4Y8mViwycblIAUu
P0p3tjz2fF85TM650YkrqylHx3E70x2JVEcoy0Dj+koRZaraYF0R7h/Blatp6MLczK/AHsU+gssW
Jc/UoY4ffrLiox3MOgOTvcCjqsiTWU0dJDcmceSkvUSEAhbWtzeIVv30fVXAIhEbTwvvFr6O5jTE
72qQG7SDh6+I8aqXRkJuYf/fMJ4XZp4Xg8aWd/2Bc+OaD9Ktb9e2mKwWS2CjfBkDkzjhEj7XfKhF
UTS8D05ahdhkGNPmfwWkKFlWTa3SpTG37oYhyqp0Nlb+jH9zlwafFnf4Ln3FF1qTwgvU0dQPmDcc
+WFO0tNHmyCxbojrzQmJ6Vta1wSrpxZz9Zet+xZAQVvlhySAYLk3L7jkj3RlqFb3F1DS0GA2xORL
rHk4uwUlSYRop/Awds9KxB+/PiU4Y72NDRCALQxVnMDMJvgYhopv2UuVrszGkEc7bbxybskk2eo8
1m82qDNLDCJ9oPBlX6Oot14Ou1PqQH9Z7sjCvtoXw8sAjkv/5/jUcQdJKAQuukwF18djNMar8f2l
4rYwifff7P1HDHszOe7DewIgjBe8I3dPZj93P7ipxWx1YWWpOgM83Tbuk5JbJ2Eu1myD2Xb55UFV
IwNkTY/G4skNDlDaB+ur4kVUXhfjxZ8oMk4NZtq0lo6jYYIszUXk9fxnIUJfMPdbd/H568LLLqQY
Kv6K7zicIcId4HvgUZbuF2I5Uk22L5wDGhKmKR6v/duOpFNfk4aDeNnx8c7qsY7iDeqa2m1HM8uE
HPx/zkRW3GmyaSfBDps9BzTHtY7LjJr9IX10htHUhRx9eVoqjpp6hYy67qsJ0KqvLfeOFQGqUVNM
DYuf28hXk9KRMcq9L/91r672YTNlaDZWnygCGGY1dkAsZjEwxFLAJKpe47/7tAX6xh0slIt4t5fV
6BEHQOGSl+TZ7ppPDR97HeMhoGc9vQ7MyrodgdLKC8ycHDarop1bn6wkg5am7IddGIZ7fbxRxn0O
OT6RRS/pDZ0crmPGkXP1T8R7vpOoGWPHjrKH4QvWAsajbXefR3YWe/5lBswfHg33fKmpzKFelCyf
8w/TFuk/JU4Aw7EfK2tIBJOjSZ4cFMfN5cvQJS8GG/OQzMQ/DF/QbHRLfdqPUNqXl4VjCi6PFO2P
iYfq2YxSIbqxHyiLg65hRh5E3Nr2pRixk6ML/DgiXFG3UAVsai4gNqpgsbDdU26A7BXCYjVF1hdG
UkusBxdxJFmfFtS6l9abXfLS/QsYk/vu2qppEYQRsR5P8CPBhdHexIxvPyvegxWyHFh1+p+JlzHv
Xn52mkOc40N66O/+OuugH8n6Di423/3eLRLkXpiz9HK+FhD/KsP4896RL6V2/qoVdG50aKGLXhNB
gT2PIV6UDiAW4iZU6BfzeHfTPDVaXG5/ko7QPZWePD0tdpA0kJNo6C9bofIFSrrLyCX1Y45r2c+L
jyr8MX1p18zVvjhL5sBRFl0BPA6bFcrvIH/0Xv36vnKhxpv3f0dVrFNdp+3xoRhvypT0GD7rDqcE
/nN2ccd/5wg49xyUsNHx6vxEKCfKJyYxNrXNlbCI37rzZT5LMQbTUCXH6BO4jZ/gKJSRzFujLAy7
D2KM3vD7Kexspao/CP0wzsboRCg7fnWn3zguurnyeEh317xiczhVV2oiiLiddNBEwMQu26gCLUdE
46WD9HjoVKFPKc5H1OFuFSmFgxSfqwgQhvlqAe/hm6WciqAAp5okSj7T4+2/8xLDp0NRzhmPpVQk
bySGfqgsY45XL1sUXqmXjnif+en1zkMOeFw2URprkENg+lvCQOh3JtHA6uLRe3iJcRqz4Q1dH1WZ
VfS1OUzwEV7HzD87iU9+gnZMDR6OjUhQ3j2jMh353EjkWqjDAz7FB5Bn3a9TjquN7QVXChTeTGXS
P1fvp9seEdpPgQ507eDFKdLd/q/jENq9C/zBLParTQZC0mMdPQSi9gM8npfrRile0DBIqims59h+
QhzsMRWfHAzmYCWJp3QP6k0aGhl6b/zxr2s+s9CaWI3rQQwHeuvbAOPI3Acnu5G6bdDR4FyVYt8Q
Go8f5i331SeewvtkMMLLgH9MBHCDmzTj/1rhKJ7gHsh3qzk+V9QOLFTHd3OtgZq8e0kbaOO47Y4u
3SKgB+XCVPRSHs7rvtDT/lpBX6bpvLlWVcYhh/cy3uUc9K26enSYvNc5mrznsdWHe2KLGc3P0LtW
fB3QRWFT94p71ma8TNH+/5ZX8B+2vEtJ8qINun73cPsWB8qM0rJoOnipSrha7ki/CvLwkPdKuB/H
GnVQfOPuMkCqcAty1mAgUL7s1mqF+5gF8P7HxP+Be13F1UAnDO8DnB5MldMN1WceWAe+3lx8rVhp
g7+uXO+rD8fjd3yV0o+K3y2MV4631xHxXhjrE3KHgbTK5/rvj59f6OcAA4nNj8WqLLvjefLmj5W8
YECrAldyhEkBncLc4sP0VhahBDGolUTiFJo3J2rgy58RT1JxE9OKXFgs0dC67xXd8y9gbLu1dZsr
NEgK6ZApN0pM5eTJ3IrSiWejdjRYow6HP/bJxWsOFQNSwH1vkcNKQtlrPk48lLdYQ8qxatrVOlO9
rDOHIUWdx1VsLycxH4m22Y0Hy+Ri/vFw56haXHBHD78TsFRY5VVW4jPtxwRcpgiVGBK2tcOReXnr
ZcL7ktORfWh95zra7VKEzNh9YYfGEdTBidkiyrHGTR3NubLolAKjVgMY2QszklIjaksKH2l3l8wg
LglkGjURqZQ6RTo7ceKPBSecHvRT+gv3LyCi0Rk1I5AhhwknbH1r1sW6zfZoY9g6Q3y29BDi+X3l
/E7KMKTgm62c1ow7/rktj+NZreo4BzGaaBsGh3WMQ9o7/J6dyVcf69B/bFmKIKHKZsqtzptl0wmi
DeveMbykPHEqQPEYI+QE95lbP7wlnOuAddAhex3DC9SBEIW7MaZjcfWgoBzGX2cAVXd4HCpacGaf
ULOetWazT08XY2nNP3mqbbaauDbxst2x95CfWgF5MRkX04WD6/D7E7GwEBnZ38AS5vEjE37kTUao
cd3/Ou14vVy5uYA6Wl35VnOA+OdGQeXpON2QuJan2f5xxE7UG1wjSRDVdf6/Xnx7HvHat3YMzpLc
I5MF4gqI7eCx1ig3Dxku6h8u8teWw8Kshs50AyRhTnKTY00nyDAgAH/NdcUw9JUSFvt3nfvQF1K+
N7da7K4Ofm7weYjOabJLM1QToW70XgE0AYNqpKF1c0o7eoPTTs3AeWf8u1jHhylryD6vt4AG+DpN
heMzVQnj2Y95Vvn7uPiWnflNcUCiVRXWCK7zjU+T1tL8lNefvGkZhJdj+GC+BzLSimPwltBa9Boh
tEvHSn2LXpDfNsDN6UDbEqPwVZDm/WHu3mPSsnz+ItYwF8gckCOmh2VMAmnLduap7wmefEca3tVS
wT7J5V6ApyokI+ohUx2MBAku2wMQwocLEpyQIcucHUG+nsWKm6dXHvOxjpbZoibHQh8fGFLQWRbj
SgSbBxNScPHkKDUsol2C1k9ZLy6/0kxtYKbfuYj9yZ84yAgE+hp3yHejQ9yRmApfFpqH8bKgXKjr
GopQ19zwdjfEOEpoVBbBfERIOuvgUKOi6c2xsKIC8URWr838Rv8zq+VuBOY/r5QkU0m1bvm3IQwF
Kkyc76VuNrf+WD+1LCqLDgcobRn3YW/0NdrAG+Lu/DgfQ7TZamaBJylwTXpOrlRWwPaziFF/ODcF
slCGYLtSjRp8kfjIQjv0udN4u4TMNc1auknu8246o1K0RlLDWm3Q5ZegE+KQJQpVnpXBqvY1HUM+
eYp+sosTi6FHdKYbpkzzNw581kT9hQcaT985ezQ+QPE5Bx3Sn6Jf5A5sXyY0QlwbQMH9nVuX6FFY
B5VG/AGn6S4fntDWadlDN03uvN7k5WSBCrLmLsdysv6DI2eeo08x31BlBY1CHFz2HY9CXo7bKjsf
0Cx+May3slIhLrtoiZiJhfIA5yklu90hIzRXCNTUqc0hJm36FiR9zgA+5HAN/ZpE8+E23SCV4Rz2
l5LRGBlJRUqrJGeXUUGayUitHvIoWWRljP7cVS9iMF21ki+tO3Ned1m1TkVCS5NUEEH+XTmsFsep
6ASeiw1KKBtFLMdYB9A6FV1RuTE1rUlbMrSIHd+paTtEZwkBkVtpYfALQSxkHfw3EmU4vrVu7F16
Ww/evsAyN/0xczal7fNj+ANzepYWG0swMDIVrbsW4vlgcXZUvTwARJB27ywLw21kQIyAjLrdT+7G
HTSsmaOdcDh8G4FwzeJa9Q6e/cOtK9TCwubdaIAvDkAB79jxf7jQ9eBjnmSonYOoQjTM7mX2N7zi
9CA/AXxsmyz1TE3AJLbTRt4aC/h3X+vsabnYOFpYufMsET1Hbg88FU3CCkMkvBcmnyqmE+IK0hDy
JVtSYWpbdWk+KeCxC1GaqkT+QHZy2nGrjb0oVGH+DMeMLatdI3LxPZC9j0T09hBmsScy5gD4nYWz
9qD5SOlxxo/HWnrnI+iQot74dLysrrKuj4R//Dc6L+y/rZYxUAUIkMoPNX9c+IG8kTNJTi0sRlJ4
ag4oYol/KCQUSuBQ+jhQopamOpH11UghnH6UYbOBqqPYi/p/0rzMC2gte/cOf+3d8dkvv3AKbEhC
oh8wrnmO/YnVgNl7mwmUP7ZUeIJhlq/YBV/9ZZ3abBS2AsIGakRMQSmxgHj2AC2kN6Ib7dRfGtXx
0e5jWFxitzk726REK4KPPelNIuaH0DMuW9lRb78ihADn6cAR7s//I0mBZam4Y6IASC0cMJZrr6B3
sIDs+wKy8nlKmh0ATo/APZTTMAE58oBf0PewWLT/L2TAGf5eMzLsThMon+pFAGbC1Pe3TK06mNTs
99Sd35i/KcPF95WbU976F9i0X9DaV4W/l/0c1xwgb8DgXXSYtCcccUZPNzm0vjhjRXKWED7SDa2g
i/WSpMrw1Q0LxxM85xrMe3RzlrZOeYX22CspAiKHZVUGu1lq1/EtMaTbVM+OzzUxpjRjJS0qijG2
TXLZmSioPMzaqPybX7UFAbvjVszbeIsG84HjUnj/UHfOzzyhIpvLDfcBa8o6XDfnzgMJC9gYfy0i
Y6k0F+BiAtk/FYw/hTJcRK9khjpnrW12D56n8zuAnTz3Z5VTD7X9rWhnI/Bf3I+j2tsIEpTpX0fh
yCFLME6OSFXf8hd/pTgCwcJXShMqe8IEobwoMbkncyjmahLaWEq2C/Tf7IPpgsZj60H5qNAf766g
K0GelwOuWA7RCWWtVoGkVstloUxNgeuntfEbAPKMT9WD/xjaCC+Mc9wClDvd7qHrH+ZlWKBS1Yq8
GVcDYHiUhhycWXgqpNdbiUCcNydiDOcEHGr1FE73dk0kwEYe/zELo891AMw4RzpYabDX4wMoKwiC
oJP0lB7XZHtEfu49RrrNsubXU/gAv+89NBXHc68YJlGAnRWFLzE2iWuxwqSxg9KebF8ccJQRN8km
H02ipS3P3zVzDu7CicHs2EkyqYy9zVDz0vUs6VDWMzDTg8z8twd1O2FUnBDCHClcN7tfR2wgYH+/
+cjWeDKRF8oEygvwIfY22WyJFMcNU8++LHTTEodk7e2mqVaeokFYbOuOxK1L64+4BZrNpZTE2bEO
SuYmQfx69IvlWMLc1MZ1VG13XM0Vv1voK80W2Q2KCdOYeSWv51UiJbvWKu0vqxpkLU0YmvugXGsm
0m6hew+tBC9cbQ9VQcxvDox3xVgL1l2ZH+apcnliZIHSfvmqMVz2qG1fXTqy7WPRmc+e6aZgKsKA
eSh13E2ZEv9pVRWCiaUbrXxQk+tE2pCwTyx9nAkVkqsbYtC5OSSw6zid0W//qjuJo04Fg08wnCjK
oLct0FPLJBQgC5/Ii5W1dCSmdoUnNPT83MEmz9+E3HxANao8jrX1OdCkfQSkhNDVUWroWNisEnyi
/YWVe1EFYiCY4rsaS7CowziWyyBjlpR4ueTYu54PvvAczLBFqRAcnMP9GVevjcWZMglJZLIsq0Ie
fiBmXzbxBivg3FFD0jsRk6d/6p7E5u29kRjZ9XziVgUrW05TOQxJ+wCNqlbIX1m9ZHEyAGno5lOC
97zTGflhZYCUseOtdcVS1/1RLtKk1+coUGIbDT3Z8JvYYnNTUJA8yHbi1z9XR0XD+MNc6CEiOapR
Ln2dJi2jDny6XsOUQalJROymtDhdQTcAsCCcB1rvPlT8tpLLFdpwzbTKC4K2Y1a1vZKHi+b+/7Ty
NfdcZwbK52LjmuYLbnLZRMjiqxxIGWyJ7Zq/5cvn4ml2PXBN9TgeInoUhmOeHEQWVoLaMewCsLLN
WGzmOmt9LjZTlck2oOOx8M+PKW9dflVrNRBPi9JKaGsn6TGX8Bh5UqvVFOIZQJfmoq+p1zb/8SuH
fYw1tQNd9BZJq7CJReofRS247kMrn2rOr1JH48eJ0ROuwqgiUEwUNxgBGB/3BS1oyGmU3UP4SfVZ
1STQTxtWoSB5VeWjqIqEKyFE2eexDNwWInhXXpA5AqzWRMvPhMjgSv44neyBhBsZnH7fbEWAAyCk
S86b58sIv3ChtR8b1Yq3CN9X5W2mYAixQHY6ysBNYdgF0at3JDmsA4h8aCcJlirEfVIYg2w2bX2j
Jy9LKF95YU13jTuRDd9vtlVVWzawGFcY5aFowJNsJYcqKkUfj50YL+CdDNPGXugLufX/EJFmi3gc
Ghzc8+1HXiKBF7J6t6WhO28T//OAVVSkMbU5hmHrsAwXjN7AfPTkuthceHibLXWW2j9uwCW5rnbi
7+QVpkgDP21ctCATud7LRyRdY4Rm+35wNDArcpA6X9yAHORHAdATfOtY40MNQZn7831VTwW7FcVo
hGUG9dDjgZou25xboMqXegupRu8Qm3KYUObCc0Oh1PSP1N2ONAZpB3TtExsuTa68e3eGVdhkp+pi
+OYDQdxKsgLnq2wqv9ZODSxzaGb//EBx7Xr6KN+vAIYcKCwHJBmwY3UU8ZFcuXp98FWlsriRtKLV
AEuPc1f+zO+bDS2yeyhyAV55uKCaLbSDal0JElDw2twylX1C81LBmym7U1wYTdNucMeqin5A4zvm
1N/Z+p+i34AWcY5T6Jz4Lp2PD7tudKyh82lB9PKAt3uXKmfO+BiNmOoWH4Gw1hgkbxwdcKs+mdSu
NxRq67UWvfAf/pj3a74pN1i8a0gDQCIyLt/wrHugzrWu4LXSFJ+s53R8DKgHzlVyR+QSHLN76mM/
dKg/E/mcOLKEeAnjV1xX8iHKN0oc0M9RqYn3IRAgsCFqaMnY/ssAHCb+muUgGSF6MXVxuKnJPIwR
YFd1Z6QySGjmFfG7gZTp4/t+7Io2rilRDo1PkT2PTB9snjPSB3JaTAQHeLr6zOxyL+2ImKOqAfzr
cNEs/eYRqEa1n5O90fUJuqgTdUKPzx93ZTy/J2X7N11zmbqId9thmrxOc1L/zaX1p7N/cUbE9i0C
jM8enwO5WJOXscsaqBEflkhJt/2ePNouD0poCb8UT7w9JD3+HfwhcPJHhjLcQzYNT9VWr0ThqBPa
3Y8pMijZmDDZKsgqoO683fgA+51OQFXuPgb8vVGJIfs5YOk43JeIVL6k60ZtVdmm8R3lFVmkH4SG
vJqsTrPPVA11rn9h3CTNhtOKIvUTMlgfrEHirIzb55GjstqSVPVnWTfeqZ66uQh/rJJ0F/9vnHvf
CeNZhIkEpR/+WfifoWKYP053C5tBVgGMwiSKgOZ+AYL46tRtLwVuq0HevLF2QowZAaTiG/jt1Sy/
z5c7/7Zj4x+fxK1NeV9eh74DV0LsH9ZndL9dAObG8mTX/RxTVAsCTRrq/5YD/L8ECj6DqHlB2RUk
5R8auUZYJM48PiAOjvFZXezG/kMv3CizFOt+MwLwQ5Mlg8tkuV8Jm5fQaYE8IPmx2mFw5jNWxATL
fuyKDiOBP/He01Tu/hxTqgRBgOPOX+rLGeUFLu+SdhYU7UQ8ivAkEgLTB2NCnyTmJ7cTnIsgrHMS
fi63nB8K6mvFZZmdEbvM17mVSPPwOl3BJ5KYdAt/n1uxwS2+MH0Jw9c+RZ6wAXyVsaLIMNF8RLvn
ubhfhepqwiifgkowoE4BB5CDv0nXJS7LYjsaT2pczrEximYRGDGZqaT7TdSkQrWvhIVrIawMy8Fk
5GRd9T8SAl8Qpd6XmHXlVxyPDC36l89kZ/y2qSWSC2FoFMq2ZH7b+VrnJiNGfHpbcFfG5KPu7F7X
UBtIWpXg41HtG60Aza56Uyz4aJK6ijiW18gt/zzLP35y4PJrJ7Y4//D7g4CYK8EWfksROK/eesB5
KqtsdSAVAkYRYE1iBnPxemE/eOnuKuUu2HPfKVXyK2LXimsRXp7yJQxfCzRl7WMBrxEWraUCHMrL
l82/c0qV9ZqiT23Q++HsjXazLaGVZTBCI9CnAjOFo/y97ZS5hVRG5xPL0nVorykSJnl9lb5HT1AJ
41ujb7n6TELgqYW27Qgvovi6xcGXRSf5OMXcCjckwHn8l14fM+liA5WvfsUk1XKGUOwtMJpA9m9O
EB1VpPZFVDqip276zcMjj1lVz7VLct67rQhT8fIJlG/UEh7+Bc5qzwacEGX+kVdOSDeqFTdEv6Ng
4YLWaKBWx8ha4ibfD97npDSXvDE0m0zcAHXWhUqyQKlNZIE6xuxL9TmaojB31AX8l6szP53M6EJk
Uxk3fgS5UiC5Tt2UZOHy90Ilhbo+9YUceXsghSVwOpxexEQY7XZG1bMano8b1E/jJigF8yrD2C74
OMQORBOd20Nb63LimBmC5mLEpPXPj97mLLilRmi2/Ot4hEemj17RKxdbVoykAMR9faxCGt+Q1033
ga8KmCpYbiJIH3trZF7Jy4am4zgdCw1yuDB1UMaSZrIRRrzGVeU2MLTrrc3dbgLbk042mqogqmys
U+KkyxCdUGH/boGfF/7M/hyEgYeJxVzgkzk8vCvd5oBrbRtyU3BnANA6oUfq7qrjWHVxnvxL9Liv
WzO/qZySv4pPWhkFsEaCuO60/Is9CMJE8LyMEk1JuMnGvMPWFErxtZLR4/V61LV8pD06BD2EedlJ
omubDPD2Wm8S85TsMpltECR9llZASeXzy2yperYkamRaalKO45c/7/yC559EyA4quKuRsk7zV4nW
qc1Q6QeM0N5rESLZGFfBGL11yksXVHDVtuVFmOwbaLd68Ti2pgwoeUZe91HOoFiFTvmyrSJTH6AZ
CW4u44yfTGZ3QRolql/7FdYxIsILu8Nnu7ZXe53eVGtx8wY1UWuQpCewpnYeWuWVuaUrBDM1FUnT
obCUKJaPpD8TkRRB+fIHZpwKDDlfyYZ8zOvhpMo8JnVDIUl4+elcOJFLUn8+rt3CYX7R279X8230
cMgCLTe4cSefWbhVV9myp5sL9poX7cKxCeGpQIc8cdl+/LCGES9VtWVgq5ANmbc8yqwHnovpmjp5
hIah52SnaPyzCXHxjqIDJ3vlo6Qte7zM5OoOdFS14Bqd9c8t/O1aLuQfzyCiDxZKeFFbFMAJ30Zr
gTuxdsNl1Vwur6RoEUrTs7zT9N5fkHneFWPn2Lictg07TgAuGE34DAiZ3bIKvgMsr7J2WnkznaFb
2p6wl3dZzrqNbUVCIEAXpd5H7vafZQxoPJqSbwzXNRP0dh+uBXb/vDcVWmMcZOs69ISMw7JloRZ9
JfDq72Ser4OgfP3dJQlo3E32FSwJYwcQLLJ6tPPnPgDSZcOlVC5RS0dnLMi1RYDoJTGmj5We2RBc
k4wA9bKKWo4Lrv9Bj5Bh4E5+JrYB+6pSQ/i87Ry4bHjyNNe3ZQCBZDtZ5zqJCqXn9TKMC+EixV3a
eaFvTJaTrGXp1YjufLAWWYKA8AGBtlJdL/VYRiiFFNYOB/jRqqkocltr40SvgbJoQkipKM5SBmUa
oCXb8oYvnDaSxbh+m8fKIGZYhqk6Kctz4gWI2FfsWBhFml52Gw5j8D0mfYWIyRxOmtPrtB6mm8ue
lQ3nhgPIx2RWzRg2QFPsRpYEJRNr1bz81/tyvJeQxzkRmgRc+QQjxB9y6AeB3XEoH0caPfNnfwRf
zoT6zKugdatfsE42PFf77OzNzCnyiBKcuWTRd1rrY5pfcKjqyBAk/uOq4m465CIgRZxATpwS2zYu
oMao7ADforuRxF8nBVn1KGtaiCesemRuU/onpx4ZmjMkA9aUZwuQtAtzGiIFfazsPFo16Aq5BwQx
4L5roM9gugoUPxdw3LP+SppXDL7qcVVgn7O/movGa+qtiV9iGVHhGk1jVLO8q/11DSRsRfOAjj7S
7LQY87O9E5HB8Rep5WKrzuG1odxq8d5evdB1iZfgVMGmSWoaYkQ5nF3qPmiFqaVvMWqZ2S8taEUl
cS4sfmSKmqoo0qKa3e8OZxlwesDlx8RQMwHLXJWMrUqSlXEm3xUAjaOiyxoshxJiKiNz72abjzQt
2T2BreCMe0gKK5q34YFRozftvJRQIWlZbZOTWo07Ddv5vqX/2ZMsNngSUlc0lCqqIBUQma3F8rD9
obApJsufggd/wEEjwhqDJw9CAxqWJc/+z3qyWJ1jo8eQ29Zk/7IPJzc/IqE49cwsk+viqB73nJLs
1ss1/G7RHl+/F/Ka/fUrycr5EGD1kbdaFeYgriiD//7/MXbilBT469y5lHCCtqjqxxCBF5K2IcYT
xF/JRa7/Vmhgx5rhwpQy4TKZ/RRWRXlZ7T0KwWFwutX6YOOFXxNV/UcD7n1aEErxt7swtVvI7SEe
XOXBwmdtBVT62DDUdaLr1pjDmTTbnsbPerI1Qv7v4s2D7jtch0d/sRV6Nj7omCFpppFuGWJs724i
YR1x6O2tYpmEQKuEcogyikNEnYmRJ7K0yf5o8TAznxETvF1DbTMzWjHPLAR0MGG/kmr7TsNgK1Xk
UJMNocY1kF871smJSF4ZMByCHIImoLjXOK1LSCU2BWuEkIIPVZbQ7Fgi+R+hE+br41SShxihvSTy
Ph4TlTATNRX26EDYxBF+3SmJolTD6+Wj5clU2KORPWRHNA2laEk4t4Ny5+ZhfeARqRg+0seAMJCC
LKfsNfOyrWuHHTfqA9EKAfNNe4mECU+FoFqNnA5CMmdtW012n5gyttuavzLs7zothD+dS0iWDtZt
B4TUVCAVhPHvzMTI7m+9Z8QD4RWHgw5nhQyVxbtRt5thl9KAklrsPPiq1cGLwiYVCVr3mTpyDSb8
BNCRjMX7pTHW45bOG+OzOpsuFCFYISSnEduKzkH2f6ZxBIV+fBXkUkKJf2vrmTBu5aS/xXNorklc
cq0tkO3bbgjSY69BV/Dpx8MqyDFbdBl6yxLiFALOn+1GrTCvG0rZXcR6q9iz1ZRS/irDQDbcAj5S
NU5wyKvrqhmFs680hVpXujXKGLaYNuv3+iTuN/mAqziNhLPF1gqpsEv9imojLzAwwAs8gKRIkQso
nSc78t4n7ZsIu687ZhPdh9vPqpjxW2uwuWvieNxMexmxGOv3fKMXxTk6eqlZuk6UNHsKki0+9Mi/
VRYBe7MZfBONhPj66va2f70SYZ2cOH+ORsnpaHOi2Er0kTc5T0z1LaRXuJAMda3RBiNTDpsAE+Rt
3ZSeWeSOSa9LZkmC1FxlZUAXU5werAleSJNBjPlRyV9Ctvs94rv5eVM0PZDOZ5yeFLA41vRNmvLV
xAuXvHlcIxdi/Fi0X53Bcxr8QTWuVsobJxKXA3+57cqtX4+Hx/lt8SDVwGtyHRGrWCkIFzUfkHN/
ddhYcC4+yM9pOJnlr6/rBSvZdZ1DB50LpeHEwPm7El9A8foOArnEK3fuBnE76WNndhwpeeEY0wti
Xm28LVy3lLfBVszaIWAB1jcoMwt5fcYcsGSqPFL4LPBB/UB1wlipnfnsBJ7WvMS9kpaU8q2gOrLr
HjqB9pNoZXTDHt9RkwKdFjbD16yQGqKI6bcLssW9Xlv/hGXLUhX75OIXOApuQa8gPlbdZRYD21Vw
kSm5jOca6ARmEoBXBKuebQ3J3bnvVfJRjb0CPqQDtQLmQrrYD/slKZMvh6S+AS2uf3SjSkEmgDiA
cvYcW6/65avBy3bHNId7anKZ03nPUbuMegzAvX2GHg2meIocpjRjBkMpfGisc5iiqHa4vPxbs7vc
I69g0nc72zfqmzLHFAlgT2SRhl0icDxEsVtdEUDcBS41ekGL8UNQQ/nbvhj+Ooi87LYgQxLVmWV8
YerqZdWfe3F0L3DcRl3xF9elzguUcgaNxIkxS7S+C+Qdu0yTyKDlQ6ujMoS0D6z8zqgKiYaw6w4u
qVfi3xnlS2OtJEPSJfbNCCjTv6YkvmkdR1iIWEzJjZnMzO108A8vctgjq0tX2H3lr1pxCqMv7DjX
Ilbo+Z3kGCfUkPFI0BNSv+mk9iUO9aSb76uBKOf9dFCyUjpnyBtmdAVZ9U3/2zqRQ6kN/NS6azLb
u4ohG+rBt+DpI32HbPXoRoQLEQWP+YxiecmiGzdq6qVmdL2dexCZQ6p6NiUR9bRlfT1ceB9vmfnk
CfwEU/8mYehEsWMCI9HEN7uo0GP3rM+1k3+jO6qczwwNwnDk53FghOe3ghfCIDwrPFm22YbqSHfs
1OjEWh+zdxdXn0DfRYdck8QiDI1Gl01WkUBjTOtGpBCAs/pUBzcio8V4f//PYYCeVeZkcRVAuoVP
wSX8W1H7weq8FsmsPU0ZQCygu4CHLdUzEndH1DKO3BDTY7jpESwqP4jODe+xlWTWh3x0F4UbOjsn
SLKftlDjlheGX3oIMEH4lN4ei+GPtqph2znfrb/7hhRydKCjzuGvzfOr47RU8+WcobOcu/U3LhEH
9mTef+yNCy8GXr14KSCFJJJ5jAt0PDr604H4XvEgku3mRe3z02DUU/rlcgcdL5umd8yxHduk7i6+
ENcvHzliOh/7VhVSpjdXiRrBNaz1haKaYJhTybzarImgsBy1flIT9UQ2NzRLNoUOEUJVwz8Z3HW2
gpCEXQDN0jfRXuUGz6BAd9UdYmvui0Rl4EZu5ck16bv34DghAL7Fwu6gRbKOAm2aEOIqYFEXLo+d
xXWFEZEBHBZlb8O9QdAtH3WcpPGritiirKrCNmj43PFWzszWT3BLjaCnqBd636xco0xugP6Y1yOU
y6V7TPlFes57zCd5PDw2wijsV8heUNFDZDNJWe9DiKfNj+2tmoP+SCW20ULRUWaC9Qd6GnH/PWkQ
Ye5FdPy01wuisIA9tF67R5vhrDZ0tMq4X8bskgjMQvm3AbWmmTKkrjhyddryeu142pY6T6rab16h
m40NcyAvRuK/gSfifn38psxImGrM2teQIIhbaJeRu/n5eazuTGqYeYWkYKM2MKOxQfMI4KixCMOj
ThTFEgDR5uJKPazPzltgRquQ/dkxFsmTQbxpey/1vISC45G3wKntYduDTQRLYHg70IGkbaQz3hXD
DUxhz9fVga5qP5iqPqO646dPapcQui1PjwsGwDxdXS5b3HB6tk0Sv8nVxhQOQGkuzLZwD+oGF77G
HjseyBw3m0ePxqs9x8SlO0xgmFDpnjIfkLceuPkoEUIdRcCJXw1y3g78fYHuZVOFoyfK4ex7KpK+
AIRxVuEWn8NZx+Bx0BDTcKj5Y/V2UdWH/ChJzZ43yqA9dNUit5GM/0hQgI+i0YzuIl5RculG1GBO
eGzTx0y/SrWeORbOvTkj0wOLU1AjigwIRoQbL3a66SOdjBkkf7kLHDVjX7CmTYFMrkx6upSpXXsO
I+os0CUL6Xhv14AzV2FFP9jWTlM9JfIRfLCgFVookfCHXOslZmDIsRItnx+Hff7kNOtSZCDh76eA
q6KckH1B1VzoyNzqeLNon3BXSRURgt8IbzTSZ/97NmU5R0Usa+9WcwETfA10WSEj8SGANbQuBklp
m8mG8VrYS+TfPM33/GaH+tK9uLrqpx49iUmQFVBUrJ9yf6zDp3zMQAIE2tiQKg820KXoyuV/IQ/T
WEl/Jc4RDBBQosjV14hg6L42SEDmFd8cgAc7bbJB6NXlYMjllT1Rt8L6HaW94wkmY7XeNYtci/sx
c3fUKBLhpABX5Eu4ZGlAAY8rki4mcjrghho4irbohBI5PpebDXNWyuywZ4aA3Tlp5QhsqNCi0IET
zy7fkbwKwms1bsB42FNOxyBbj6a5nYOlfk/knsT177duR5rfUp7clEiVrSzFZN/8Okp/axGZy/Vy
pGA+ocMBl9J64aKN+rLlhUiyyvuNH9ThMliW8lb84YjkinBwsVWEzFfHmTfK1ij10o7hdNK8cfpa
zkJI1m6OOmyS+EDxLZH1pSbcBOq9SW4ZqoYpU0bWFEEI9HX6olu7sJgixgORvHG5cU3EjQ4mtweu
Ux7bGt9hNVdlL1Yd8E3IutYGDrEoXN3iHtQURVMFHT2EzZ+lv5+hlxHwz7eZztDxB14Zbp0veVni
Ek71990OaAUk6u5fHBM8XGVQP/4wOvA6V5VhyaxC7AjifVGJ3W8NisXFXq61gWuGnTRpHEzU8HoT
Kg9ISsLSMGlz3WKw68mW6BW+49hdlIrpZ5zuMbofO8Ez/GR1hkMotV4AEwg+OtPishtN5W+49H6m
7oimJqF5L+HtWE47MccieaX2rRPGJCQ8dE1mRiuJbchDhNJ8YDKMQgJa9vTvewmSYIYR2tJ9cS5s
eZGcaFZCypePhS8vTLfotsIxmoLFlOxbe9V1KK8Z87hJEXC8FYQTSVM6PWZu/d6xQITx2MYe4v3i
9MrQ4e4w0Qhbkve6gyQugN7zwPOnJ0CnpBGOTsg23YCs5O07U+wshBNSSOp1ulGLL3QiQpCgg6uv
+iis2r2/9bkBr2o3NOz6a8S20BU7XEGxTJP7Q7jK5V8mDdNeXQVbdrIDmqBGzECF3grhBT+Y280T
+oOoUnt37Ncvni3eXA0zPgogAW9b54CpGtCWEY+D4urMI9hM0Rifz5zWGrRS4hnLdYGf4ffWHFw7
3zY2q2+I9X5yHBYXPzpLMiO+JA2/r4RSGFZFCgl6NC6h5eKjmerON0+QWQy3iSPDHy1lDRmC2BQk
6Yr+r4R8nTZUXn9JHz/lBc7/FCE76MgBYLtjOe7UqUj4GSdrqg6Wy8UlYRVWh3zK8eqvE4W7kwv0
A+QQMX9l5XIuBPbSLdZ//pN9h/7JhWQEbpCKsRvb2zTKbj+yYwOhs299sRE4OIMVUGDoHapHOcxW
5h6R5gtLi/KUcis/6bQJFPyFskdXl8f6qe3CE4j+pOd5Ex4gOwAvL4XvP81AGZZWLiZNIsjYLnNM
g57n0CyssIU0QRcZ2KERkTrPsY2Z+Nivjjq542O1MOa5F1jX2F2BJBiAjwGrNADn8f2KwQaMYCsm
FLFl5KdTcTXN59+1UBIia5PKaxUuGYdmcoaRdenhg2K+sddeD8qArNY6Oub4ME61MoWg5975AUy5
oUW+9HcQSPTHokDvzN6/CmRroA1h+sImDUxPFDrOIuG+t3F0Ej0qNEH+HdVaEXbArHcVDGGpIpWd
K0mbcvw24SaZg9cLIDF9JM+SWOhJ2tjY7EjjPuyDQPvp0m1I/bD0Rw4SpNbeAMRzlgXJwJaZ2gup
gBRXtyYRq28MW/Lsd2zfYY6EbDYMum8r4S2+XavMskCj35plmFze054lKAf4rk3ovwxzdDpTCjwU
LmS+p9iFvIV8RcNgAoIAX9NW9Sec4r8YG8460QTJuabYLmaMiP80KDYPucuDSud5sen0o3moEhtO
+j8b0FBye9Nw/DhGKLT7JKTX79VEg0ZYFl91pf6YOXbcCdmNBYHfKm0N1jrqLRxKKscfiy0IYw3d
HsnKhM0Qh2wyhsdGGrdqCpXSrgg1IUZQizhx5HqXhpbmoy1ENtneMCKc7L7zxh1ulbdfJyTMm/T7
aFqs8HgAWTr26SG4mW0stYQOfyQAxiihUN2D+HzwsKJMxPWblJmvPKthEruLjifMntzIr7eMWKN1
ZpJDSqjXpeTp19ig6zchVXZ81aixGnPX3KuOItfcStx/3QMe6TihfCv1ZR1FlYLv4P2Rf7su2k7k
/LAZEJmH7j+2y0Pm4quf/F8u/XR14ZHgR6seouAqcUnjwDQGgSuOdkuIvZdrZ04SkreVIwZ6PDwb
b7945R835xKp6PZZc3SGs6yRWZsYH1k9Yd6zwfI1bwezGPcUL2qHF9cWHA5OIjsjsOv0jlV6i9+p
eCL/pcI1e7sgVolYP/+QnPPjVsp6TCJ3BLhge3H39WYBeCYOShpAQxvtvQAgiIEpuDyUMIrgFv6n
7y1HCV+gYwxmva1qLwLIZZxNqrJ61+t4jDVyl4jAIZYGIqMmj5d7M7meqI43rmIRs0qzApAslW5p
sFdWekp2E0ACSsFu8XdsC4YikbOUFHraNzusbWQdtN6VzWvUCqsCVLHJ860RoSgQy7WEcOQf4A79
BdUIXedYWuiQRYKXWDaS0vt4zktKMe0foydmSvo4b86F/cv6LDZvGKfKxhgdgLdicrIdFioTZy51
2ksa68EWD5pJc1HlRAiJ2QbWeiv6Ck1SiwUeAxcRu8ZG+LsehDBAdsKWkLzr1hcO9Qj6G/+rMeva
UybjPuVtrel0eHr0R6IqoVtaWPnZP3cN8GWxuRE8OCxkMUjDnQmkD2K25aeT8IKSjtmw7/ZLV9mz
NJarmbQpFy8NFHul8KBkfFKQRKnpd7esFcjmfxQuf8vI6bZaq9mriI0Wxgtdfr7Yw8PFKiBPo8JB
DkkJX94EcuBsjlggfggHUNDfdXxInnXsoJjBLkom810Dqy78KdX+bYrfmfY2Yw893uvM+SooYLAm
oVZJ/pYJEdpg+RiXz2jNHEHXlNDalaW/COfjLNFXxR4VaRqCF4uvMM8sDSPgEiop1ydrNK+8SUrp
hrpRL8aXX2ghFRkNNLgxhYERX8urcL1WlKtOw/AjtofY0rGkDLcwrFFmXBilajAC2vJXmj2B/FES
l07JpGpmWJovbAgzvMP/iM5u/oMRkfb1gTIgXRp0KgmiOizvopjJsDcKcWBPCVZLiH2ppitFnGhs
D2GYXmYLwcj/CpRO0a4DR+l/Dl1rwAu+w+3yTRLGB0Ef/tj8LD0sdFZ7A/Zxwm18zbLxjkuGbxne
80w6nORvH/U0VV/k2/bwHgSY9DhK2l6wF9xgqptTTCxtAdPRzjD8oAInGn2WfQrT/Nha9eTCCrDf
R7sIFRNb42ZvjBIH6inhpPlqng0XRHl9+dQbL8KvcxjXpySeJfN4j0h2dbJ5g1HYLJz4kzf1LQ/j
qNFwzUqbk2sJAJN2QAZQeNhx9VSgwldeqSqN0cyGToYd5LdanRh2Ng/Qc+dQO8LNcgosFAGQZvOD
ws18N2T4L2dBe+yGmevkFy0l+BNqJc7CMOCtfssQ8JrJGqC2qNZn3nycKc1GMzVjHmi7hzmDk/zC
aSUeeggEI5OZF4xgByhNgiAs1msebm+axvvB/AWvtzqIDnHdF81ANQTpxsR3eY8rxiN66WuKn2Jj
gc/SbC6nnLQmNjT3X1PC3ttl7vBljaQZAzmM7jV/saVnWG5s78pMLg75k2djfDs/7XkUHskarKku
rplILcx3piOHfcZGMaCzviZ5NgXKSkyTwleJAciCqoMFDti8/LoVAhSRZGJG2Dm26XqXfcGC+Cor
aPcPx2MqF+tR3oG5hIaXDsyUaKimcKWDXZabUJEAv/sylc5YTBmChNHZ0FmK50o4A0v59SRjS0jI
07srzRCtcoNgWbmitwKOi4iDcHme8uc4s7SDfXukEo9zztsgTb2Dv8pWjipsGekxOOZgxDmC2DXd
AKOHi4URCPl4brsAWCsxZZ8MQukMUMStJ+fuq2u/eWwAL3/k74PFPh1o661Cq7KE7oFn49eNOz/G
s12eZkq5fmLTOl5xwCRmO+qf3VS3KwScKnzMBGzMeLdH9bYZldJPeVJwteH/p/+t9X2rpFHlYNF0
lnfv4XqK26xi1WiqFPUClDy76iubmg0k1A2A+Ypr1VTiaNJQtwjDyIj8Z0tEtu1JtfwZG8m8pzD1
tNBmuG0azFzAq3cOt6B5GdSSmu8UxxfHp8ymV9monmD5kiMngQd+BIqPac54K8hLVJQ+SbRA3OwA
AnBhOzxMPdvSHwfks6T6w+AL86NpGMwszmWCcte4fkqF8N6jWAORS1m2FB7kNcgbm6rb1rlRrkuw
5jHpHjxz5vCSgTLo8ITOIRs3CsfAQeVvb3BEgiIAPYTwusE1W4Xtfk1ZkFSv1SI2sjz/V4+52dra
I4tpAm19A6sfYDyNwVswGxFCax3bNdh2T6e3ttRqfgG8Ki+dv1OhTO15AOovOVCYtlND0JOS4kxo
z+h3TZ41eolStXP5tBkFP5mhsGUrNTyZNUNPCkvw5az1y0bZ39qScgpwnohEE+KbO2T9U1dDBoiH
OG12Nm+AojoNAkPXOiTtTzwkmzzwHAFhWqwKoB3wXPznIKPBzH8SAwdQXyAPg0IeSATHUIo+LWQH
6Q4ie96LyPXK1dHjqaHlpIW11bxeQHqOlrHA8IFb1cTBSuN1+aEexEG2wppIqWsomKoGQuo/XBEb
t+XJ4CjNbagjULZ47HeOjycQh8YhwU//f2OTnDoFWtiMzpIRvG3IK9nktBpvcl1BN6maPDIrwMOi
E09PWaUJwPU05duPOuCL28O51etaxmrajaWK2G7j91qFHHAPsrhzRujXa9vXYkLlwhqfXBKlBIkX
Kg1GJIowwsLqu1yBDn98eOZeltJXdCGByUa922MsaEMLjqkM3GjBUn0TlCopySSo1Jr+xW9VJXxW
6GUWnyJJ1ZlGhq3HiaWKuX/ZIVACCvT+IQg/AOAWa6L8bN4TPDxaK+UYpolucnK30jIwtMjUxWcR
mOcakdtGpQUA7N9SZ+q2Ts4mzqm7bx7iUSr+k+Qoaurd8zWhuM2f/j8Ni8Zgj24sSOO8mSkDknk8
L8EvAFFjxF+7yb4So8yR+iUT9hgp87x8B5xxZKAra/ApIHzxU1lSrEb35Mat5UaN/E9lkEb3P7Z7
Jm6zGBkslcoROq/6pvjfiRUS3Q5Au062c5q376D55LZiKS/Ct5WXEuWy8HlhsbDNo7Hf3tyq5+Ex
/pJpb+VK2qIXhlRjvYOFiOPBmy1+Xd1LAwvS9csf1LAWmxH30g0fmAw7KK90AM6nZ/MRw9UgJio8
qBIXLXvY3LSrfeLdoaaBHIhldcFR4RLQQ9OnOhjnKJGzW9NdNyZNv+oWa4Zl2OV5889btNRXvPFk
+AahWKstVzKqjv88NU1RBNMofyJdSttP4/4qGvEKkmTT201shkDr3n17Zg51jJ+iniTtbW72p7Df
XRY/HM9CJJqryDh5Zca3lXmcnrNMme5B2hi4WJ+5SvqpTBVdvhm4xUXaB//RVVvlVh9HPVpkTI7h
omWdlMpo1Q71FZS4lhH7epW4FDTkILux2SPi+WmwQggvWyow+X9urUBC36spf+I4gdbsSZbrV7ax
jmSuNvf63dxx/gHUws6W5FmjxxfhIeUAAzrivp/LWq/WxFnJLkplattlebyel5WvU0Xa5kQqFdjw
T/mp0O1DcmcFHIolA4HY5kebwsGKd+Mnq74lrn2SRekdPFYYvvMkDtxjyLIJDpRFVZ1xwwjXgUy0
RFRgHG3nswlHlSW3F6lsNk0LXhuwSDlc6VIqLk4iFbAK9S/Q3SOwqjOjOSPzFkzepeER5YYJeFjO
eYkfEa7mAtugDRgo6OWKKGodd7nRnBB/zK6/Vw4CrgdYGwG/QOs2R2OY/f6OhszSPE2Ne+YHe7wd
KpBwjQLwSxr9XHT78QVnxKhfpqBbRHoMqwiOlCm2Iq9VVjirOTXwvCwJvq7eBRAP2JEbGD/JJMa/
3OTUgOJOHtPRdFQ1ZMLH2NcV8FMzMRKR31Tlful51oaxYu7HmQ0V0PcXdvfOf02oqAH6l6HMyIyJ
IvtYY/E9Iqzf+WNJVACygI92IazRRI51gW9fwU3lsloS0wmUWaa+6ILXJk7TIZdpa+sTe5oMX/FM
aPz+jRknoXy7NhtRivOwf1BdnxwTspRymqlv96Kfn+05rFIxLgQYqNoKvazr8c0Sm5ICJwtCtr1Y
8UqA5nKgbkvuV966AmJbAIptSJ2AIH+b9tFRbcU8OAae2z9OU4eCmK20o12AXMAZXJhMNMEwMsga
DknC0GKGj+QSSYTtIzhjK9FiaV828ZwmhBlr1r7FITYXCy+9LgF51hl/Qy4e5IBuPBjse5I0r9zO
P2CgUBb9akzoiS+dAmJPHrAl7cwt0d+QDScMGwek7J2kscZyPvOKSKYZtOaELEEJnBSEF06DaGh0
PQlxbPnqTSbPObcWF5aPnKXm7jY48qcJxQKk2eAC0r3PaQAoBUHdkIbJFh+MFmkVrS/oONSqTKyD
Mo8fPz+F2ZtHdgkLMr9XzyEwR6SZqgXl4s8ueilIi1FHcY74rnnbDsorC99CmNajQbICUbRwvLua
z3gsBzWSQzyxPvW2EFymHNZ1GfJTmhIiKp2HCNoY1tcmtEQLyCxkqiYWSUllnyuDuZ4jxSw9r/LX
lrW2flWOizrV862NZWaBVkPTY2L3q0sY/2kPESynfTYEytQ1kqZdPp8JIMQ17zxMfuJa8nUvzhkm
Ya/TGipRlLEdQAPjew/ZCpHXlseoOX8Hnx0b54boFxkFSfbclVWGqw3w0qHjXuFQMTt8mqErQlAJ
s6nK8Mt0+g9NbLerer3yVPn9zgeg9xpDSxzTf/eTYBL/naVWChumqoBieth9Hyjjg5EJZtfZgVvh
ri9W+zDfVxK/dGT2qCdgiZz1qCRa5ceREDmKT4GRUiBTTyGFGY78yZmvnVds3uY13GUyZcdcu3PY
vWfmeCAF89TPHOYIYmnZGTcjILhFasdvvJQf0AFCf+PGSC4ctjXhYvQSLC6rTW28EN8L7WG6vhPp
yXeawJag8yVtb/hIGGFc4rGRLZlG/H29Aa6kGIMjlaqLG2PoZ5yuRx9T3RWDTMN9/bjg7PUax8gf
y0hLfGgVWGaaJxO+1wJlSuj99hy+3mfHHg7ZkAlW+HI7aCUnVRfysFHlUmkO6OA590JDdz6I3HyT
nhaF9WotmntrUHnDvuWmfJXgYwiJaKtg0ntchyc4sYWJlVdfHc2h0nK1jPtNws8RmOJlXZzYUleq
2eiiKkakgy1FrWA6QrrMYufsys/3OW6dCWeoTmNx0t8FHzzICMrDR9bUdatyy9ArhwD32kclbv1V
Q75ldT1qMEF7tRB7h0G+7D/9xqB+Xl8QvDhhjS0rVbSCAFJFDZaW1SdTCZ6aiZEZlXw3D7UYD1kM
n9WM5UpT+PiAQqMADR9jwMCMlNl1RLY85xtUsETjWK3OvtWteLtFEDdiVbXZaVRxF+ohJl5Mu59J
5mpTiBexjvxVcC/U4Fy2+99ky+BQpFtWYIzAuYXqdgq+cimaG14KWtHF62R+l44L+4JdINfAVQ/Z
S21F1j6xHqUya8jxITHMskUihANr5NggWJaEc+6dFiiWa0aEpywHKbzkGQG9PdVHtBocgDl7xY12
+TxHVtyL5qFTs/Pef8rNU/pwwehiQiQ5dnE5WnE6J7mXaT7P8+cwPsz04nDOSj5SwI9KTUl2U24w
+8r26Jj+xOuUz6YbhRTp934FfN+N01H3eS7YlwWHyBm7vicEbwbWv9JDL4XMxYrcVe2a0A4OIbI/
7bOmawM0CL8GHveOXZ4DTO2eMVn9mXftq/IVG0EjWXNThoVfVzwkAujIaBhuI1MeiEv24yZWifDW
ow4GsFwTyV08pjM9Yp2LI0qm3g66JFdyq2/yYj4N0hBndlx1l6Gm+eYHPldEowC9u0dHsuGGDlt5
99vwOywvNPIWASkT7f9j9lHA/JQp72fp3zL7ta+XyoVFRt1+vaIWvKz8lj8TbCA8qVomRj2fFSP2
t8x/L23g4ATFIwbF7WB1fkxp3ZxyVnuAiytx7n43whiT6d97XPqgfHGFztAdNQ+WWWeYXnSyecdT
gvoK67SGikZfmF/Mr3BlxV+Q59+lkGV9REERspnqFmnzdyWR7Kqo2nSKtiNTQdyxCVpZPc1UannE
/SpLHcn+rTMsFt8JeTJ+Lq9EXzERKRjkfFQkzJz+ZrmA2Lpa4cMKGr9BZnt6QXeEZOqOchumCup1
vxnK9JNiYb68FaMj0QYA4eo80GkoKuHIz9c/8qQCFP5l9KGQWgL0L60slpVK4YJvEIuQhfhzlRsH
YykxZ9Enyt5YXuj4n27XUk73LYOGM2qJwjkqH/2eMDTH/TPuclhRCiqT6CoX2Ps8dPzjmRNl6DQD
cAWTx1B3qIgCt7DhJaqJxM+VOLgASkeAYE2jQ7n9z/yQqrqVpiVbcCg78AdgrQKnoADwdzT8Eb0X
0/fLQeQhxNymisaCRLKtL0kc8S146RHp0DB4S6+rFvplcDBg+q7EU9NNFk0I4dW+LALHVGMPC4m2
HKqGZ6h811zEi6o2fS2PfZ20TxolNSJ9hhIrPrTvn8vpMCCh0e/cM1FDolr+HcI/Oqaea3gt5AoT
hk/kX04llBnOvuOkYGOCn/ErbQ79OOkKdG5yYRrHyHAdokoB67YZBqB4G/duIvL7Lt7Y+X9E9sky
1iCyNTbXI3gBkItaMt7zbTsRZLgyYY35YnAq+j9nskO4G95O9G7IsqljNPGb89H71esT35FwHRMZ
chVlfHtXLsYzGRqmx0OVbswpoNU30f78b1Odm1nL562vJ21WCm+zy7R6IL3PhzTwqOzKU8cURZME
wiyEltLCnPF32qBjNeqziaEI0Tn2cHFtqLg9iywJG9e3Hr5SrNA6jHinkoZnYmlSuRxKbcoibrFl
8Ob11YayNWPswR3PAO+ER3b5pqNAeLUjETL3q+x4dphsgImXolbD3YPUkKbkm+R8luxcPbLeAD2U
/wief6eciY+xRrbpbVPLVthFXol91DJu7zrtzMrPKVeuRDyMpaBTiNyNAtcwUK7t+CDO1PsmnHE4
LcK8k0xcyT8WqUIfVEcLBF1ugqSAGOYBFO3z9pjVq60emJaF1t00feuom/rI8VWXqS3v7pTpay3h
qXSAgkalFV4MiLbHDbW8p3L3kcSFHyAaiNyM1nRaTIJ5d2w1Zf9lbOhZCDTO2teFExHe1uF4a7kM
eZNBwEDZF6LVWeiWY4ACzMX8bt/UBXKb4F651cmjH8fkIK/BY0sGR83Rr+ZwvySCV55JXfshr3PR
eIxjQN6brYlmxq5E+LF7aeDQcmQbBLmITpskjqEC2N4xyOJd1X0Zxfda8oe9mjduJAC9pnik/bnn
jg5MJwFcN4BLhZLwZi8zFGyl5x05xVGBP2IlWK8cRpw+ufCvJPR+ln2Re9X7rxnFgWWuAZ1osKTa
OPNTdzJKlH6T3pwiICAh4hwIi+6wXtHSqMv5ARc1LG4nUk4kZbp3+tUCCWbAgHqqX96c/yDpddhI
f4d7BNoOiNU3cHc5xqEIjLucCcU+g0ZhRgKKc9bqpNX2QEQ5Y+lQxjLwbmkd5qjPPMvz7fHku27S
6TcahTD4HIABrfqVsPXSUa/Jd9FJawMxmy1DWKNOa6zoDlfD7rUnBzxwlskLxz7j8Do4N/f1YceI
fCVpeK0b/I+5VCb/8Jsj+tJJJ1e1ASFqYuTnGpjWxqcuamClvLoG9V9MXNzRFSzWdWkfUHuoTjUy
IEy57npLO/OkmanIuCOHTVRs8ZmgTIEmcnIE2Hf4+RoL24svKeUlP+KiIz/3uKr4I5DV0MCVei3W
gO4PU10LQv0sClu62RmLbQ1oeYXLOc0ZRemv1KPZ2H9ignAQSN9JgRhlYg08uKA0c7Tyt8CJjTqz
P+bsWGQC4cUUxEI2cuYxi9f90GvbQ77isG8YEgjN4k0IABs5IzXL05W/h4fYplc3Ntk3uDF/DPIx
Vbxab0LFQie73oTq2gJNY/YZaQ85D5CV5qNcQbMluoHILZFatN6HNCxoZQv9PrNCyZ1LQLzCfmOH
Mnre/hsdHYSkji/Rp0GePzTsM00JVYggIqd0CFg4FGuTNUkCOoEVJ+gn8wJAHK/s0iNegbbjNSL2
Mn5JivyJvduKnZphuoycQGFpRce5log/gfW1AY3hhQPnN9F1gw//sKsHEsa4juSp1Jdx6NQ1x/hy
VUfqTO9ycK/mzN1saw1QsNxmbX2XvR0auAQ2W4uq3RaCTdfZTjfQR4xMWupZkZG37whtuHh8zxts
2S8b7Xo2HlVnIBDhMLbSJOkARgfcTuz+Ber2nswcPoZ1jE7PkF6wKNDnZl9wgzF4C1w5lKi7wu0O
FkSBe/N/bfyCfHMjRspZCoKdHV0rB4tEHLeZO82xqeIlmDPGc0kUoMmEamH1+cDVtvlMd003CxuS
mN7aK86Mx72Ju+eAyUZ9RO6mPGszh84hCM47RjnKhsfWE8qyWYBVcoKQ9gSHN5Iq6X1VR99h6+xu
vBbQJ2v+0sPWrXMoO3CPywHoDO9Px7z5MmeNuG5XZfMpxjUElobgXufFCTuDKSzrtXbdzUQvCwP+
Ql8tFYJjG1vfiS04L43nEoDlWingCJJH/l8sUnqpNKnYw7wEmcTutH5PMV0qddvtqf6dliND/9js
hRQPjgZQI58P7tb41p4nW3EnZb5rG1MnsIExfgu/NLrTejp3AC0/PQuxT6i2EXjNmJs5hLr7Z9FU
NAbiP6nWwMnC8MuOo46bRJyjNB4EqAy/t3yhy3Bt9gN1VoIZeDdzF+MWyaPITSncFOmfZS/zoR00
gVtGjGPXMnEkbSNgF06BF98n4Xy+O9+NPis3+cS4AUwKY02wuveb4k9sLtXHZxmhN7tvnsI4lcSX
/r5XSMMit7UMXi9RLk/QQoQ+Q1YeKC/WxRMxgHwymLZwufyqFRFzXEKMVESwDOF0g+gOiVxeihKO
3ZByY2Wtlv8VhM9+HBQ2BS/U9/znzgoLfKqNWDWIKWbgQdfA3ucKttUUnkOJNDHin2okKu5nmzEY
Ju4hkDC9WAMEWMHqfnkMjq/pvrRXvJGHFX/PFx6XU+E1/Jaq7AQiFGLHhcCkC80ykgKLG9ifGagY
YBrPo2RoupQKZ2JB9FjY1a6wzyoAhbX8G3vnHorrTxzNC+T2q7FQGJwzL1CeXpvu19LAb58HCFzK
EBBqr599LgMhfinbtYoSegEHm0/nk9Bytpg9WrF7Mw5kWnw6bnie03T++0YKpn20+wywzgv748GH
bGNYQXTNyvT5XXiaAw8ekN4i7KgZcuiXTEMIZlSphHV4HDKAGzmgK/6LEgji/93S/Xb/xKSU5pvV
Vnw+aKx0xLeE/q3143WNY65/XIWd/H+4SsdjACYNDDNdCWmzk+CU+JRU1CALek0MfkhkhTxN9DLH
KOnBdiPHYurdXisIBghwqqZiAzSK5loKD1At7xAZj97YA32dZ7OfEeN28xkgrvQxILW28dT53w6B
EtMZsELo3ZfbqaWx1k5tX/hsIby0q5ZNsEKuKnEPbo4nEifxvXalgrMborrOI2Bo5iU/YJLFdn6v
rroiiTLC8mGh1ebXdIKtdziYvnsCf0fNPen60kOolAI9Eg1AkIk/dd41s4KOjz08FyOuSb1GPwHY
jO900xQqcJzO+yAIXLDrBQKU2KfzD+2ZMNsqaLCcszMZd60U0JekAjVY5wAkuEHL0VPKZ5TlPnwN
o9npmB4yyYvNmzo4FZZ6VzJHQ2JynehyZ3lulDSwkRS586CvhnV4Qzduq6FfrnPvxCmWxX8y0XhF
viiu5YBl+SBja8ShTbi+0hexPMnKPguPu70sNv4ZB+r2n3Sc6f7tNXGiRPlMVlJKPU+E/LkTpA6Y
g8nxKY7aK7NX/4rtwjix+oZtCTqwfpUwBp2Fx4gnssQTWcXInaJI5MeqnvnF5iT+soncOA1nmBe7
blQN8FBVi88wL9mrroJefpaoLg1WeZgbdoVVaVQ0jPLGCPnshzSWn1+tioPfWChJjEQSFTzhajuY
YDtvjjfx4zszmsOnWqjjSIlfqs5I0T8PptMi3zxTkMBCFAXRaGTxmLABtyQxsOmthgO9lrFBkscP
bi0ssOXP6KUqa4BNWzCJXLyPX+u+6gCerEOQSvhMNQrrTDuo5B/eaN9gxCnmChK090Tp6gpSmoDw
64iDoCkYyIRwqAeycQOApviAfjPnrSFJgc/bjVI+j4R2mx5ajqFJcUf9EHKffo0ZSn8Ocq5b6whe
VWPutZkfvGLla+SR7oLwVANk/01QvaNNa09jnQOnkTNSG7K4ymVVw/Ogrs4+9Xv1xQihv/b/MVpL
tNXQA2E9siYbxbbo0BKVYvAGj1GN8WN36ZrNmHk5RKdm+ngF3BorW4eUiaboh32pfkGqaQKJ2BVg
XTi8Aa2U1JOa67JIiL42kioTJV01VQLAeNUj2EdC3R8PFHsFRxJHmdA6EXwCSRWxKEUCZjgI9W/P
nZRSpRBpHX5UH4VBB3RT9RK2DLmTAhPIutGNJHE9H4dg/V/PDpACzASiiIhyZDDxcB0okARz94J3
JftHGIGPBaTuSJ/GqFDJO1ld7cpaiCDQZQNY+RMpwsO/w9WByCqSFQh49aaxrBye3ixWlfh4qJQd
rJHisc3J5k6D/FSp7Hk40oF3BugWMf8gz/ryBMsQW254ZmTnZAqqqvg2DAyHSLV/KB5TzqammdT/
uLNHr/ACroKUQ9JSDheRvRWy+A1D9Sa62nImViTCot8Ku6S0ELYC83KI8eHR86ip20QbbR4W0wYY
gc4QYQSov+oo7MmZHAeyN+2JOi/kFfXkupeMCeT1Lv3f7XvEVb4Yt6ZWxI7O9rBGGQSinl748uv5
ehsfY3RLClVF7EEWdT+dJuQusGNfrUoeiS/sNrNyd7Wdth7eAMz8Rk24o9sN9QK3AV77i4V5LVHE
AuTjOnLsDYcIzkYDYFjApOlee6WZVM4ToTuJiFlRBWYWjeky1YgqCex+w5FOL+/9vN0Zb8Aem504
AQnxewMrWZGPZCTxzG5JQWdyc/AvJXrFHsU78sV+k92NjALIwX50U1Es/po0SkSIShDpedhgZY6w
h62xR7YA6AJ2KeLwqWALepfLtAsQUgKbpZlRD4ExJqi7hWxffAy/uozf59yy3F5fYI1+Box3HCBS
BZHr/09z++mSS6XMvcNcqv0yiiiIk/3avEY3u6ofTU3y0CaKAxrspPqaEhdB/TCR7f2uGOlLBVrV
jQH7dUe6ueKJ6PrCrSLboGe0t6F7UXewo5N9R5Vz4sFVaNwdRlU2pndB4tilEbEDun4PpGDU9oNe
FZ/InmWbrtgFDa8skEZOcPMjkMqrPUp2MSHO0n4QlatVtV97t4K+OU8VTNv3UQFJ6f4ixNiH8pDO
CElMShmvqCLAYYJ69n96E0rpgq5SjDBzwdiWSpItxtMRwi5zOOn7ps0PzP66M5CfpSBI8sL9rbZy
FSh9BYR9Efbke5yblfr4+ks7GKUIG76e9EoXJ/TJp1I1MXozLiz4T9BC+TBvJt6u1+0Z8k0VMS3p
7vsfPzEVpBw97XsjQl5tIGhjz3JwpzXPxT66N2TLyt/WSsbaMxAlV+WBKpoc9qz8xlWgkxanT+EH
TtLfomOakfClj6UhCoqAEKUucVnvMgui6trMN5iFy+nindSw+1gEBVE9L7goaexYPA7ghp0g6Mp8
qi1tBu0Gpb8vA00PHN+Wf8sxSoaWkxYhPKmyA1v4Pbl9cheQ06s3bMLGo5G3vQborO67UeAxbPSe
qikOK7yMcyj5Ff5gOX544wQ4NM2wZRXB6EwqJfjX4kqTmva4PkY8mVqxUeqsRrA96vqoObDir2PU
7gPqVK6Gyp0RYTfwWnfqth18yiyLY1mIWK36d4lh66Si8gIrSVx2Cw5xLznERJV58uR82yNVQfZg
IdgYxbzglzXd0+qZDOqOGFKe43PKMx9K0akwcketpvMbsZAiQLOeo9msZi3c7FXfP/O5jW6ZclnG
ffh6Zg4AqmyNHgY49OdC1BW8LlVifwtYuULlYWem/BzCXItkXeQ6dgekn+pUZrwXDRV8wI+vQLEv
vIcXUxubTttA79dSBXyq2cvojl49dJM+9KeQr+ohbO3+KAEtiFIpE8PDQuuV8ZJ8KlqrYsV1zzoo
BmmjujrJgOiyTVTIsAXSV96zSBFkXFZorAGTLUaGWhSxS+f4PEfak+JGcPWweJVitpSoh7JehBPl
UUjTI3iEEaVKVgRIMxyjJy2xhsMiCA+JCBySf043kPCkgGXHSQe53/HAGJjqkUCnQXQxZdn5zVDG
nN7Dx4rfasFP+89V+K7sVTFlZVeeOoB8iuBt0xCi8JeyRKvwHoMRZmDcgT3gkLKVVzjfOwg0Wtdd
I+5QRwTcZEAE5gGpvuOGR7JZUqxUhI6bstQma+WUw31SqnoV45rViSI1U/HTtHbZaJmsVfJr8mDp
Rq5uB5gZWmCbsHDmabCqmi4zxmwT8xEnONOgvkmJJb9H/sIESWHE5Pq0/Kj1Iz8qxX+0/6xW9VC9
/ZRCaxosF0UFMGl+ZGZMsCVm3Ea4SdzCRn/em11CrbgntRt2Yt8OIK5NfZXa8mF/wC0mA4KWRqYG
Krip75C80/8lQobjqVmYtv7bXqUXWLhRYkYgPOq0x8KJji0v0h7LNqXXacHSryS5G4wnuIXDPI3l
3dMvaWrmOFLzFCNNXdHuBJ1P/36p/6MDsy0VZ2/SGMW0QoYNX9BmDVsedErWFhF3rSU7Km29MA8n
C7hWjz0XByp477MNya30nsFm5U7+Nbf+AxAJ7PMYQtz8/DG/dYH++EfEXBB+z8Nd+S12iP+HR4yj
PiDLXoB0C/emiUa0ScI6m3Ds/WJIp+4gCSyKo5Y/r0xqklzz+LcQ6ZqsULFvJNFfl7sD7K5npjdC
YjiGEjZ3dgZ1wV9Y7Po1LGOQ5DaQ2I+RkECl0E5Uw6SKX3tlryHd0B3GG9CNxb9eNKy7HfVacnYw
/R+8P4Hw0pvOmWzEw/Re1k3lcfCFb2kifxGF78SL16uJrBa5xAMnDii8Xf4qTZfP7aiC5QewoDpV
3sbAZtqR/F08CvwUrgd7WY1Ht9VNHxjmpsgcBajZ7y5OoXNGmki3NbyYftQeNclaIYht2525iyV5
/sbsHiEwszK09H+qsKSqAQQE93PjuWvSolprkppIzTPvICPmPN0Krw9QO1fqBNbgIUqI03MCoYGc
NR/DpC83GGIVbjrdI+oY9nEl3K591N+3kqcR8G9A2Z3Xnb1pQNz45I7dWuKlzVpyOYPdK74RB1kR
W7oRycRdXxCji7Iri9HokKMM8LTtKGrI8npEM5koT0Yl3H2kSybMzy5DVFwZQEBHcL/C180pUdD1
aIVwbIdak/fcyBtu/3KkERb/Qtw0QHE5zJUA1neGJg5U/opzX8SFL0/CV1FzG1ML7kr3bsTuAqWl
7Km19OPoIr3O0eolvVpcohYFH6jK9QPQ6zd3sEBMprb7o64gCH1YngDsOnBNNTjcosTAAh9dpwoE
Wk037BgPgSWVtfxt3i2euHY0BpabrMYndS6rndQ4rEHh6+BwKdYW2WOe2CSNrFH2bVzJHCV6nbr+
h6uOPnRF5VkNH2RYPyiYykDRtQNzVLNPCBjp52FZFGRsW9uXNML/MrRckvkZ+TwyHAMrkGN0vQNp
mz+223oDa8FDWgRlg736/77T5UFo3UJOrVokv4ikTCwpts0254Y2maUvuWMskQy0dDeF7n2Jc/jA
72qXia3ff+hMdUFlUBPRySinqwlOeisbiVBg/rZ2wpqkOjtBe6Spb+WO8fAR4bnmmaBcoBEoaG0l
8TelEsHC7nHMelfqD21mMrQFyRWvng31NgbiDLbdHzRCd1p52JIwjaWq6sl5d3v5+GYv4RJGEKr4
ZNLN3ktZk4PFBsgNwI0IQ6CmNNfENrx5FW/bJkNi07/zblKFz4JojPDQJAXr2J8bvhTs8r5u6Rpb
uWMHXOsmyKKH2H/uNjl7tUcR8BqWhNeyTfqxkLe4/ntsnKYWFv69b/ZLywbXeROaMOaqjIYRAvVu
bNbt929V4T7e3/2o/CSc6tJP2VFKwv+j/W0hZDukj1ExskMbvts4FKmbTL20LHZzptE2/fiFWylf
gq4Tienz6ZOsLW6JUvQQ9DYuWr6+Pc+naal1KKE7FuJzX/Y5vVdmgs2Fp7tbSY/Q93Zbg/w79WMB
LjR8TnP+WeYkj6RIom9GnkbF5pjC3/D4jJ+sVLGtKxQ1e2TGDVUI0FVmeEIEGEx8AfzTIDmVOABo
UD0fVKckBhMUv256lVK5fIPR5pilEzscffEUlSoXfT2SYiKXml8oV0sBU6GCVls9SQN+GZcVjG4U
tq8IFC9lajNhWMJvXDIlyAlCewPr4Bmi8dg+I1xxlZz/zHd6X8YgwssonSY5rsf4OnubRQyY/0oi
uEtrk3zSvKGR7FfZie7TzXHSemAIjgC1XjyCUVVjSWtZ4sGy9An+CRHEVR/ebq/r/oNYE1NhxDgF
YAe19qcqVXnmhl+ho9c5DjzPPIOtopCsZ1Iu6NCgFzD2HJ//4ryIx4NUK2fd/YVaxf41FeulOUTW
NbRBENgg6XH2zHUVSLbdBvw5YW5wuts++9gGZWfArC80jFJbiMIWaP8z2XyrI6J9QwjXKRtjv6yt
rgueC+FyMdYhtEjnzXdKY7rZQeu1EtMpIpYa3iuMc50u+ONvb8+rMxxSE/x8/yevm860ikf7/eAg
MfwPkzDdyLLxjKYoptV2jsK/xsSnVgZ18dnMnTDkVnHyTu6mZxq7VqMP6tWJF5N2dZKKFoV/P6j0
GSZg1dyCmi8ZThq+Pi2TGzk/Z1LwcuHCUen6oO9ISGHhCj7ZjiP8rBm+TOTaTmxEk/Zn9U/0mEfV
/hipRiE0Ukd3r88iojFjNDbW8cpuBGDodc+xKRsHzuY3nB5yiw5RL2QsQw0yg8csqk8aDWUGyTT2
eiyoS1TXVx+OcoPi7q8Iy85NS6pcU98Un+5l0S3jbTHzBWBnCb1KlLMpCfu2Wi3WbH8Nj/gd2Olr
hl+/mz/Wb4ghFHYpH0Z0+0nvWcy4mn/ZlHVFykPWJ5B7IKgosgklKuWze/lAQlcxdo9kBqVOaAIs
dZAIA1jA5qHlrJqgcf4zYCpvzJk4RMr4fe1h4ahxeMOD600WdiITcN4BjRsF0ocaAjnSs98rVJ6V
OnDxdE7VOmTU7atyVc8zK/zs9AFKpNBgx3Yp85aOeHtkRoGOE4jHnO9loROU1lWN4Eg4Mm6XoKNR
5oZSeI5a7C7SyQuYX/J0nKIwA70Pc7D+HeeQhhGv/P2wy8YPhF61Z/a1ZUPh9vn1d6q51LMrJsA5
Pb4L3UyTBeNVs8QBrTarayZKXzh1R5+scu7OY5gom9Rz+8DRM3zhQYMGW8ZjdwT7/P5eR3O0SxY5
F+yjQG7/zJzr7FoAz9RWx0U9j3uIMDmnzG6WKx4MqXSUJgq+1yeiuQAS3lIp37Sbp1O5dBRLukYR
Dt8RNi/SS+ahz8Vd2NkRDYhUZXgRKV6wysWADOF6GVMe1e07WFwpM76CqXl8fgxWFXIclxfMHC6u
MCWrwfigoOaiMSCmMi52yu1OZbfrMWMlkLRqflPXh8aLSMXL9bpBsIoGKt72S4fjbC8zSU9QchMA
cLKQlpA9fonuAYt9nacTEwJuqKtLLkPthoZn9MW9tiaPlG9z5p6JQeFi+0cdGxsb3VGTim4IN9Iu
R+UzOsknOazBMNMht5a4UR6yvPniaQIBYkJNEMzFJUsgGUOTV4JHMpFtUT1JUjCf/kfRoKwMrMVt
bhKf3lty2IYoz52DKJ3fHfzDQQ3sy1SFO3GjthDo/wJWyJLp5xF1nNS0X+An3Hd8RqYNM3yA7Cru
jmu6ObhkCOnLssIa/A7JhYrvJZ2ZipSVu+HTKGWAInqpOn0XnJahLGjHE7wNb7bdYpVOrasdkUP+
ay6DeryT5iEz/dbH4i8xvFmTXNDrkfqJXghoEKjwI2jY4GGs381F3Wtdb71biwfa530TXLpkI/v1
6ts/W37vw2wsXe/Gw9S2d4RUeoIK0krL8RInxltUDKLeaHoVpTfpyYDt+CXF8e9j0g/VAAvd7gem
tB0mhpe9Ibma5gP7t/QUUTh55mBEKdKzhiquNa29D2JkPR3ms+x8/jrqOHff8on2qgm9DRGE3KoR
6g7r5fVFpp8STwLEH3bN9auseqIROE8EWmUutGL5nT4pew/1hD0IBSx69J/hVswTlqtQFNzoJW5k
uyshsvPnelEpWFPPiLZfXGJOjgjdaQLzYwkYqg5LLflzGlld/sW7M+tDQbnWJY/laZcQWxpVDE35
HcEJe6v8P1j1mlKSwtk0h6AWPoAI1voJe6Vq3T3XqX9wWb773FTaojvyB9KRL/+WYWm37cH2Mu7k
qP5i30KbhV8S5cA2YK/arxCIWxYgqjIO/wGoePZfrEyQ1DFbs29vjdmHjj5HJ08/RWrOqcMJKxyG
KTCz+rpGgrW5eZyRuHu16tUcMBR+4L5g4XNLlFyX8yUCvniQRsMIgSBQbvaN5wBuNtXUsAMC8GPx
C5Dz8c818/zgfQ6lJQDv8Ibe2y44JXTkreN4PnqXci7S7w8a8FEiYOZHK1tVShAtE9e4xGWDIFUq
ZXAtVNIi6ZHCIQrMSR28f6KMJsRZM2HdHo/E3pNUCt2bM/UnqpXycdrh2bTvhUVcBb+v6XohXrWS
8r9l2Jo9aIQd0b1yp3KVFP3QOHFF4EV8FjQ8ommfVI8bi/mUkpzJIa7adcsxaUHEt6Tr2rH4fBL7
kXXIFnzAIarJn/FzUb68HJVcUB66GCShAmvxmQ8BDouIXA80eotcPJXWsqAVPzElxFoU6nJNENpX
JZK3pbuqOGxlceFIYHudk11Kk4SlWAgVFaakUAAN1GMkueWRBIk607ajWfBfAPys6LJLMfC0s/wh
qJdoTNttj/8peloMwP2RGjZm7HWw8x12ySWmzt7u9uY7kQCfmosR6WXhc3G5rE0L499I2KivzYt4
8bSigZZklG/jWKDRYZWvHSFuxhr12nco35UhEyBixZLAmSRq9/3QeY1bef1nszK2oggmQSkRP8iZ
JlCiWJ+FURQEfwmztxPOcG6gELcjLq8b5Dk8GbanLyYAYGZCeuLI6BgUgIbfme5dQf1fAXw0OLiX
VgbgzU5l9XR7fcqqV2I5G3QNDBCvJV7Ahacz+H9UEhXyd1A1MvXsQK4zBx7g1pweAquMOznHIBwU
6Os3CoAsX6JN248B4oEv3xVP6G4sOdH4bVLwKne1dLd0c9Iza2U55FnpvXJlecCqmaolbP4Hpbb+
kwQs0GwQDo0jozDT1weLC73zFW2vMDirjeVXU6H/SxflDiNCmZdAEyzt9Pu49XH31d3QG98vP8+l
eXRzFT9Uo7jRgDIWgsQb0IL/p18ihF3/GcSao3Q6SyG2gwG8gHp9GiXDNxxaxsL570NpaSv0Z4yj
rn5MSLJuwROC6z/dVC3chUjFh2s4JugbReOJTDV1Cj3zRp0gm74sk1ITxmPjJkiR4aGv1KEt3zhb
H4XRgryZmEWRS3+RsL4JBkt8bvgu4ScvJDy/4fC8381PkvOJ2H3QyrZ7Sw+//hN6TyfI+tSebOSW
X6sVoV6i9IKNum49ScGUK7a2Pbg0Go4GuoJhaRuH/Wr0JPtOzmSd2CuvqGCg3WcwBKKdTBizXhew
znmpvveCcfzIKCXdy16AxbE8hLOcbaQB+tUTaqShlnjyLBQutRPhVZu72sWUZWy/6l1i1X4hGRek
7P31K0Zq0pDl+fKd/+YXLoYjCagKykpVEA07ooy4InnGl9pxZceCHw08vx9WVdCZAflwprz+jnYW
9yt+MhCaw9mMH5GAxtthtpGNRlaLf9Mza2AprdX5+wPxHsWBs6NEWpHvzWHwwWQXHlqPH97TiXBI
4ACBcMta3hQ/y1rReILNrWXaCTWteJbDq0OyS5xq44hLplgzgXySdNUxXAHuG1+UIb8NrLWmwElo
O7XFCrzqOZLy56wnULJ5b2ev9NbGFDrNaj4NEMwqgIKKnQwpvnoe9h52EziwHrKt4Lkal+utdzkF
uvGy2wRzEZ4DpSRghLT3Hk4TxhLNUvBcPRHSpmwUFjw1liRzS+JDYin26d4E7SRa8fqVnuijNgOs
HzCbm/E6LVTRYYnEVYcBWVXRgcvdvcrhaMM6hNpw85f6T3okTOXyv29AMW6f7A59Zn1Hfig+2o9q
yW7uGpJtcLWT+K8D5hhQNDmhaMR44uoAZPamL5ELmbTIQvfZc9onRi4G0mMnhxRGhiHzP5ecO/V8
jYC9Ow6gPD27jGI9nVG3K6aw1jOE7eIEiE32KPv4VnMTFcV63N7pgGcfQhvZpdTQFt1jQqdUu2mq
FW3Kr7IrXMxRmitwGI59SUP8yMsAmUvof117NOfH3GxQyFvVdRp3jDq7IkTFHevDOPKQqOjBICez
6ktR5L0+JHdRF0NAiV4UPEx6jrLT/4b1+04P6bklPcppsgYMip6X+KZnyire7NRoLnRdqDKeXqw6
MqhTC18Zj7HuvhMIxXoxES/cpUW/7U33qHcGGQKGPMxtQBMJRydZgUYBWOWmWaOoyO9+tXBVbieb
NWkTCbO6EuqIgrEp/3uNXUUX3LTUPKrQ9o0yFdOLNtfeW9FpjS/SAmxGSWTDiZcUqURqXIz2H1fI
cyOPiDyBpsFq5TPmJdZ5clr4nsfMn+GzQGuLkZaT6v6S1EqVM/6VDm6fRd2c1s1EDE1BaieIA2cU
R6stMn6ioYtsxNiiaGymKuesiw8itGByMMhZhxmpwNVFo4h7W8wz9an1dqll1UL7k/01xcKYuAdd
lSjPj1rgOm2UF0iVrFijDQ/Z4gDY0HExe+yp0JfjoCIKkZt200cO6MsMIBao9AAWkZ/td9nT+P6t
+KFZ0DUtNXrae7MSz42WONhMZ3KBQgEi8xw+fsBMz6h6FtOcKCe3XN3PTUEhE1gX83oEI6n+Chwz
6wdrVGj8GkWAap1fi+ggUVlP9L9IX0jwBRSaWUiZH8mQS3ci18INdOuMTEheFneew53ijkzcGfuw
/6Men5cOFjYsIRiBIq8W76SDg0HyDMhrfmoqisiRBIR7RTGfxBDiqhAp0xOcFqAFngLyKhw1O+4L
WQBO4mNYDxQ/R975XFC4Om2kIoYn/Bc3kfMB9yqNuwMZp1SvrJyKbLk8M8/qDVD8o30eOyN04lIn
B/qYab10nzk0Xc4OO9ImQKXqDIU3SyW02ygSqS1lWb+Q9msFoyg+0vw+S0+VhZlJdGylj1aUdmD/
fkdlvc2ELbdQlh7J57/gIvhQjrpwVtXwXAXclSIEggiJG9Ql0yoDbUz+Bjl+UBEN27RPlWfX84Fk
RmrxDDrvN+YHRuKJArPiz5bcUM6w7A4SnQiryc/WZGNpdZZHP5Eu3sgkhOUaAX831ILpmsmH42Iu
xjO7Et12euH8wRW7MZNC73hQLI57h6LpAI6bvcuQ3MONs+xH7uT346paWbC1ya+uAs1BN9/ShkDP
is6FNZYrIxzWKSzfqb+ihRYjXsEX9ViEGcydUdDrp353b2ALg/cIKKbnV4xQiCgkL8+zbu7zhCYw
u6Lmib4F/KonBHD2RkXTiqQavAu0fbgSv1rBLanwYc4kzlnweMxKARFkcr4YDnW9tuEULIJySNS8
vVmWlJRZChuN0RIYvbd4f4GdvxHdutswnVdVusMHRsZnz8x7npldxRG3cfxryCVWFJbTDsoAtgj7
+po9qmS7N8E4OezxIYO4IfPmV43lL4kDLrCcFgi8jGMbJ9ItwVtl/WuFzl3a2NkEYAOJ1zo6BWA/
PCdEszTZlQpR8PP7zAElgOGFfIXXgXdB2Th5w9zMW13aFD9zx9GuO6iDjzclgb1Lq9cKdiIsrzkX
cB6v6ryQm/N9XY8Qq9GlNTKadZQG7pZ/ff/3T6ZWc9tuhAt5vueqZ8mgEuPrSmvT8eRS6JhFfQMc
5W6iaeXcAjLQZRWDP531Dpk4BjHxRRsz7T0rWMZjF5TvdxuVV1/6N7DWW61vgc2roq17l/8zytfQ
gkQeOKunOdEZY75ekFzUnQNr8BjQvA30iLIfhmKUknYUha0iljMmuo4yUSESXXHxxsyBlB7pfBHr
n1KYA1532/ifLPedCok5pSLZhStg6GcNovMPXJGhFbgrBmraqOvUuCZOywVkpx5CFOpvkNwCfXOq
Lygjg8e99T2pF+FJJ8hHqTbUDnpgPNwNgA8dQwWjymlWXSR9GPwkTYsjA+H+N7pmcIutrIksE15M
usT1d+CIaoDW8O/Q4x393W35seQIE94dgiy53ReEYVh2v7mH59uewQ1UAP1s3tQTcxhWAEfnglvK
euwc94YcWrgn2OS5SNdOd3At3rxbCmPXC0AIJe4j3S1kN8FlaJ/CnG+x6Lf2IVTbMihqMxAoKwmD
e/5ePViVpEXOn4d2HEoL1D14JGYW09Vg8SANLgIOUyzM1mxBzeoxfund20/Q7pTO7E2l58upSakq
TBibWL++cfuVQYiqUKSgrKOlYBqb9rq+nCHI6ZnEHLb7GvelV2jy+onoKsCzCGVtPTtRNILV74S3
DN1d5VmgzVSxYWzKeJg/wBgfwEQHrShkmDajrK3XFYPvtghwVDT1Yat6X5ZEEdYXgNHxaVN6uNMT
CA48m7T5TIWaBaqZZLaMoTAAjNiuMRm76P3Pb2lwtDJyBjU+t9CS7ggO+O5DnizC1zLycXU6TPok
v7e9nBXPFiTaY1Zru6MZoFT72R5Ksig9HXR3DqopZ/U9+BpZp+HdVS/BpckMzXZV06sukouqLlk/
M7TNUvFQ5WaMe7I7X0omx9pOe0/xOHLsKaDkjLuDrfqK4o+1l7vqswyA2wSDV8Baw5a0XjlwtzSS
2RXXFRPdy4f8FyNquu06p32nn+uHincRsY4WIfnKowvNW0gqk0Pq06vYHuLU+5rhs+766EsVZ2TX
rcWfru5JVprK7CX1yYjsgqo5okT11g8UDLlztWTn6fPU1zpo6E6F4WmvFHF/1ZdQhAAaljahzt8R
7Jy/zmc4Jvxv2v+n/XnHqmnbEZCLxqlBB4FusuygUydUlc/ZzvNU3YU0znFMeNU6YBEyd3sJK59q
rihVsU5t12MoDfnILsNVtFNLFu+W7ilOIB4Tjt8fuuI2//enjiIDjwBlG8rc0Zw4pquPqkpX/BzP
K5PMD7d2JhGut31n6oJUzboGJ6xLt3wuhTpLLUwchK1Z/eqZLKumpFlr3zzwE5TtCnhu7ITVq1Ra
vrcJbioQZwR2X5sMVGuRj1GXo1C6Hr5gqeM777gCQpL4vvc9ukoNWvsi6V39gyDOB4R2iEQK4aLX
dv/4YRHQXE4EbSQ6nNG1YMNA9WquiADHvArbb9Xwc0+sXeQmRN+L0ATiAH2UHRbmeeljObMADy80
MqoW3qXbisJhT/wB41I7ED9fhRwhuM+wGlsD9O1mgNgmonLdL5aw9fyjWBy9uCMQcENc+TVFligl
XqptKcQP4DRP7gL+YO1pSdLVb4neaD2p60dTplSOqrzS+CQ7Q55zpXA3LoNexZil3lQ67Q1XPKUt
AZBxrUQa6JUbZWwu9S8y5lISSstvlzhKZ9Xw9VzuuHrLuFjWYzIagDcGigmrjGyKkCZQovPaP7mr
5DoA6lqjnTBmjnMPN+58B9GxJQQWZnPVzpF4wY5PxLjoj0iQVjqIlcIu87Yp/Xds1fYw7Dj4IlGL
8cP83V7jrsmuGnQ0XatGAm9yULDb7tgshpwt+UTUa8wCnCTIuL3Bx6EtwljogoKPxg0yDtkGgYLF
mHcLOzN/fIoQjNRxBJL2A2hikv2eJbKM2tOAk834R0PTADn0Oxohs8wHIQiaBSsOgqW3eX0rOWQN
ZNLz64sHU1nGEDJYGwAqRwEvKxcuPRm5ONLCeQO+bS+Fcu0q4Qe3muIhmC3tNFxla8sO0IOG8cZ2
e7iIIjlUcMZzDrahEVxW6saoS3XxjA4z8Z8t8G174RdlOFkV74ljmazr3d+aDadnVgKpE+Gtn2dr
BXzYeBkDei2Q6LNQe5Mo+q8s9UuT1mo821XCDirav5bt/mSWAfdd1RrMDxX+AvhX5dw829kh8z/Z
xPLibGLCIjj/rqU/0HPRfAB1H8yF9JnoH6N80cIsQMkwCDrTGYy8IZgOHO4OGErV9m0g+7uPo+M+
CBJSwgafWWSVB/+Eo2ae3tZPmijiwldPQiri5SodB+SoVsAbLTGDMspP6x5a8j2cf/Pb0iNxcwSP
wRDdSPuLG0Wmr2o7c6Ql2YTMeJONkcavpKlh5t8JHLZW6qFlct6atVLmD6aQGgxO+bAEUQKuaeZt
FSFZIy54m8SSd9Uj9Y/1qnYOwEuZy9nZTFN+yQNrsaDZXn2Bt50gWcIe5fWReOyVAv4cKj5Gy0XP
GXSKZ/Bc5HxMEV2hEMVdvn88euI0g/efJtNymaIzwkzORFBp7KIQOHyAZDapD1O3z7KCBu9xTKl0
QqwsQAmnH2qij4sJoVe37vifB9y+OwLOCGlVesa8ZZSkkZ//lMUuvcteBHtPAt4Ji9KOjnF3Yq0o
t1eUvO0xgw8yBMpD78KviRRJ252eLvp2L5vLTkrQhZK/y8lUinh+N5W8yEtMOOJqaa80+kld1wIO
Z+86yMHgKl+6XdD04GpDpb/0SavI3kKmJiUxvDdVdvs0rNNgadA71Ze4BZ2KiI+ppjMY33MDhI/t
dEGgCbRnuoZ1e7OJvcFQt2JXiTQEz3pNDLokab0rhuzqC/ozZhAmnh4Ieh+YZKyv6g3L5Mc7Z3bg
uJWDAW+bhx8duZH1ycaMnT78gtNP430cfFS89F80Edxjgfku2uUQLLgTGHMyc80/0Ub0N9t19QHG
bv9UgCCCuX8X8yYXxlRqe2f1llKVoxDxuHbBNa3sMzKB7qYqgZrEYO1uVb47VrPHaILRUPaF34nf
jo4Y5tM7WeUMuv9vjfduXRcFy26+MlO0h5cNtwlZ8vMKqurNAlHB3NmQdE7FGgaV7mNMDDmzDCUV
Wb9yqBPUmhy/zs93WZCSv3WNJgk5kBLYliWwSMVXSa5Daigk6w0U/NufNwHRuj/CR+wh1mDDjw7x
uBDYvHZ7+DmJJ+FaTXdpBJ3XgZZhwfpe/mbhogtYcjsmo8vKyawVLW/0gLg4IzMlcBARlquNf6SV
G4hQmXZGOuw09DJQM8EYel0XnrrsgrA1lpa9pMgpgQV9OIKYHc2ZfMWQgaZ5BBssj0x9Ul6nGt0D
DEtZoA459EYd8tNplWOYdZ47/HQL3fm/Y1fAyDZKi7vsK/j1J+kZ37+jk+RrlPMlFntjpR2xqt8W
blfb8W7sFW3+Aae3De26IajVXhWFAhJTmrxQTvq44dVeu1gYjQ6r3n7TBmxwX9gWu4Eahwg/9SXC
EFMfonVKRpKjhujDr0gij6yEkPoFjJU9TV/fqCEPKuLNY8ytFpyNb0lPqUMzmFdWNR7uLchm425q
mDrhc7/iAyus3CXOpIqIXg1Ie9AIvqKeUshVzPxRE8kjWNkSMLEzeKq6Ueovcxd0f875mrR7RDTQ
C5K81Y2kqRtt1VzV65IoWDi2ZvLwrCi+ogr7X84AP88r+F4hXP8kxVsxDAiZhX3OhM7kJ7SjBikp
TSmowM4Ep1ryBeJ8L1OISwYY9XW0Xxqeo8cO7+yNs0KFrk4GkEpMn0OSYJUsZPNH3WKUA7mlf0ew
rZw2ofdqe3OgsB2jolSVznUoSUIBL4q2FoYynhSlUKCKNDbG0WJQrvzo3TFdR9WYTWadssDaPl7L
9vwFgoaPl1xZ1Z88dI6BnockmS6AXKAvLdMS4YuqZayxPUOoLVDpWCAM+NbjsMCZE78hibs41f7H
D6K2tJ672ZYfGJ98aBb0dIdoyVfCKcW0RNPTuk9pIQ6iUkCXpGz2WHz2XtEpGf61UYPfoPVuME7i
Plp7jCzbdFKOTmcn2vfA4favrCbVIOoOmHcxRm7SC+4/TpReyoBMGWK58hFEYb2rAj0fSzOqXwcl
Ih88wxYomXd2+/8g+p/EeAnDw87ILXHhIn4PLL3D9uEhrdwXyc5jRVfCBC+ncNMYm8dkTdiTr8oM
tm3nrPVuBcH8VyrtQTKm1RiwLxfe0H5bCv1jNU54AQgBh6zFAyREd9jk707xYzg211hIkVTQmcmy
KOWavF4JLof2omW/e+NtZW13/FUka9UezWkRn1tUidFS65c6GJfy0YeJ7clMWllfo4oclzthUzP7
99FMbD4BHQiGqlTaas4I/pWuMB1vXzdROv1Tt5THmAAMnGVYM1O11TeN1CPi/NlHge4hAjSvtFtx
B96qfHND080LTuHl5x/exYKthaTUR29QrfXhEA0H4Qlfrj6C6tcpXfYlncMTJbrk4PFBHSQ/pi2m
gsm0eHjNHGd0/YZd1NOYFiIDg9o8K/0vLFdA6zGWGBsJquvMt9Erl5HI/VVYcbJN1wI74TlwQ40v
M8J3EFHwAii7JYyrLNYX5EsF4BRHu59Du+bxI1L5NwOksUho6V4RzLI/dgiXW2FKFYuw+Ady4Zo7
ja54fB4cSTlk61FyMYD81lrjil5DGu/JHm0ioVfsySIsQSVAN4rfqB2vwi6u/suX6UeoCUECfo4P
/h+mHmLx2M5JAIYeUhg6OsRQ6WeogCQvoRTSpzaeZO6qpego+p4CTuXL5XMnQNRiG8BkSfp2EAeD
dFBGTUATbW4oa2vIkDpSbVHYfWki+43SScSRnbsrhi1nMhOX43UryOg2s8imI4+nslPw92aiaOqK
9nTCETja7N3upCov3Tb+Z5VLvcAG3VyPvh2L6X2PfRHSbH6IoOJK27yvbkW5WtA8xddaflGWgsaP
miyxN/4mdmOP6b2vwzdjCf8FF+v+vZZrLeSPpfMcpDpOe1YURqGkIJZ/qCU9zhvNEj0IwviGKPw1
knn1+dkTTsckXyri26oF0lBPzKyteZmyPEhEBBaI3fNDt79L5Pf7qg32Nr5wononKTTuKRGTI7yQ
5m6wRch8tA2OlOZAUiMSfZuUssMD3R6dI9YpFTTK2r5xYvJMbiHcS5jkJozp2giJ2bSFx7grZhAH
vFl/s3+0/f2wkx6rCcQHlO6sGLhAuyIz7RdCtlFAKm5r6wVfcnIBbZ0OG0qeceqTtRSqWVJta004
VXffnniDaC9MuuYCC76CGNzcqzRjsaAHm0bx2Y1+Vcn3p4TmZ6EsHOHnMfVbJSogMPKhWizSoRz9
x8i32KS0c7CX+pB0D7dXUFnCqLPu7yXZSXgnSHQcsoHGvojNW7RMlD0s0bBb/n0WOgp+E/DfmDbz
iKoL4u4UAFtvlpEixGIzQ7qHV8ktxIrSwVXSEu6mWghOZXu8XOWc86GnhIGU+2fTD1g3CxnA/zrk
iUTFU8DrQqOpBlzl6u0fPS/aqrL9ri+H5qz7+YesqSY0/4Gv8NDnYAA5U5YsFzqQh7NvcRUaVTHc
//byA679mWRL8xzIR1IQdzlFfebMUBg1TeMCUQlRpLC7NZp1uic+rEA7QBL570ZKZjroXWDzEisk
Yv2cCNXb4RazAsXBWZCLvE6l/0ogJA/Xv7wLRPz57ukb8wRuXD1AAHkPpWi2WuvhXDYCaddJJY58
Ut6JW6tEHmPqA7TloM3k6RS3bBLckJ6iBhSCr+JW+MJ2EBtz8UR/qio2uEmLv3F3b25Ma1DpEgFO
2KLy/7jakExpx8ykWLkT4SoTbg+oFds6E4DldmV1qA2hWen51dQ+SUpEhPAYjyaieLbKR8/9j6CQ
kjCuhOOHejH/CO/iQvDAeoem/CI0JdOgGNKgzketaHz6REhyqWmdafSef7s0lJD2A1Q99zK75pXE
o9YewN3aTMdarZuExBDUTSTKrZqa8eJDBgCW5OjZCbRsVsgDRG6BOghCz7XuUNZXofUsYaVyyvGf
nBZyrSwqXg0nyQBy5UXkFc8Eowa2r3pxzS06L2AKS+VQpCKdw/YXa9nwI1UZIzG+hEEd89tPOpxS
RNgpqcyXWoQf1w0pEXccyYhyStDgwMwN3xUYm5A30nHmA+NiHJv8dfVyeroJRCvnAAaUoZfxlnot
BPRvfpaavGUDJLsZMZBJCpL8pPKAVYA4O1/Hd6bUz5rIPZYTFmNUHFFHOFptDX1iejoAauiwvFfp
kebO3ljgzSBBEO/ZkRU4kSvYR7CU3q12LMsHX9C9hylXhxlvh+L1brdg17CtfD7li++DD/IqReDs
HHYIaG1rHwlUaIz5dp5+p062VLKeTJME8podQr1Y/zjt9n5594f8W/dFPIHM3QFTtN/qZObPGme5
zkhsoPR3z0Zp2vffENUqkE2k/Qui6XU3VAGGRa2jkiD7+3vHTU2BozpYP5ZGnZ5W1tuOnigCoxMn
hH9zg2q6NCS4s+Ts9y+eELsYu8arnwuXHoaXiip3nqKIUXKRvYH/c9ea5SAtNFuKX4BOJQMt/tBw
rIiZGkOYe0gQtaoxsfod5S4bTSp4cYzoHZWfR7daneKvAcXGIK6w4ClFxWgU4/T89FgrPNncKXwu
9wJ1yTfEGvmFguAj2ZB4wRjfl5GAn4uRjmL7fp0eITs7wdo1PPXshquwWSOIM5AorznaYIt2PVut
6UCzG/I4rxpJ2Mv/w1wa3nl9ILY+gfmbZlOg3T/sQeyC05U5bxojdzAtFDj7iYTOSYK0TtWg2w58
kgq3Kapy+m1aQWmdUb3HG92lQEOfRHqxs72i5iKigmnGArdJKKpz2wW7J4qf9qatKzFV6bGfrzcA
HExb4QIryX5qqK/M0alLyqHC15pAR2oYeKZKIS4G38hs3USC20fLMTpcyynPHgIVFmZDyICks0GV
KU4J5uZtOlFJnGr44Zd4AGeQDSmHy3HWEWm28VxckhRvXrLqXOFYHR9SOif680LOyXk8TmuQR5HU
Brt94fzJNKYg13/etO+cIG02vOh6EctRpUk1DDQ0lBuB15U12YNib3bP2pUu7Y9XRVC4D8DyMigd
n+VGUhky8Yb7mWa2ulCt5jxmDr4geDZkjtdqH12l0rCoYoMx+DNLBzR0uniJQ5RCksCwLs3n7i2c
yEu/xmggKNgQD36AejlcoxNc9KHGd/5Juzgu6QZso16GJiY32ESVKafsakxngFwq1DFzgcpD117T
bganybi7J7FhrKejMZEhRUN0VfjM9EXGxHBqC86JV9e1D8vYN3OaBnNudMXpuEZQkN0WVgEmkoj3
FGxGSJaSYY/SljI+Z3Or2ZLrJCToPZQmez6r6zV210SPhn7dJ7KCpT+9P6aBighAmFOqz9RWb0os
R3PA6ZwdNl79SNOdnEBEwQCgtFxXx/1awb0+CwLhDInUwdKYPmiv/OwWIrIiuptpG9Qjo9WocQmw
d+pLDvDxnuo7cH0L6xFXNnD9BQY0aYBR4QJe5qityfL6ZQ2swvh5i9hcPENFbALRuOwaomm464Yi
XYGYxU4aTrJAckDtP2dSyRnWv7Ecj7xpKP1QSxZWhI7tNCOmv62V1uaCXnFHOlTaE/q8jl8Zhznw
Bme6FKPolnmG/5xJINJQO9v8Z28lIjE+B2fsFbEWrrNqHFsbJMz50SDSrNSeFtY1PUSyfZQBIZCS
/Mu4DE1z5GjihR8RZtCytVCNdNCqwaJ0+wtBPgIsMHpxN/D3+EcYKI7qUirN4Uf6tInM0JIY2G82
1yqnKhe8CMRnBQ7TM3TpJM5KCX1Zz9P/YmKXkbJNyW6F6g4JhODlGdsRD8OXlI08N3xgJpB0D/x2
Pq7E4+qjpPNGHBRBj8lyVhesY2+QIlFFu5c4hD0iRfuKo5Q8FI9shlOxdvarHIFNs+yv9EPw9nA1
qUS3y7ybwd6WNSZ31KJZiseE1EMhCxzGobs5Bq3Z+4n2jdnzi3wJt6J/QYJg9CPnyT+L7/9IjpuJ
O8KrdX4eYgRytyygqRuX0t7y2yhmzXcfFilTXfNM6VZbLI9q4IZnnPMu2LmhLPkohqBx8gsUOaLy
+jJt13qtCH7shNA3jFyKxOahszCVp0bR5nnk5952rxzu9m7WtuVgWWkQmNkPHYCYguYEiUlE2qPU
niEMlIKRU6/+rCSj0jX6/BEzt7uM6V5IjOF+Q2JP2dRUp77lTg6b4yY3XNDWGWosb1UL4F6K36hf
FspQxXg/99EZw/ynxh8+C+TjnpNprLZf9jDR6ajvJxApWw3AiIs8YxlRKc9MzksDsq3s22/9LFxU
DIIpZHE+a03PHFUJwogtTLhpyWDUzkKxv3+TXUlYDQ+xY6BY2h/2vgIxSXKGghgoFsl5VVbEjSmM
xHgcBWX1sGjVrnhfdxIy0M5vOUiZiiAsPzg68zwi42qu75AY14zAoJuMNPZqXX4jbu7ppkXyrA/x
LveiIGUEWeqOtO8wRq5A24dpBSLuNx6ykPK1kTRZgsMeIugd73rDsCiU2wdupz62z/JBLS6ZKJO/
iheulBZG0w5eR9eE2my3RX2F2SFAIsBf8GMUK4IMBqtAoA1eDBH4lORrEx+7pebG5VcnkmmY7l0k
4MSST7tq77Q2gHTMB/JhLU6g+PX0j9fUT7/Gn4dM6Zk6i1+6k9lOUs79o0++cQKC81pgooQmOq4y
qwM/ENAx8nNncOOhAsYI129gDjZjKL0gU+uNk/hcGi5yPTDiayOUTj6whXxUFlAGYkc9FcQLh6+O
5zC/E0jO60n5vLCXN4wf5z5sH97/kQypWmyCfIC/SA8IB2nSSAq+8Zo8xBEjmGI4Qrf1cvpgO68b
dt773gL3/gcgLjgszxih6M7gPjVjaleWcMdNRgmNFn5YZJVzdocCIqs/sInl5Tutjqp1rSIGUOyW
tktqa/QSs89sKa7hOThD2sz+frbxluf5DOzZ+OsY+GS3n10SwqZHCA17D0x8GPa5QYBF9KmOUiAM
DgjDfE5pwSWgT/FXctsKveVPoOEcUYmKHKeVZTZ3wW9bNuR5x2Hnn8JzzGL7jLNba8HhMaqC8ZzM
LU9Xkjk7cPPR16rqi74NPeqqDrlga28E75Oz1unRwDepD2zyd6Y6dQQUxUq55S8Fhe0R5dMThLvY
bTPXRSktVYunxs+lVSHvKQTv5adxMSyFm+XVBS7cOM9ZDD5N7eVlYqxphvFAooyjKLA2h2dChy+w
/9ZA+ITKabo6Cv9MrNFXzsoMd4fwAymIjSF4GWt1gVYwpz+1RPTh8Qgv7gmBPBmUzO/Id7A41I4e
qA4vYmG1rlpKu+MGpnCN4QMqMN2u0nhpL1+vuLSRbKkt2OQo+w6mG0S/hQ9CKpITDkKd9g/WfX61
eilcFxAmLGltIKsgOt2YaCHIQIgE5ifhkJEXGJg7RaVMcR8b9w4j26nSzVx35mr6bbcBdWtLLFj/
ieKyqXVOxmv8jE9R9nQ46YU5o//9qEXOMb1EorbOIwveN5bjvSIWs8SN8cQZ4J3LdiGUik/oAjwH
43iSRJGCGSq894fC+sagku0aQTCp2emjbPQOv+06T2eAwuWBYDg2KlTi4Lmfqv6c9JElmO6ymiCk
/5le91TrXZ8zjLlqrNj/eZfEkKUQLBVZeiCrzC0OhA/GD9dB++LTZFE4Go7rQmWBqW1umQcWvdD3
jFvBmcGduXzWG3sZucVrE8HbtSMNb1cwa2Aoz7qNu7A7CZCjofoKwGZuKcbAVex4xNX0l33dYZ9b
Z5jJetobcBVdU4uBVwSuK5AHQwW0AErjMamCKxGNI98tpT/EqmB8XfIu8V85753Fi8ifJG3KzRAL
vT7H1wqAkmRjcqxlCwE6Ak13VYAJrW9zN3OmoWPmlAUdR6TC4i5NGP3ukjengotxIjdghsBkR9XK
ZzPRBYI27fjYhGzaNGQIKS3+J9E99BppU9Ct45p7ucAcbUV4X59CARFStjvr7vQjdVeqP1950EK1
jme+6l6TowZDT4o3Pzw18XeVMVzIyYj6OJThLPUAaOmSwOZglSp8FusccjVBUcR9JiV6zdjWl532
6J86Wi8ZtrO9daRzZK4czrvtrf9TkTaoz2We+H6QOeMCZJqpdkSk8R0gH4L10k0xGJB/M4LTvZs6
7lMPzwi6pn748oDzW76SMdW6dunpl45eON0zURWH2VnRoP53n9S1E6vkBG4TROt2fc55pKUIDiQX
qEcXeIw4mHXO91qgA4H7q97/ai0P+AFYHstCkropwmL6qZ3AUhqchHJJS+Gj5OIcl2fhSfkuZ44J
s+IUY51O1KeFyMUFX37LDLzuU/X8hhiDaQpd6NA7El7jBFVsefCkQotB3bJqoiRx23toF8CIaKOB
1JXbwDT9Z78HrPZmZVSj/OYW804YLpbVJqLkGw3cgrs6GW+CLWfpBtNvdmwVjB1wGTZqEn0LAw2e
d6sYnNnvRk7iOBRrWTwiP5aJ7be5LNdZxcpdgfVbcQuWxV9BvbW2cqPompY4OUlSNN5uh9FbNc49
QNygkvp/Up8ugIMDrXUeadXvggI5ywUqr4BF7b5TMptnvC44crv9Q9DvUmXKByGijBcgnOF32tE/
+uPBmo4yj8Y4JbwpWBmLpeBAnDOpJxLqs3RDw0G7sVT79mLpnfx64OgGWZJqVZYsEo247Bzlqa/o
k55jQgR1cuR5saOq96UshoZTReT4+bF3lUztyMUejBkC4CGpjY4iJQbYl7wJ7LpZdHT8xf4j1Dgm
O9xckOpADXYB2DZO936k10Ed7cz0o7F9G3OLbA+B1ADeltw6Z9LDu1J0Cpn9XnDw/pC2dQEo0FtL
udrncHrFklqEMoY8jCVpBA+viFv5jAY/6wCw0WxvRWIuLblE4zr2AOSsQnsz2303w6JvaAHkLR3z
RVPD72kGgkS3bdq23xxDyzYfBKdmuFBX57RhltmaKLH+PTYVraSO8aSv/7uaA5qDtRnAWBCo4KXx
Pm1IpkDf5WaT+JFvW/DLJVgV9WQciaueCSoN8Oypkpks76lOseyG7AclC6nslbdfkMfVt5DVbb29
xxXvO3iTHc7IqXCL7MAhM7YLmZ50KOdWNf9xyVj8sEtlkS9MjgA65QKWFfBcURSTUNno7HdoVJh5
0lCAXR6MPYJROa9JijgXeX2TWYoGECWbtxrTxQlDOSpWK4gAYXtvVq9pu+QyrXgFodams6ZE9F+e
vO5cfFPrQGoBn7K7t+RH7WHmsn3s3XFq6IrqQJubZ1nKrIXdc7cLfyzI7Vy9mKqsNN6UP6J6l55Z
cP/EBvdF5TH0sl/vZswJ8pzTcc7VBpGV6KLNuQLAZMKSVNX2P+kFhDnW2HnVkG8guoeAhpHFzATu
vqsF3tXuDsQcrlxOPzF9HrxxOO2eb9a4nclleFcI2li2/T8EvhutU6UejC+lz/XkO8GysPRFEQHf
NGYznQEf9JblVvEezP8H5fo2yoH9kmYNbNVj3Fm/74w+l8K4W/2GvSafzDjQ1MK46rriR5LLW73z
nBQu+zWDXuVRFheaOvAiJUw3nnYh24LjxF/XCM+RlD7CssmvBCzK9wgHRVvB99pLWjGgS/NU6YC3
tzyVETKKhdzSBFVVycQHyxAJbpPwA/ETA0yjXKyAvScCAnBEU5a/EqbUwmys0+Vz2lSySvx+dLDO
OiopvYZABpbII8xSmOyA6mN8EdHjMZenDDtAZcZeBJ5Ilk+6Q7BC49fuDUhVWUn2ya95lKMSbmc9
PdS73YIpuoID6dDaEjfw5gkXwKh+BdY43wrGUcZMb/AKAsbEqX0BebG+c2dRRZ/ck0jy8zRIGIaG
gsUfzQk0YPFuhrQHbQbFmaw12Bw9kHzAStF3GGepWHBksKuKDwKkTE35bzWS8my0i2B6flqQg8WW
kZBDp1EdZAYhBY964s8+648XPB+Qbz3avH+SuiTl3eShhHkF4rNZYcRfPy5//JPvQaihTLaRVuNM
DxxnqiJwyHIGgYjnkCu6H9YBf36Kx+9yg2JmIqrS4KlrFNzSb9bug4GXhdmU5qmTu3DlNXgZqht0
3h9wfKEaohgQM34my/STea9o7lBZx4jIFrTo0qp1q6e92k2mjqc82qghvonrLnhL+ai1sba8zfwW
oyHzEHwIl+PYWNOpOBZExKadwB4x96lXAXATBZwkLwQqLXLovQvAx0L+hwmyZKF4WcHr1UPw/YS0
TcIlFx7iNJMy9Sa18g/iKIbmSVLYkRSrKVSjdMVkILJaJ1JzzeDZXmR3RbVVK4s2rCzk4JqCCB8T
3ZXiq5Wmtx4NYSBncelnXCfd7Lqy1wTeW91pYkaFSGOVLOL3io8GuG7N9ns1F4vb6atMzSfZNP/4
NNojKF+yVQxFI9nQSxdUywp2C01TTGzg5F5L8+sYFXzWvHuOK0OeozsFXzZQ9YKAr1cBCZkY7Gi6
gLLhJlfrZqIvoPBtUnu8xrghF1oknny8wO6lGjhKj4+WwGLdTvM+TLlVZvQ+IbZtf/ItKdTj3A9w
reikk+eUdNzcGnOUHDjtX6sEKnFzqewcrQkjTF4zfnE/dExdo1YyUUVCw33LYpXtRthabf4bcYyx
YKJQNNDok/07PMmwhP1XBGZi7qIF7KOZbvZQYFBJaWys4+PCWSfZ4bTrpb7Pi0AnyIvtrGaIu+Rc
DPSMdUtOyOxerlZ3xjOLQGPm4uFJfAIpSTfvSqol5snknmb+Is3JYS1KQhyezOimf+68x1GqYUF1
qKyftx7eqVqRb62KBDQRWvLeTbT8NkUOtRUy/94BZxYv7rXVI8AtQc8FtzvRiADitSFmX2725Jzi
rw/7u2WeQG1OiuOdylT5cpi7dbONN/ENg68aSqADwXO+zl3+6hedXJNcfjYWW4tq7a3+iIDkfWtq
2sG2vCoE5LPByl4qZXS3Zbeq/ntlS61gDaJJ2VI/FNiwSBLRqekJcf9MzQKOGBalFSk6XhG4+9zj
BdylT5SAR1WH8LBd9Ps1jZb3SjkYUcR/sEQhy6GHvFuoA4I2fKi540G0b3ljuQU/FcHp0epBuvgU
uN7XjrFzbqi4/okU1rf6g7w6DTQmckOJNUa+0pgrLxY0l7Z85s6n/di6hSpYqhdyJvucPZGkIHPT
fnr9lD9012E1LemBWy0JRUWcNQzH2sStoJPInQwsS18dABC5GYF56p0d0X8VueHgZsrtFnCzpwse
tCQ/6GfOqYFud4zqSBaybzvp0hX4Ki4uIOoKoOn0f57zA7Yu703l9Zqxp+1mEztumdYJauw4v3vk
3SGE2vaPfo7YoUEUXvPI3z1RGYJjdJ33Vi0YHJRFxaiLZ/17khSwzQVzU4gAeOO/5bJWf7At8ho7
v8gSkcPUyDiRz65YZdKko0zhP1GeDARFSXoXu5jrGthrOUf8qgwYSHjLOdWv/H2hGFZHiqVs8Dx8
fHGXEn4vfXp0IUJZzYXwVN9G9O+plECt8G2xYwl60ScAwdZkTKEM+5QTQj0WfFsDPc9JfSuUrQkR
NucdHvXbD2LanOdel7jxQGDqDDkQ4/AKgYhJBUHgg0GWzaAbm8kKbGfOwxgmvB1Dc3LAuC3JyGGm
ODjKYwQY7jTncS/L0yFDbVs45b3g4z0Ps4rme4JQ/C27sk97xdnv832CoaB7M4Tn1uJH8I1VB2o/
9jCkUypnYmHCmOmgA8hHeD0Noo8VOxo87FTkOMQpsU+bT8NYCkQ6XreJiY4eYfi39I1+IpQJ6/d5
kg9f6gr8tVZywK+xFxLTMJm/2jPOaDdYn8/CD6sntOBVzGs5BPcNv4mwLhx7JrmVPEwOoJDRkWeC
QRxwzqIC8oN2g4Ew1EC/uLLC6YuPu3YDFJBbn3iwcdq/TrtxninvnOf+3CVkTmDkIs+DQhVnd+Xg
Og34I0VYn7ED4SgsST4WXNZ6YbmS/bQ01rit/WobEfRM1apFUxF8iKI22OqKTryAgnMTCHrHUwp7
nMIq62V9R6tcwhj8JPThcaIClAdvLkbizWIYZ0CCj7p+A5x3B28sOdR0iE3IkikiyiN61BTI1xlA
Kfv/86grVCs0CKv795NXqBImaAq7tu5w48Iutm1XDorNuzhyFUgy44wGrwkvX3qQB/lBskVJeoxx
NDTBxGZFYZifpMwekI7V1dgqa5XX5LrbIOb/xruyxoflDTWVPDD+KhfBtPTsKDTLYD+PKf61hndI
Ku36JjMFLWFOswdT5WfFvOhxmgH3Elw9ziriL5c+GXroVkDpxbtrYMPLOZPNpVr7AR5Rw8tOXnzk
P3yPsqmlpHrv9dNB5xXMP+LhbHz6JCljDuZsag1i5x/1tiqj5WwP44x65SVzUXoqwiRUzgOtoGPl
EkfxzM6BGsk2QNSWIse+hygs4G7zodWqlodR8X4Ua3ye4SUn2cRTsjNMAQbCpm0l4QbBWwPER8Os
XL74e67CYZMFyEYMZBj3IN+VltEop1+cEo7WbtaIJ72tJmotylyuwU6IrZJr3UwZ1+TmZ4kmD7xl
u1hF594JnroOzzzHqlodmYwuTULdXh4uGNpV4TDfb2gjzePnHcqD97k76qjB0BUC4MezAelIQE7N
vjojLWtQoeMB/tj8H3ITges1IJ5+hi+nsrk4xr1JlgM57tDwAXivItjng8ZwMAPqZG2LSGjMVTGd
ZUxLmaqr2G5o0ZrkqznQZcvCT6un45dmFbS9dUAEk+g4f4u/VSw0uKevWSS35ITOd8ePvbnHMxMY
NiYolQTYxQfJKTvsxupaOgIowkNSSYKKCevXtWdIsOPZV6f3jOudtHe+09J44f0sArfc2X2JRs2w
bs3+fwPaoF1osQd8SuCFL1vYBtCzQLYyaFGo++4+KTNjryt4UpKgAS31AQksBnU7TAVeFYqcoqpW
J3clPXRYCIzkymrSjh7x5+TVqd5/Q5JxzzGYeWxpZpodygnJaSVr4pkMEUloevPizGrhK1sOfTtH
w0JyWVbGbENFZF+h0KIkOWH7d0RLKeWf9sSaI5gJnuExhviUrrvdURS/yDpGYS0lPCrprAqclG6f
EL+6G2y8+B2xSJsFdpSk4lkHA4l9f/vCWnYmx+htS049D0RT3JuijPnni2vIZf59B2EzEzSUGKkk
EhtPOr7gYPSkknbIu7FWS/2j6FG4YtR0MrOBDIntpZEMCOGzbd/TxEixkluu/40nuoy6i6oZ/PQV
AiPlkiFbtQLGoSiHeCkPgdY3P6yfmFUvKKOcWJQj1HkMVejs08ajBn6mxMHUG9HQwy7hmvez26VQ
KKrn6A4HfrxKST1u7ZlbFJCDq2C/eCfMmdcdbLdbYjWAAWr8GTUjCU/KZorHDkRvo0iMxLhRh+p1
3Ei5r5Ce9bafIJRKGFtdXIglkxx5LzO7Ai1LwrhRZVoBxriizCZ5cCYtJy/iqfKecsll1PYYKeGM
70iUWBcyhpIGkipClnZEqXqK1YFPz62OwJOccEb69U5NuLTUkzyUMZqDnklNBIE81eVazimimRdP
NinAOS7/dcNlA8UWcKNPjuAZPF67IkpOJk7UZTBGyhImqY3sZ077A5D5fOLDTQwx/6rwuS/uisaB
CdZD2OrKlNTOgbdIoq/2jca9JU8qob6QKvIelQwwCDnIajfC3uKyB30K35ujCtIUctc6xazJoV0c
qJk2K1Y/UhHcNAao4kEfammA/JwqLLIS9FP9am8fVPFbnvQTqjpEDd6ERjKJQwIYZi6/imqGuLuS
OFEa/KTvqVZpFEP5L4T9FHAmV3Xs1PmK0t0UmirduBAc5xzaICHqxaU+qXW6JtLPbxZcUyGA2fAA
YyGnCVNFkFzTRB75hSVhnXVjLp8PwI37/GqqmDqQHgSf2Gc2IF8fjgdC7FlUpnJlSrIdGvGBdB2K
50zhG7XiDhgETOOjvDJRtalKI0X9kZNnPJyaYgweqZ3w4hTuWyGZByp3t3J1luMDad30IzkO6Cck
OUMtWVkQjlGLwCvmj08v3scnmscDx2ctPekZTBaEOS/K5ZYYR3ayCW5bAN+37y49xfxbOvmL6T0u
4ysPPTRgRQim2wqCCAn8ST25ZAxSwqkN/L3SSlguPn1AgxMEH9AKIQeo98N9ndHXd5D9y9fEgn9s
YWisSD1h8eNmeo6t442RNF5j0IZpTrO5Z9u8jcPah8LctaBTPuEOj4bOcanWPMDDI276lJX5jZwI
zxRyb1s+B/JxVq+iAMgw3XFiIaQLrmzVDlRqLHFGYCcJjonKQhwtez5XJm47ze2DxoXevq8o1Zra
nB+ukM3Xo6IibTSdnUSZrBm511Kv2z3/AjRAWiG6RCFtz6WwprU5mY5CdL4riYyzbdHojrHAARNv
ryrRMLKMMUBXur8Us74NzUYFL6tU3CE1VbSe/YCndW97M/PHRuPfRBYqWrgo4nf7LJuF5OLS2YJL
3Ufnlq1b2VF4oVGryClWclJEnxeBdq6+Q6brdgeIc4+rw58lxf9tGrlOq+sM95GBmj8Zljsi7w3+
lkw1RdSa1e+/Q0vcGW+eyMYIAQCSI9p+9bu2Fzvg34SLYoZf5ooaZujwl2nzRR39zi84G5SW7jqi
XadOxtR/Xoe+xf0EmammHqqYpGOSJ/OxLHkjsN1VEnfkVDSJgV1VzP36a+c8iug6vEn/xAHmdOrn
8Naer8DHfxlZgRilOmT4BDKSdOmtde7iNOjlqQ11A+BRqKCt6beKcfkIdkMSd1IYA0uLCunduzyC
2kv6SnNaV70iPaYnS0ifpcp86YRdUSpv9KV+0GbRMhVT0wFg0l4ozQvAGP+FZT9KnIWnUb29OeeZ
JwnM41QSVsVYTGx7sMCvIvPZJgvJZhlUUpZ0FYxlINDr1FAbq6MqsNE9d8gluZP3uMrPjv1TDNEf
QCR2D/VyhmrKl2o7N25/gzbldEoiYQrCU3W0PDtOlkPYYtf4dqg794HjLZgZwhkHdnQYiDDrSG4Y
/19/OC1vMPXptkx/PSYynVog1TbW2byy0gMMNre9CRIL0mRr7rIdlsL3X+TWO1mnlinCgPWm1Zld
lMWVsLGjN49+wgmLK1NP60i48Bz67k1pSHJ9PntUULmZqXht0hjlyTHfKDY8ybI+Cf8Tn3Qz1u4Y
7T/XBBG5rTNOe/RMj+uacYxkB9namuU9UxSAE8x1r1RvTkq3G9WjxynXYpx/F2sYj0Njpb34jwE+
cbAitHrmPNtU54M0hf5DoAihW8kqLeJ5zUrJ0bY7hWUcXr24v3jaYVozEM/6uEFCKsBc8bt/C3Np
pH7VUq5AaqYb8WSmf73Qurft2Gdow9LSX988eQ7ra5CmbbCUEabvPmXgDRcq2BfhbUfwwOkPrfw5
8eu74Ij1COZzdEBu+41QwYY5qV0R2HPd96Mf5akp+oyqlNpxMALLiIo8Z0zlk4pCsbw8EXuNqxE1
tRLIZUlx5VFI1839B64C/8wC5YCvwwQ8It/pr3lsylbJuPc+48c7JT67tkLrsx0/smBNwTYwSZLC
/zDZ5LBFu/wLpaDFHccHHTOTlZG1sFqAuaohFd5Jid3s1bvkZrhg3d1ohJ6jAmnjzPZFEVNms/O7
JxmhFcTTwTZfxK7lstPtTUcMbrVLMROUfl8OXrW9CR6BifXWBJUR3hnJx8KExxAWUtTGzoeotBpC
hymVfOuL/gJavdqL7/UX1AwudT07D4AZKdxGS+UZQKyMndWga4DaWqZ2vSw60hlzBe1d2hLolGRb
z5kouwMjzlwofxf25xXW/+cWsQ+vbeTI+wCPJUr+6vaqd2W6IMn8PhtQZ14AAYmnA8XF1+qaDzMr
DWAzR0d3ISUEZAlfH+7yOZVhYnGSGHcRluszyBqJG39Myotz5Rt2fC1V/DeBoVRoPcihjBjwz086
YSrkv6Et9q+Z8VoFS0My/N8sJydmD5d9NLWkUIvCIGTjZd+dq2WYt7j93z0/7l2QypLgSJFIYmX7
IhUmVrfmOQ9GWDl9i8767G68rFhi4wkKwWLv52pD0ITTK2JQ0iP4Ps6vHFNc9ru354sLTvaftJiY
ZGup12tLjYs5l7i+gy/VLpb3AJlgCDsDdFXxtKMV8yj8VmRIIno+8jiakp7WeYpDisei/H+qAeNx
0CYOuqyB8NHEyeXB0ctTjq1ww/GmwHWZ8f9Xplf93bnjsQZJF/2ffM50kBKQR+ZZHaXzrFzxKHvk
WPZq5ZDS3FrrxbByQ2D7y6zm0H/nlDDRAUsGVbSuuOmRS5mAXGbkSUj1j9nust5h9ZiAgdL3OIPP
EDaXwfNdijQl6Fl1hiEFIgZCsiNoqzddvqUJjElmyzM/Ra1IG4sKmW2WXNuQDrrUaoA5ezMSJA1V
zKqTAtGVHAJKr0ze1LFqKp9HDbjt+cu6kS+itWK9prtJ5gGkRsQkhz9ggzhmpcu1tL/kwrppiSB5
cyr/bW47gUCvcLlB336+LUcrHekU4Bh36q6nWPIc4pmNERRZptV8FSzts8j2JYfg2ndOQHqg2+V0
Slo9YAL3+93oSQtfx3cSh1swYwBSckyDO7s2lJ8n/43EJLW4rpG/Osvx1eA7j+g7kDKfq56vSAVP
EIX7sLuxKgvQTPkh41UaAOCVtr7x7BwtSotqMDI6Fvc+ZeCEyPX/wMZSu4QxNKdaLikxafXPsj5e
qYeT55sclKUqzpH4ESQIhbE1B7hwlwDJSZDpSRwAk5lS+tp33l1LljgLvSjc8qB53b76CTWh/nuW
79ZRGXuXuu7TF30Z/ykwkIOEulaJNVC/aJtA+W+nmrUw8xsz9QMIDSx/Wzp87H9qCWeGHuLhTuSA
jLxU+Ykg4r5oDCD4VxCMMwy2/UKiOtmJyZOO+drcMYRFFl3TLSmsOmIJLcfRQVR+mUkFu2ym2YgM
srVgzKIJV9/mzMvTFk/UncP/p35upY3MBsW+kaAjHKPdbSrPlyLQUw/lq4OKmZpxk1zJU9ywLtZ9
ID/ZXgRTJ/PsLGpEVBHGfATPkL2Rfd0NcOcY72rN/iQJy0m8JYxdHxeFxHzWjWcHTUFisCvbeR+v
e1UhNsSifj3/SV9S25pfGjX3UyB9QdW1QFZYlUkpG8vIx1WGaQiU00BVduX7D2Wosoc/WM4ns1QO
tmi8zesfVFxmhK13YCk5z5W6H7Mhbz7LbwCiFLpfsOoCGXzJsWsML3cTqP+1LRyT+pwanjIQ/dCg
lvlQNgQRToMRLoa+w9aCvWt7N4BLExgbzb1wlC3/7MsyiiqPKlbLZ2xo78BruhVMsD/9snSx5bVF
bYc4zZA8V0bqBnxX+Rul9v5zR7wmWwPk/CF1MbIWk5k/L8HR0g5BBowMDYuZ6IINg4a8wMiHIXI2
MVTNUbGvXDQoWBACF9c9+2kFVFlYOT5CtTwhnBQiOUz5MpfdpTBvhQLMU0hS6Zn9oIa00gDtwbqp
9pUkNcDbcK0orv/8GAqnP6HfAXfxuOPY2EObhzXEuh67U5Lkuum545CB4QkZjgum6cuBRIZER/tJ
Y+rlbmeATLz1VlMOPcA6fro8xg/2hhUFh+pVQo4OTCiwKroq8NIpZz9KhdaDzcJYg6rQfZLijeHr
zBjrC+SP6jVAqN2qbl0RUyzmh8k6DXtwhft4ZrbGmo5M8r+0B+6wfNh0EyRFzYsn+zIDr3QJFZvq
rq/OJDmI7ySFYsZ3tAXechsNKft1pbLJBk/3FhHG/8XR1YpK1caO5SkRNRTaIymjWI42VfqVOezg
/PbRJxkLTZsFqE9sENE+3SXG21shODj/lKQH+cz17FbsIPQF6HQmJLIM/U+JKej19P2qkefrjYOm
pWwryBfN4iaAjdkfUqqxRuJCMi3oP89wxu5dxzrI+H7cZPCalCtFMWjal0wjO+gSZuWvia64jX1L
rKQ2YJI3a1s8ADEW2Xbhnrb+qrsbUf/KzzWWRyrqLD39XqYpJWZGggPmJYhsNlpmPA4mP7Bazasj
LhWk0pNJDDCRyYLmIVtIH94xACkao/f7de92g5oA9PcNfVXt1701Q7I+Rseq/YPt3bRgkP/2XAjt
JAZFD0ZYlZDHNlRWNLgd1LmMWCKJ0siIE/EHvJ+Rhv10G8FxA6tdhvo7eA/qMk0lM/K3k2ir7XS3
jxKSHEGK1dHVnE7E/T4PAvCUeOxZpypTOXm2Gon0g9yo07XvDsY/Wt5bE2oKVkNjP07Qan/7gTe0
hBrNynuMyd/0tb/zkB52t5aiP2fvMznvnylW/adVTEXOIrscR06bhxsakxmBXpoj/aMzwcVY9ECI
D71Z6CRLU3V5cKEUzNBN4DnPvOOkvlqfQHiFNBCTbFSLoeYOE8mehkbTwMHRyXXyvdfG9MaBw+Tk
Z8rKUhr2kCLHacTshZhfnU9n5FafhwEEqy2505gjqn3oAZIfDJF04+zdw/WlqIoni+Xj0LLf5EfQ
ZLhAeVXbvhKgvNhwwDLFw7c4N24EQ51MtPmpFr+/p6VPBADpCpI/6hM84zIfy4L8WvAn4Yhrw0xS
/RPe5S1YXfJtGpf+gqsFMLq9+csY/Q4nsypLLsqKilno3aWXHECudNPoDsXkDtxvTwdSK4HWT4VF
Pf2vv/cUOXv/y673+KXflcEt6oJJrkgecBc4poMGe+bF6EZyIujBRPggPNSk+tPSWvnChrAfv750
TCRUdcB57EoexcCfrUfTwUXZPvwMKjDLtLXVjBfCzG6F4NoYEup2kZFCYJH1u7dvN8KaijJP29pB
az1N8QirUauT6plVbRac2W/qp5oOCyaDg6Zjk1fraPyEriwsyrY428GROdJM/dp64CcxVoyueTrJ
nWANHnOVIY1Efpm3mFCvUbuKeOlOkiBu/NQDtCoz5Mw5f4gA8KQikDfB6fOjjKGpdBsk/3CiaxMP
3uXvwdN004ljq9YFc6oHMNLwiz9SmaJWEabZ2J+JazvJmo4XQBrfjbs5yyC19kx3XsLzUCD9mjbh
W+dUUQIfe819WshiVDmFZ+sRKOM+Oy22ZR52gxW3yvvzYL0odde65uIZBMZPK0KUhYhUryjwMbee
+guqiRAjQPpacbgaA7+OaXZOEA1PvNqWekxiCsxQ326gtacq0n9QZws9SCBMDmX4+jl8kmh09cpd
BzunJryz4konDHmKeC0jKpyVMV3/kYLVCz/x1GRK3HjeaFyNFpIGIZ/IR09yeQAK8InIx1pgv/qR
CpUr2YLUg0iN73pegyCvYlgpEV7Lq6TijEMn65FZxE9iNfE9onI31lbFLWIHgo+hobC8HmLVDiFG
KkBYUP1le5tIc9sJ0QhhxZJnNqp5fcOqBQ5t31vHhVWpppdGbPcT1Akjl446ieJnmBg/psg+FT3u
eLKlM75G3aee6LxT11aoOrOwCymUBJJe6WUql24KftY0CC3yuVfegXqcbkc+8Y42OSn7tXwZ3T1n
o9YnUNAMTU0Fk2TVkRzKoVlAOKyjw5euIo+EoZuBbrixw6Tzgq/isWnaaBpZCHHaa8OVvTnFeXiz
ZOc2zfx0Nkj48JJQb502qJdJ38q51i98e9V6/wcVZqQCOQ/Pw5pGSqiw5ejUCsjbtW3ML3gxP+zP
Hhq3EE+bVyEu2hyClv5lYnuazyncBcT90u1cdoi4zcx5Ve1UW9PvntnCrxocr7JWkgRyFmepdOvH
dqko8pB5DmA/Nszx89Qzt1NDjrztlb+zwYqI0Hrf0WuNGSRnorKPHjZhqrDAyEAfnX/SebGmuoop
WqVXUz5wBAoa1cAfFKtn0z4B99P2zIIx947bBOUW/5Epwdsu4YtvLKGSSZB+Jl0mIDk/7AGDqMCM
BCwRoZRuHRpxIGSW9yDXTXnvUYMUAlQ4Bw+aR67ay4v9hLX07uC6E9CLtVF9HEp9f+xTfeFU4Qj1
qBTKhqirsxsMhIFPlqmIunE3qm3TomLJtSaLy2+Nx3STrm/CwUui1o6HpDhmsx/8eWcBBvWg3vtV
JCkdn7vp//sLlNf/5w6jINYl5IcyS/c79iet7sKwEt+4PPB/aiASqe22ZJe2Jz30TJnjyRC+cJJu
Z54z4avlNXJBAYDjIfw90HQ3IK5VhOq2c6YU1n3sszDFuHsEh9ZNzN7HkiGGeAkr5pUjKebAWFeA
qLBJiM/Uqt5YL6CVheYTAra3w4XfjsCgFBEEUjh61Ytobpo/u2mDexwBezZprM/EjfhkVSWCfYnc
xcNtEgMT1LsU8AyVsGWIUktvNU5NNybf1rDlNV/CTYQVXTN1zsXiVHVOb7PuZh9CtAKT2sBTmZtR
qOMxoQgLe9vBse3b5xZWMCXocLNF2RgxcocnGrOj+Iuk2OifF+b3jKC4zwiIirXv6Q4RJorAps/t
NJgHr6/oT+Qroq2+D5Wxrkv7MaQ5EjRPXmL8O7b8RSQkHkwtEziHZtT1RJDXy9EVLwNYWcNRRV4F
aCVroydR3NKKf+/9/C428bJCNJOtiC7ZqsHqpTFckW/85Ubzx3WfQGFOuiMebapPEx8U+KRT7SeD
g70optfpCXyVZlFdxsK5rA3F6uDrQODSNO36T9GNs+eSdpA0OQTl4kNny+IF486FIuseI/HdOPD1
a4jOxIfW0ENvgqB1Zm7yPVYnlFYKYdUJ9Rd9ogv+zMla2IS4SlvdNmjDE1UJ90sU5RDRwuA8/3Yd
FO4yQyd02N6VXIDv4BjhXmT1kJ4QCQENQ2HcCEIlLwjZJs/9gcqs+rcnVP3xmg+fIrq6B2wn78VL
kfAAvZMUDrtZt/ATe4aQbUv3sJIyXtOilLImrdpgne/2HWuBTnVaexUe+vW+KgohGm5RcA5BWO4l
U2we9xgv0L4chrbMpqTG4NIkclS5D5EniiYNo2M6sYZj64CZI4qHv0O23MZtOEmrVegbmN5L4jFx
QTBNR3h/vVswHovZyaGaQ8Znpj7Dn6YaFkUtXoDJNg1kFX0amZFN+0edRuTHhaxGhOoPAeaHTMCH
DrzUqUdQxmP+ZoEdo7z9HzlUh8srYmMtpEjI6MPah/fCXLIjxZwQgBQzjcQyP1QPWNGsnJh7QvfN
AIbyaftnHxEHplj1wnGxzxMHsqPmuAtwVZLvBvIm5h0H/y2jMlWgi3aT+XV0OINORmAQSEc2p3S7
hfYTXcy9iOJ1kuw/SeYbZYCZUytioWf2DA14eLl2YgU8XEpInGsH96H8oHz+2NAfmwhTv552mDj/
HBC8C+qYMeV3kzS9+JEfQcX36g8RBMs0/3q79bDqT3No0wxP7tbde53uaJRwMxAp9+HUCgrhVbt5
6sLTrgtmGVRfOZgtXDi7E5/YOVGIYKUOvXAFvfOwpdLXwhb4En50GRd+/TeSJHgntImTUNPWdVPZ
pvn8N5nNcsSJV5LYVDKJFp2DcX+HQKwZE8Paa3a8e8yF+pEYHwPWRsf8KvXKAMaC0eLffo2fLkS0
BLSF7qV4d9g0SgCDBN8uxxBAau6IQ9rh9d8j8jgfpwnRdJmg1Co98bZ6PGLnIUu7BPX6B5ngLb4L
5rwKvnW4+X3e6XoY3+zK00OZhzyILK9N15Y3I7oV5wCeXMTbetHubB0qcDLkM5dKqeiUnMauzkLN
SYbDUBxD+IHmeTxtxKlpuS6ir8Icn/uaPbwqmunWHgAg6K7Ik39Kidsh/g9Xn6Pwc2E3MO67OGEy
FPGEzugcdQO9MWuymWeFcUPoF3Ia67NHr5IAzSGF0Z8trlQgUKof5xz5UgN5QurdpmybyIGCkoMX
D1mDTDsOu7bbzYu7F7w2lKVqZ2uqkTxbt5BxnOl48/ERNXPYCtjr329i9lX4NAINXpi3g6lHepzZ
9VQCPps/8Lbs80X6oE9FDELK1kGqmTapN2G8ZzDbsI9T/kLYtO0rNHA8Yy3viecYtlaYezB/I6E8
8aBGyHwiAGrTsWnvHNFqxr9jKxzQpre3beDBlAWoPf0V+mYkpgj6No33HVGtIvtIxhktehMIl+lY
QhWOjZFwIEbZSqJfF1HfaJyTGFutBRap8iZ0kMipqb7fakF7NPb/jiI7XmRnxIxIiNQi90TkQTGH
/vX6LWswGxxl6T+wC9C1Lqui1sAmF8lBNB8CPKygZgjP/h/7eSXtwSMnydzOutZzPYXc3Kgam/eZ
YE/uh40OHiwACwvLy6TYr+P15zeLLMRXXSn0SnLACNxJ9n/tiAXf87LnILEINXvcX2l/pulMEBJ+
+mDt7dQmYeniuNs61+7C17vGbbSKvfZd14/JHk64lZnQCAZevExp9Vnp/2geHuSIBYKb94sfXPY1
iV/XV8NZnl7d6tA/0gH+XBwKf/g0idL1jZVEVVuNXx3V8+klqJQ9DXu+ti+ioBPvIN7dBEV3aJmT
iIeTuHbYviBNYe2Q4cA4ZNgyyVt2EQuzKeW/uyVJgWaiXE8v/kKk6QqTWhgFVEEKEYxv1EI8dOgV
hQOzwCPpUw3mC7PqJqqBjY8pMEvFK5eprb80GCzGgtrOPGP+jow/rysfkoeXBzhwJbsTJKw09wnE
2ltv+b8vteQRvEJDkUiVfuUguS0l16QqC6I9DKpDKqWTjJK18Pw6OWosMBEUdzt0ihQrRDU3r0g9
EaH3F5Cw89+jk4uCOfqPW6J0srYjw34KNERb59/+nIg2Uaht1HP0SWpWslP+ueCVp7VoqTBgADjb
vHaMaUXjkSQKCUWn0lMUZT6GAUy4myb+Ha0BJsSknUMVKK6gBCiiXTtcRTvW4HFARX7s354ndDxO
46sC3wZVU5bzBAsUj0A2uPNLmAzCZrpaMCMI0ulBKfEg/Xgq33BQvLAr7PKe7QjeOxEk0gbnwYWc
+Hj4CxfM3/CFSaX0eK1991bcCtdEdQpjGZ5cOY9pyApMeri0Sr06PehgrWSQS1WQvwazh6F29Iyf
3NdJsMZcjmXGbPcOAjqynRz+MBqVpxVGIv4nXWbXKABOy8Q3GA16Dgo5QGfmgGcC/Eafwki4+RnL
J23BUN/vQ2QonkWCPqk2e89KojT84Z5t1Kn+sGAjAAjEc69ASk5nNdMUpLvLcVv8F7xMMwlBdsnH
VXV4WQ9e8PCzOprzmBSjt4mstYZfFv8k/+0kyuDeuWQ7eQw/C9SZBWDHssAs004BzLHzh6wGfTWH
JN8fU+CYLckc/Kw2Px1KIxvwoi3tpex1WJni2u+wShQEqQ4BeUukoHuWtKJGJ5/qcgSTLKxXuwU2
cS2gZ0C4fW12Rx4KoqZ5gQfwOSOA2fsZ1Y3WUv0rdM8CP+Vb57loaIBJtNMm9mSyHd+JdyIyQcog
jtUPz8gf6TcFJOtxZzCAuSVDekpzRtfzSUiV/okSVkaWmXsD6zIrJMRMQhXdwneR8Yei5uj19sdO
f8oADw1oYhnHeU5IYwNT+v8g6B9jZlSP+DocFo3EqpST3qYovtQFP4w8dAvCODlIcBiJnwBtLa+W
5KP4XfB9rD+Uuwm4wTQLBYxGohshpG6r+FIcSpuOnbLySgU9OaFSwfnduXtDY2PHiqp5F1co0kOm
MzRBJEsts7fxALpec/ZIZ0lN3HGQ4Hst44FyUf+iwT+vNWxqL7gphG1qXVJ9M6v3UqCRRqnNBVRd
FvSedn8RDUr8H76CUXjg3C9Mqibw/1qNXzxpuklkzF29mYJNI0UVvn2KYLMv3xQ9kLzUs9mE1c5R
4Hp2Fz9giUxcXona2G4OostLobu/IBI2AwVUDIGENJkx0xbDm3ziY90hi2QNqnAUsyRcRcSri/7V
e6ttdszfb+4AQ6WeL7PAeQKIU1I3fLneDVihdBdR97rOnlpknQx/eh8MOv2owfWtCk1GThkwOdPZ
Xq4dUHa2f/7TbJiLY9GSmJ0gGaDL4PwFBRgk3QnkE3lOTU1xs9TFmczRpQMkJPEsQ5tS27sEv4bI
4nUAJplBy6mlpXEOq+oJ3z8HTdNhTBfDZ8vq3N1vfGefi3Dw8tLo6J8oAC8ePpAmXjc6aRcloqFO
DtTVwplFOsaPjcsdyQwDqdOsn3dKnaPFnG9ThoA78RgimYjH9bjBnbmuCfMkQmkHjMABqYvO0gpx
UpxicFTJ7+tVU5jx6erkJh7f1x87gY7zHl7sNEfJh8O593Woyt8wifmMGquuYTIPDhzzj+OoxH9p
3d/yPMMmTaNGtCyPxgdSkZRihQ6N+gibqj3hUtNj2w6+/8M3LJREefjCEkh3VATA9KBjZp7HJpSV
BUpzkhwLReEceQ8NB/qLrr20jhVNN+jj4SkmaevhxyqPsYCWlxhYR/RoeW9vS0olNja7k8GpdbUt
swYU80vrxAeHTilQQp/RwPfl1FLhmNW2fTIsb9aX2HMpgkIAjmMpfOeObz5bDylE8FgbYwlsM7EU
L2KhgIJmzBAuWMn9PD4HEHnlOgyNm4B5pLC6s+yquHLhGgis+tSdfpmHqqXpsydXQ6gk7MWSq9f8
WnjkTW95QUM5qRTSkeGnC4s5mcBPfpAKaEC/bItZ12qOeaR0TEPa0SzJh6gSlXGlDFAkIdQaMB3w
eOksm6rzAijhNOkUI8d+hx7VymUJVq3BkPnjnkD3lGXFsTbEKE6jwVOn1tjWayBYpBTsJMaWvz3q
ZPmclmnBlTyGgTpnNGHVi3TgwjM3RkdE9U9x/WEarPCUo4TS5u4scwiYYinGS7OUf6yYvibCNngf
g8n71EfGlrsBpFtUvXnaPvi7pPU25+MsA2fkJICeVptt56oriA7gFoSmwLb9lJ82j+ttBr0gumxD
2+x67N3cFIv9iAuC0d/OA33TzY8VICMltnwR4j6O+elwZxkHyNinpX+QYFxevGi3foggb04kXX/O
eO+JH7KB6Vla91hvgohXAHfPw6MquzWi1TuXHw9+HiobxGwyM4NEh1DMP+Fko2JeoevpufF8KdzK
elk8iZTa+3YQ9W+q7ahuEw5XOq3v9sW6BVAQWPTiOw8sYTPkG/y3yuwgqauwwtBdvrcb8VICW4c6
AioNL5mv41dJN0q2sjMtlfD8Lq7gLy4GdkcFckKCgho9wTTPvDLzLNwwwLM/vyq1gTcpr0PrJ8sk
wLEtRjhn2bNbYtirp3ASF+q22ZYcy2f/s2auWxe7XV0YNS0M9lh7JisxkGnGV7iJiBOcRax2csLe
Xy/jfOCE0b567ytKHrK+0HsHrPh2KohgLavqYj+x89kwFbG7n3PHNvpOIchc1gsR0SKpjTJOqejU
Ly+9rilM7sn4Hke0LMK3btjTbgI90NpHLFLVEWLwTEkSiuyOv+UYapzVbfVG3q934SPiKiAggjWz
0onPKk2Y5px5w7bNPtwQ1B0pDnGliAD86PEThFeEkCmCwC7xb1WlTucloFIOidl9Hav2iNjyy8UX
zCmGVLQ2YQ1TjqtOKZK7OwzEtcD1RRSv39NkrLmh31tWCcY9lFEkTW4n2mw+jLn9nmLznhh2kbfd
xSthugZaKjIrSiUfFQ2P2Y80j59IRp6GBLJ42GPE1loY+miTvIHyVKdyOaq6WpxGYoyUWw9FfDyJ
14nXPekiONK0N/YtqMCJVWH3cQ4EMNPW0v0+XSghpTkNKekmD12uhVcZTrSUfeMkdbv4QXXGEg8c
6uBGfFF5MsV8NNlrtGPv1TBuzTO2P1XMGt6RVBT3iJX7ot7xEcTBA4UJ3KmmHdH9ZhUcBVTFl5RT
DHZBwnNcK4fZjDD+lAHGGHBp2iP8odVlTFikxRF7dqEGpkFqY/sSvZlNG7l/4IndP4y40rLUjo2h
qFXiVr97V7tyINYxXvRo8wTVlS/zcPavWZw6du47KXLM30XLW00qZQR9+YYZzOPC8bpfZUskib6u
U/3SkZTHvWZRCT9BqgGo105PY6jkLfIiLsW34FZAwIIJ608MVMNRVjOcoWB2YozmD4pWZqmuvgyt
5sRmEhmi6EDC4TByTdnqNEDR07P+MzvA2aPBg1P8yGHWteiHe/up+PJF4OtkdilBjb/vJ+HHXZbH
ySH43Ja3IqS1WsTZy6Cd+lWdqoiwUXMEkzzf3zInEvD2YYYOSyF45nAnQhsYDHYcdvyGJr0ihBhA
7vu1giVrqn9GeHFZHSWKHGC60+t0qPB/mhsGfGW+s3DjuE4yNjCXZ6ItI+YfkfcgKDjmBCLhHljG
5AnP/6Vrrwm7ZzM5/NXmIt0hscfh3WMAuwuA3H3Ir7FuTaJlntPfclxwujQydPzdhwgEaBlnYwaN
uqYxpUa//32J7UQU/5uI8xqJp/2nfbun2OR6koQH/tLuORVZNlPDNig6hqCldfqKTXfvidxPUp42
77IAFpJ6LEPIW1jU6p3LERTiCveJl94EPUiOA3K2VMQaqwgOfP5LcTsx1ZFX5oVCSDci/x/1mNyT
rTF0vJYZG+mb824WtE7zzEN+akFKI96QwFNXaFrg/IDvj2GFXkpVqDRjPUD6vU4VfCPKi/G3dEFp
IzNsK6jilQNeZ2Je4Xr7h7oj0IBVOhn+UI7/rhUESeyExdX5FPDWfMRlCtoBn5cDGN4IWANN5GHO
4rQLylWLh259BAgxlkE1/2FDKO/Db+IzrzsJo0FdIsmZ4pi05Gx918aCwSKy7AnzD+7zt36YSMj4
rBOAsL3tAU2y60coOrZ3xQ57o9xwMsfQ7vSqfdBc/y5mcNkdBxOf7v7ULNf3gRTZHmxZkjts+KlK
KQ/NkVrfedHt/RsTg6YDbSePMPu+Kr690f87ZBZK/KGhVvHo6v0thb/+x5zooj0Qs+utgpaCsUl+
sPag3iLOT+tw7L2pRz0QCoYR+QEqKDR4YZ9U1Hyw24f+OTBSkaXa66hVfQ5njYxSWX8SHSK40hrd
W34z2NS8Z6dBoC6Jss/tiQCROQhHCYttZoZOtsrpzZ3ILHm6fnN3ttBLt2sl+M416QO+bOw8ziYz
ZEfEGPmhJKA7B1+jiIkq3mMTXWfHrXuTkvv2QQgSfz0+lTq/wQN/MbbfQYs5JjEKRadDcdkfJSlz
c9yW2Kxw8aa5ggtI1H7ZAy3L8aj6zAgyCHn3lNRcNM88TVFW+3TFC82OpWJJzeXsf7HvT2B3DZx8
HbXJKcBWstAwN/+KR5xzIa3XAUN+14BB7aHZjQySAHgg1waIT3z0bf9J6y2Wi7SgetYuifyLnwXG
4chtgAot+O32k2Mbay/rEDIMWjALy+GNv2nL2SQwVJiJuK4CbEVTQuV21IHAs9EHZl5768jCgGo0
WjR/Rd/4cyFynaAK61nQuOWeY+LFiClu9Egb+c66qcFBIYEh/gzGUeuTtPUW/bcOSSvHEL/ap8Sx
UMHOIRHLsYDENNUM1tysqkSHes3b9Z37Gl+fkuLjjrx5qAmRVNabN9XRZAKHxRxiGcnyU9YsXAfq
FALHrQTD7k7b2VHCbbWwOa1nun86P1sBwXB/C30GmNbwfcyjMEYPA5Shie94F6wLoBbNUKetwlyg
seoGGsPReKG0BZ+L5wgFqBcmq5A1837M6jd13w88vGqLpDpPqaHopmPKOkvTDIChWVZ/ZZc2eMzW
JQFP6+6huzATRE2l6tGBr0qbnvBiHtUX9r9jJMqvxnZhvx2CBU2AdT5jdCdugPnwBX/Dt3bXEm7u
+MAXHDHVhzi457t0T4z44r/ZF6Cx03Chbu6QvsoL/9urkSc4tRp8LUSmg6dXLxY0jwAG18ammZj+
PDbJ4qPFQMpOZ6rFHnygRtRmqTijNBAW6dfgP1/PFrfursSz4m2a7POnShrJEScwpPT3TJMp1cn8
Al5kyWFMGD3fk4MWqcw+0d9laxyTLso/HGJIih+GDHo5XpxGlIsw0OHwpsPB+EDlZn5mufdXy7wL
BjY6W/BksfWT9bbalL6fqmkoGrbiFTcdsTcCyC4njH54Bq4TupiAQxLgtoGUO8vnPIfIlMeCJKWH
ozpRI22WBse2lJuHZ6OBOyRQezlHP9LfJ3m43SIZK1s587cbs/ggIUwTQgN+aai49ivtzcGvXnj6
NysvgEyO5tx66QZaJjgRr5mjpkVR4BPXwSo518DG48wTrtcwr1Dil51K7naiCq7q18KJcLVYN/kS
S2ZWC/sTUKr92ImFi5KRR0oLe9+kMlGZ3KNj5exNA+Semo+O9zx7BX9+yDippWLIO8wZKb9Ic54e
+caSkT2Ibpwlayh8stEv1gdBc18f9dHhf34zuqanf8l+s8HLB5zbU+FchvmeaHi1mI6AYL/6NqGQ
QS8fFGyffByQdGKZBqhLLdhadIeexbvRA2rM8jyVpMLtk3JNgJL9a+r8Y2M1/6NcUWDKvJ07gVD4
pWPP6RXf/jOtbZVezRVdMXNfbc6xl4+ACYlDhr9h9/uVBRgkHCN184xk4KKluxSjjBTbZ07lywDM
aJYNNDzylxkY3Qq4T0dkp96MRmpYV8626Ufrhg1ClQi1BhA/REPSxOESRS0OfUOUxnrd5Y+CQEL5
JWvoH+3LY98fne4oNiIJmHnGqAV5kNb6CKQnODAZdqywdv5Y9lvRVYBD6seuPClbnkWKjdaRF2y8
6IqV5FlZvyf+OdPw7YZL7qBxlFVraoRHYIzVYIKwdxoVfxbf6uqJRqyzwID074yC47YPCbnRlpuM
kUmklP5T3USqn/hRJSW4IW1KgCc4sWt3mdHHDI3n0y3Tlb+laQ9Adr7yBsXRpoDIAm1wtQsdS4xs
DaOyn70hBcuZfzqQvoZPM6VLFDU4jnHFcpuASl5+2koSFp6kPqQ4BayH4JyKuROELF2ZPkmNiYfk
vrn+m2o6tGbZjk5n6OdZl8RDWhS7+hVS7ViXTX3ByY1nCxxU30vioeNEl0SO+RHrvPMe7xGDlFkA
rEgmCRnaGRZHQ34i0XebamniIuCFFYFSP0PsAeksBQNDkvhho11oD3Y1wr19ONPdwKtUPGdf4iy4
SNpfAIwu8KY89FXAUtYSFodp1LxUZs6LUjisNrEC7+F//K7b1XadXWQIRmSwcw5dXit0tD43bBGO
aqwavaIJyUQM7Ohkzv9rZKrTZ7g3huXCJnL0/RjDKC7gFsTqx7iq5O80WXhOLs3ZDxyz9s/57D8L
KUa7w+neeNtzkJVk1YK7KTQ1c/EyOVIlvNroLHbIekVAcBN4TH2ewaJz3pGQs3UdfRAoQVDEmwYi
A68LPzmpXmEPvf4sTX+BlUCHiLsnq35pyyX8iE7QCUmd5lllQKMwlXNyuznRxGGU975vO6sh/Lkx
Qu6c9dqXMVMX17t24Q4ugua0SdYcwezniHuos3rj6fCziSWJp3USLJhwMHgs+Q+RWWoC8OqWUEYQ
9qeKFC8Q5TuaJNkX6tEc7fE85ou5EGWhpPocOtQ6A4CcAGCqWk0aLOTxcXLY5eAzHWxe8bLo6IKe
JwbW7WWnCjsncutQPyNO24cx6cgEZQURgL/oUYNoRYYS+BZ9Nh19WvCDAWcyzjalH8ooyErKojtl
hejhDfn5txn4bagoFgb7fLQIOptLmoAIqLaRYTEO4ZqO8KQ87ZANIpnkdUMDnnw5fgQxNzXkTPtK
Fvb4klXW33m0bmgMQ2XLnh2fPuleVCU/rRdNvRNXvqvcMlJ7O5mK2Oq7yF/A+E0LRauydm0D3DR5
D3nrUuAQKif66vvA3uGb0gQglP1WzEC6PYaWAfcoNS9d5RhXMZG6AhmxpO1cPKeu5TKpte7Pox7k
jOpS32U8opS8I3NianLNWlir6o3coEctzY8F/u3AxDVw5/jhkEv1dC0m/x1nt7b24yThmOaSCEDx
yzzWkK6vNKR1FMQzN5e7Dmltbwmk10qVRU2PCAICi0Ru11MCB2T65kbHsL6UOU19hnk4Tf3xlHBi
5QcthtSD7jU0fNfk+SZLKQOx4WVLNYq9u7bSWQJIJNhyb61SDhHcniRku0LD6nCnY6MEHHj9DQVZ
a28jbZG8noPQtW4k/ZC6oP0xfR2sQ7I+dUcUeBdg1hzHiLFkh48qkjuiSYkDyvCqkKxYJKMeNSWL
IP4uQKbtufOBy2oxGfSxLIp+Kx/HHtZZz7dGYZ8u8vA/3otkNFmuVK20eY/acsRcfEULupjqjZJQ
NhpXbSqWbTehpwzZUWT+biKSxT7f3iiN+23fmgtoW4PeG1NtjI8njuOg89tfMvfbAOxe5zu3Vr2O
vJ1vhOFWjIiS6iQvetPMKDVzCn2jTLLkbq3QKHqM9UTaS6rxc+wCnq4XE66Dw4IWlTUHFSbii5cP
Lons/HenQSmYmrJPN8LtCKlzYtvCqXm0RHCVbdghKmsZJ1zRSzdZx/CPtjLsZW36XKkDHt1SYJ0q
3y6+25ux2J4+I+sDF3tXndOt+VDfOCylfGYFx7xiy+YAhgBjyM+DQfWsrWWIkn5Cf845gi5dZ57g
Cwfw/dngOC0ZAdfilc0ts3RpxT38VpvyWDwBXNfglCyCvUXT1B1uBaRCyq6FSJBaZMIeHCrOvy9N
8/GhiHkGpBc9NNdp9NJQplVwMQus8sRd++n+hxJmrUS9OEgQKPB4TXoRe7vDxGCzmUxAOYkYlzYk
yZECy5d73stQFslwMVjWc/oo2c6/husy9svzNVy2oGZZrQuwzgh74wNmHQgyhL0ylkhlK94z8uO1
SA91OYwtvajn/gV9dLakU5zX/ubGfJLOemr/ibT/B4KHnPQ/rtChGaKdvSMl8gRRMLS8pL6wc7lS
kaW+KZHcJH4faUzISTT0CvIAZDUOpAamgvfOcellhQM2E+cpaMBngBnDx1G2V5Caw+FoCrUy7vHL
m13rNeCJZXRvK9DLlGHH8sC0lMdFKKuIBTxk5iuojezdS6fIblcAxIBMdG+tR7+hDoP5Jii1DDSY
oaM48h0E4jOb3bY84A4szKpSnz/E0Z5LAuO8BvOQuM2QPh/h3KM4die0LsEY4c4Cd+4GfuLbVUPO
4KBUh88U9JdSqoBpsawgOFwQrAxxbifiJ3to+p5NRWAgbt+d4RTVufs177s7Y3F4zzGT2c5MuApO
n8Q0elNlt18Z6z4mY3noigOjNvTvCWdMkwWDCxoDNSowBQb5vyoz3m9BUJNera7Zk5giKyD5oCRJ
iYUZXX+5JVcSZU0tqMNJfa/dF4ZrcfuhWxPBgxKFvy2YW3NrSvFDisuCIOrdHOsSC6c/Ko+Z+6K4
ak1K7/7EoV5K7C5wM3G3wdvrngrNDWY0DmltK6uIIQSb0f0UDpNoetmAtYxVetr8Vr65ag2BUWHw
QwIG6Q0nR3T1wMQki14Whu7Dh71tspI36VekpMQI9Lp9tYXlfvi6iCfsxGRF5a5Ff/rhXE1BC/Xx
GUKDh0Nmeot0BNk5DdjU8NJKTICtTYmI7HAcD6lRyALyYAIdsHarUhPPcI9oVCChcu6AJRBLD3b3
OGfNVjQPD7Jf6FjhoadQJy0VGUyp0iHYKVRkDyLwLn8oJ6OT+ZCTTSwOKJGkNn49f73S/WXpMZEA
1Q8I4CovoM1tN6ZU+s7BVPPrRQCueOxtijD/GKx1m+A/yQ4KItQZ4yeSUYoc+/PW+HFBsL7ZPSuV
SBjfZH9C096/ed5DXkTcYU3ElA5I037y7KI5lZval0Io4G7Jrdnyt0rVkrElp0gRXFQpYTLIT8fl
yBrEX0eycHEgI8nZqYiiPHxzixlPjtv0D7zmAXt7DccA0DDcbUHXeKVixjGV3KPwUfm5EXsf0Y3j
NfN8DzYY5zv/NLkqoQPYvqRq23jfGjQ8MTX4ymSVfIXz0+XtxHQbJAsX2VHSB2OnFJVsmMfuzSv8
4GfuL4rw8Kw9pJAQtgFpjLCDbYjjl19TsT66ayZz2fNsle4CXblLe2k+0E0uCesBQNMT4pTIRTZH
JwMd+ld3+4tc3TImLU7ILewuQNsd3tT16zsjEf+aqDWqU/thtx9Adg910F18XN+wYfFrES7Y0Pbt
EzWjoyahPsQSNSpz3msoMx10YKOvqHVYrCD/NZj4mb0zvlLF9bpDG0j3TmvkpqXZs0rAs1gH6f2p
xvCVOm/6vG/ajm5N+3BMJEkxdWK5xSvED7zEhhHFkswsFxQvkQ83m0nEWtCNZeb6c/RT6XhAYMIq
yVv+QlCooW7jCp0Qq3WYC4BG1fDG9uz/vEYar16dWLsbqZYxOCop3VOJeFs55ItvTyyV9v2GXREh
Kt2I22fkb2h/7QvwBpEntpaXLr4N9eEI+v9EYpGPkJO9DWIeUw3BfiMMd4mu8mhslYGXDtBWCE9T
Qwdv0GFSOTV6ihtsL39x95N5SDkS+0+T15Uipw2oOThVTAM5YOUDFTz5G6XMc8iLbPjSmU4NmIqf
3Bkanzh9ghtNwIUoS+0twAbkgJK90oJ/LcrbOba9zQuBLfusMo445E64AwBNv8506fmoG6x3Qt2S
iLoqKn/htY736i+Lq4EIwkLfN9atXA6zKB6W1c9mAc86c7XzeIOhEQ4uTLL8loQeyZPsJ+EQYri3
Mn3by6gvbta+3YI0f2kqpn/iZ/J35USoN50sZsOaYqPVi5d7WuU6mlxy8Ou6TYOOrnlwAAnLmgXb
Ck7MjMV+f+KCxH5gUlDMCYS4yE6SniYZ8QcWTmnoDoQIKYLXreeTFQ7/dNdcszilUv39Whq9VMmz
IaANBk+NplI7eF5YFfOm7FttNuFIpfoEs68/xAZg2FiVziH5atNOlwMNhLXOG/oMY/3LZVG03doJ
0JVZkhSTWPi6l1xS43kz1Xdovid7w8mvCl4hdUrXrdGNdVU0liCi5yyCcq3jCX7Su/WmuBgeaeC3
l9sZetxstV4KbAksYdlnNdPCrtIkdhfgpj834iWPFVVl3153kiMFcewXaIXp1pVYXFzfMmzt3kvG
MRAZVLMOhMDllg4QcP/CmjQ/8D5nLdYiC4cn4ZlHz8zB+wjbkINFVEetFe8YyPQXas7C9wj/Nt/K
AGahkHhQRJxqfErdpfCXXt/hIVgXjJOPrqJyf8iqw0D0UTFjPGu/2S6fBmqF6zx/i7PcG6Vtg9wI
xFhJkS8MLI0oHEReh9Ix+Y6WpJX3FuHxsnWINu5xOQ2nrtBVLbW3Y0k81dx/lJRgNVWJoCiwt28p
fz6hYUsmShLewk1VKBsUk2XR9c9T0Ffc7DSFrxNe9QG51YPRwv3zbO8WMTjDK7JhHjvfc+tCEgH/
MVeshXsmB5ULxyHmQIH83YH06AaONQDh7DsZ+rsbVKTm2riLWu/vuOPUcDGTUPSiSEJ7t+I+tyPe
JlwKXD+iZ5ZxvRf1zPE61aJ1PoG6SBf1Qavq4EHqXOIf0I6PkOfCtneddB6x7fsLnEBf9Vuj7IZo
g8glM0yPhGlaAcZlGm/uvJWnyKTxB0b3rO7TO0IzCjXfqzKvPaplDHRsF8odm2Gnw3IX7KYoBePv
Sc/C0nxNgaOKJEm2pmVKjBLGXkRIdv/Zaa6ouJd94+DLCyIBNk79DByP8tJHmoudxnXqL53Pvhru
LPy4VVOBn5kDp2oQhZW9z5+M3oG1aCYhW0zrUEFmnWetzCZzHc/Y1937PXdRrLbLE2c8R2rljYKX
ufJRy0wdro+vq8WWMvO0MHmNLosqgm/1jFQce7AH7HfDFYtvsjivf2QSPNvy6rt4v4kcDI/deibh
tuJ0lnJaUCylSth5zw9aZ522aRA66ibqyi8iwK9BU8xdWW1yth+q/gFGLqphNdm6VckAxOFF17u2
98Om+IW3jO9YbHLwBbi0ncc4Ds/Epj1M6d9N8McnQ7oqKyIHiZkzjVxTZ6PZ67d+V6ck9SoXlOSE
nJHWucGruHqp10GsSkMCijov0iQAn3DP2JhPNfsgMhMGQvAWksPoKHQuEf5Zr7YNobW9YLiAW8lU
Mj1J2rLKbcfMXtCLd/oQxXrmdh6Ee1335Y/gJT20MvotkZxPzi0Zwy8b4PihQ/e3mioVrwVShVbF
x1gu8SUD8Cyzh5atZmQKLD0Z5egyKeL7gzd4M4epgfL5ktCeu8ivbM9hrSvKh1PKE+x5PhrbsOAg
AqLOO2rNKr9eHIolREwyJGo0jc7OjxDbHF6md/VDdSQEMENfb9IC89HfgF8Asi4/yuo/631EgwNB
+BNs06uwwPNekaiQPHi8t4ftzyCUe7sVGqjd6+fcy6es1Bh2qHCp+QtM6ORfTI35SU8B18sPiv50
bL/yC1r/LhVpeIWk+/Vm/4s302DjfSbYy43qYdeG3t1yUsL7wy/gIo91mBmKJdTJiFiqTSTFgK6x
xcGmnQxXksONsfmjPrs1cHiuiNB7GK++ywqnsIh4GYtARXKVh4viblxRLy+MF87wqJQ/4VY5RQW3
A+xsYeamKWQe6indnfoEKdFefizAb5OZd0jCusRlYeI73v7/i34BfKmqYZXimBcZubM5Iqi7keYw
up62lOTT7EaTqCfPm6bg/tezmKQRJ/k9HWxhVoWRcqwAxvaVUuElDuZ9djypV2zjXC2dFgca4Hrt
PCprFYz9+rC3NKHfuXvzVKAJg//O2KPpCtdhPvtWGdCcHJiIH7Lc999RCZRW8c+l81tisGLNkCtj
+BZ06Z3lVG9dZfssR6cv/fmxuXKIrbAldh6ki103yWlbQrgWMn8DITpwWmDYZz4ibiA87tMf8QwU
XfLz3LklqjcIAsOOsy5ycSZ//ZsnnZXTyGoeIHNpEsXuSqiPDoxveQ/415CeezP+tQHwCA3jCA3I
RB8GZWFJqC1RhpgYqgIPm+Kxkr7hTAYiX78U2WW3FwUbOmNs+S+rQcAvBZLWBZ4d+3DJ61UhOUN8
TSsCbgh8uLdhkqBCYzPWsRCDoJ+yf8ITRQo6HvkrqWwVqdR7d7H8bajOa7irV6TK5gETB/yn5jnM
CXpqGeYipvaSyN1VqeqjnFO50Urud7OZmZ2FikE2oXH+FOjzRoiG7ThfVPRvw3Xy7w/jbtQVNRB+
Pn9Uxyobwmfa9Q1YZ1G/Smf1DBOUXgHnczvy71ROaxMQ3BX55JFqxwHaIxolyDuRptXud2Vi3Jar
J2zu5LSiRmPfOrhAAM5agqUELZRqHoopsJI4P2nKqzOlF8nU14aLGnAcFP6MgDZreGA6n38LxNvS
1psxdtq8kiSWKyRPQFoG8cRJLTJY0me3tgfGbAX2D3ba39L+FEPicsG9uftkm0iVsbfCCDJVtrXg
x/OADsz2GcBQujx/ZYwboKN3McKTOVCdIDOQmjzwAThxfKapBBR78Eod6SP4s0wjPWncUBCd3nCs
rhPuGTsfCZnhL6vNBQPJhElgktfBu3BrKoEsz8lQwf1SaYflPLY4eQYTSH4onVtS21cvtuKdA/nD
2LODh9KrxfsbFfBNZZchIXhBXHKimHJTpVJfscn4olAXUL+y82dWZ/nJTTAUci52gApEvMxm5j2w
X430NMS8uk0lT0oH/BClHuPpKCrLY+lAIkJXs4e2ytkNGGFy/+DF3reCQmmROAoWmhuHsfBF5tWD
+CPDUMlx2PybLgkT2PwEW0kp4RYLy4hdM1flQLfculy62MXkpdq6atzxlzzhZwrmyPEzLA4t4GLu
upxLikcIECux8Fd4Epo4Qs6xPVOHiAmmtzAXQyQjvJC6ICPqeKbw887YzGRgOTnfX9apeO9rjZl9
mFcu8YLSMNV6bJv5tWaDfJ0W+K7NfYtID6CNa/HT7OXArjXSNBA6mkqYAYIjyBBZdQcfyg6///pH
OEbr+Ot/rdYFuJvzUHcjFcCAWyffyGKtlwhEk5IRmHF16ylKof7LmhxTY0aqS8QkeU84d90MFAvt
JB8lKqh89vrB5haGGVrVY3uF/ZMG+vRf3bL835ccnE7AFIdQRfHvMhY9iTIwc5dafd1UYQ0ZTwtt
W5WojfUH47M2UUjZr41jdKhYKGUJBRuu4UWCkM11rKtOtS81y61UfNr7I/fQg27NusT2572nY3MV
YUVs6YGktOVqiuxCtraPMDpVwk2QxfIL8FKg5/lxJMExFQ/9fF+wpr19fhRW/klphvYKdCFn9vdk
iykm2WEFK99NgjLkBWD1afNO6LEALI+xiBXIIOoy4GTAmfxDFcOEIqrwcBQqXlqyzb6xQepP/Npa
k/SqC7NfQA1lNtYQHFkFEcHHOImF+XBKXFnh6WFxZSfc8h3OQcZIJEWqZtpORgdf8tLtwmfvFvRg
qqKdvQtssG923lkXnhB3INCvquFMkFoKwsJFdXEdOBIua4zwyOsn+HlKfcOHM5BqyFdxR5Rj8UCl
fZg3An4j+NZaQZK5BgJItFBgAEWkInzgqppWssPf8xSgSq3dTXxCpEIw1rMmF1U9qwO1xiAgRT3C
/ZsndaDwWkmTEe8s6bCoaoQkpH+UeLsyjDKNEgedDMFMfzK7hbevtTjDUJsUDkd1b3r0osPOE51n
zIY0FgHFPIBBVPtF6EwNx3wqTLM5FEs8TsHJqruSOfrdLaC12Socq2R9TNxuEUC5tYr51ndbNo1D
qf/h9XjbUawAvwqicgPv0kIYUV9pQ0cTsxa/+m9+RVysC0TL7cU7pVriUii+D1jQUQzXqUTWAH5q
doWveT39VTvpDpmTlCUegFDdaFzE4AKtSUGIrRRv5+t4E4TZeSfV/WzWKu1+5x9rDfFa1r5RWRO+
9Gx0tSmh4PFYOD/T9ao6pddjAVqL5xysMDhTcrULOXwA9LZmYpVLmR7IQJsL/wbug6ld/6eDtpF5
v/qcIFz6LntPmF6MnAqPdKjpcNm9gwg0y9df4KADiCK3ixHuoT+QcXJyBFq/mEL+sfopPm9fMxpq
SppleseQ/piFaJokLyYbZmQ+st6xsMt3mshE9VFOZyMZZgi1iZOryxRB9nBasSkJvbOW/urC55KT
DrQHzBiyt0zNeiV5sg6Uwv6k2gXDDfBFWyHrpTn0grYdV512sh7wkODvRIZIJnb+UIsfWZ6HuhJ1
1xpt2Oul0o8ZFeLGTLzPzi20RyDXt+ekI67kyxc6oP7wsM6sS73UsHdHWMcvkPop1znQfbZB9W08
6GJy84aCTwbWrobzfujEVY3Bt1B/M2SAZM90zM/fya0E8s+O0fkYzO+weIM7eq+KZqLatkERxQgT
d9c7y45E2WQf67Jbu5u7bqPMeToV2fX8aYtsTQFz7To2mJ6jIqVkwdRQFsP0D25oK/hsMS/jHiz/
UbAbZ9eVfBrRg0bS5WqUWFRXGwxQ0Qful0GGCmCbPoV+NLQ2OB9Hh0oB7F2l8PghTcccvkGgITcG
otxFvgdOj5dQHDopP2nVLrF45WioPeDd5dZ+V1ZiR+8kAyziWsiPmQ7wbtfTco+wXtqwGbG6hm8k
nPhkfPloSl0NTj7gRk2DMJdp0y56wXxzLji0jvMD8vXSeXRPVrTwxw0ee6UWscRDx5/oL+m5INVV
xuRKXwzRQyyqjXEcEdxcccEa4TXALvXlmEgXqvEllRqgTJ+bBDnBHdgP3fwtTSjZqhaIhlgUIHFD
m0+F9LDWwkckBa9VGqUbPlYttsKpqy2FJW8kVqLokb/2IjhSw8kDuyt2ejZ/9fdYfQPo+fdLlQnx
8swczTl3Ew5utcLYnsxhTL6JzLn1AmsvBMr54/9D/HosQKQ73soAJS7/2+5oWfAGc9zx9L+TzGVk
+eLPGJXenP3D/aUCfBs5VLM+asEHanIWmRtQvsJeRw4U/e2jIq0Pyr0tlf4oHNTozsmRnSF8xwlA
xxHYeMyluFPLqnTsahobIytXvyN5i7Gt8cWonuC4NcQMsMGtrf/PtKVW4rsTikmtd/fE1oKZQ+yz
U3TK4ikPq2/aMz3KMHaLHaOKfdxKMWubyagOxJipqu4AIkQaqMBpJr6q0MOQ7qjPZxBaToVleF52
eXzr1H6v5ikoY4V0v4PG1Zsg72M/CYMI6y5zyqSJ0cssa864+Z9yOt0WwUKsEAY9NwMGy4/t+Vhv
afMziS9FIf41e77Gtv99gMg9UeXezcMJKaE8mkpOhiKyr19tle8EmhlCxPGtMMWLoDfEDcMaSd6d
HiO+CBT/RxE8NLPtE/Ymq+0J0vQsPr9/i4F1WR4OrFa1tQdvaN9hIBWIrHM9s3JiuN04N/g8LAD7
kYJsHcU0GyNwD/pJuqcjHFGZtdtAT+IezuZx7ly+goty3ATRK/O6A+9DBDx9tKtVIoUryY4DQSUz
dt3BvxOumkAYMWBAHVXTmMCTS8BJXEA8BZkRmUEfFY/EcvEWCPS5Zx3Y/Czo+O4n9v8PnZ7bhDzC
5tXFybFmMoXNxuqX/q2ri5OMQmxBDlWKLHVe2xuwrA/kKGj/BuAdYmFC6VV+I01U1r7jxx4B8P/n
eHp0wbvPzQJruPKsU2ZVzzuYz2Vn8aGCtgO9Q61NyBFWkjEposTm8ZQGm9VLryP2mr8pQ6k9naTj
fYcMATFS/qT/rCTCtPOP2al8wloycFPXiR9ZrkzvVJl2HRs32DAaWIXxRDTqJH8vxt4ounRj9i88
MkikA4qZt/7NswPBqRBqvGoZ/3RvVPpd3yPnvAjtZQJoGDRDz000SQv/c2xYlll6AaFMfv5TPkw6
IWD5ZfMd8hGDaTer3cnbTeNsR2qzb9qALFw6EV1bPb1HbuRG3U55hMQHN2Z3UPTBMbgie4OCWb8k
Z0rMsbw4Qn63Cv/UjiCyUgH/4JGuNWqstf5RVYUg/qQTK1/O2uKCTqDH1thGP4Dufazoi9zIUiwp
+05MEKirxWhweOy/eNUNRDkT3uV84PDga3Bwx/a+jT/WKx5bS+WkiuyxpGeNGc17shL/7d0Ln7CI
SMoNXvWEraqrvidDr3g4vhtBhE+TkKbIH3ftUKucDUVJm5DOfvYWGUBKECBtdrVw7kYr3kHHKlx2
FPq+U6Gcl4OLsl9dVXD3aWqLpoB6hqwT5Ck4rEHzrjsH0ddMFnYAHllQWgTc2oruPqz4TMc9EQQ5
0vxvRX12ASGuMuiIlKwJo9hgntgQMVQmdACuW6a3R3Hi5r+iZxqO0YjWiLkv/PLQVGXo/xWI4vDC
kp4bz220J22rDUwTx/U8i72HZxwWDuAxWTUyc+TbBTU3wRfqKgil2MRnKcEPPW3AGM3/IhePtVJj
Lrr4LPKyBwKE9gz9D9BwXY8X84p8E0WMvBiUel3TbqH/fTZlO0RP+nd/RGaSoWuXz9B559KaqcJG
xr3RZhfvajnmgwWmXcD9kGiWGms2aIK1unWfJBO6K/HpsL88J4bBWNGkW5Bd2pjGT0XnQBNDObs7
dX1/6QuLjoZTbQKxY8n1CXdVFkduO2Bae/z/qtO7HAsSpdSNRq4c8qsjPpy3vXVgshRGoshoVrNB
2i+yLZxXyq1IR3qXZXZG4sL1uyrir2OAhSzfCfg5+NM4LjM+LbJ/ke3BcTqLxnZsNlAOkE0ZM1PA
HRzTwBwqigL2ss++7DWW6MN6TOPiD6Wdjr6m8s42/p8+z+cjdNKYEdGpEv/DTjLjcJduDFYa5KMT
NZo48fzi+7KCyfCta2xMhzxDpANnuc6rOK9NvBeW2mppK9pHj5a2/lnBL7qPcKRQIuyGc3K5JWD1
MpJjmByLP+SrqQrmzVvrR/qktAUsCGPxiGlPohJ5rvtEmlMXBnK4o0vEwtq1HK/LChV5KkGO/mgQ
NS+gqlNtQ1tRCndvXeu1jwZu118shUqt3fEXMs9NpIuM+65iET5PuNWRxldnsLRnN8jmOX/hFaP7
+jiPq7+MYolfsS7fqXFvjDNl8iysfeWpdmSO7VwlyYCW3ggaJ+WXgRynPJQUFyZ00d7la6elyZgV
iHuLyDpVHl8u1r3qHLnzhoNdQzLf5f8aE0S5Sbpp1OZYeG8sp22SX7t00Jwt7yOvA8aVQSIsodSh
0zVnzL1uX5vPQzfqd1TPvOtt3ZcqqGxb//IdBDUAeGI9480nkZBnC2sOMcDcfUtm0Dv1AlCAHj3z
+AR/fk3bykNtF+606Nmf2RQfILFf4hV2J+w97E5JNL8QS5ilos8Aovxmt+D2xEP/U6nF1UKkIYTU
K2SJTcsfFpOdn3/5yilHRzzdBn+zsPS99np+BocqeuDtce5k4JbcXN3LfmmVK8i/RHrgVmDEmE/n
UlhFLpWeEAL8dNZCUZtqYTNZdH9l4z7J/fgTkMp//FmlPuWUPaOFJ6zIJWpTEEidFtKEzMnkUXxv
KAumhwVrSGqWZZ551oKyHLaiKx1gIF8BusNYIwJt1yf96dUmj5+RoGn90R4l9Q4LHfqjw5zTlu1l
tFiC3zNZfvJYJFtMImbERP9IxAy/7Ityhy+8eZjncTFDnXoyw4UM7iSQKIEbCsJ3onFcm1xqF32H
ByFQUOYh+qQ4y5eSLhtLU+8PPsBCKkU1e4duWHl1/F/lXabU2Y2mUEse6g9YbM6ZRD3aRDZwhutR
hnvV94iWWd4CIu7Zm1rw5L52ekhOQ+gODw9OyWcnU3atRuI0HYCyAjUoDZMKXD6zmr6V5wOqMetd
izxzJKnwBrScmijTwtrS87iFACZ0bvpRr8HK7Dp3ME9NW2sLkrahFhqk0ykXfAy8niJn8rLxQUXY
cn/Ze6BvOvKpuqr3j+4WHxCQn5IMPi93tZPVX4ao2IMmAqggqzi7U23SQRD3xvzMTQRH6D2q+qcC
nNCqjPHJqI41M9MxrdexG/pp3t/r30hPIjivnWXS7w7iyJCaclz0UPa9MuzIXT0SXoS2r7gIWsYI
dxp5VOObw1vdBLlqVyGRb7qNlfVYNYmXZjeBO+adl6fVQRY9AY6ouNgT95L+DG0zmvGE1NL4P1U5
vmxOgWWzTj1XkHBiCrhdp/OPtEe0i05i6ReDg+/nRS/UJfOCVnbRjVGaTx5tab5KKF8F2Q+F37Bl
22tAIRkdlEUeUpiNJtsf+FPi5LAtYfKCFR4mFiUiahLITm/uRn//NQp5bMKs7o7lK42zSgV7X34C
wJL9WOMukjRF3mTjDr4z+bjRxnRiHYLReNskjuWfeonwLgdcv0EF8kbr5DVNTI16XmOjV08wGTsI
BiJsKv5f26lIn4vS8JvQ/4qaCoyTCEigj5/xyPmpZayDrUek4+3s483B2vkl/zdWpIRGzutDflJL
Hc7EgFUlUxhJd48PgyPSYm4seFmQsFribTuo6KaJitRRewYxVFJa5LUAKLbXaI264qDKuLAiNKI3
1KcINBwSx5cSfqaT1SGpDSFQq4hUKvxd1/LY/HMhhuch7UVcSdKdCXoGZZgEnptMWPixBWxGbZo+
Sq9fy7VfsmbCo/+v49XZp0QeUQ65yJDkeMorFYSSjnF9Hdc+mxtrNFKyzvq+iAAOGuuzumXLC0B2
0jeXKze5qZ5Ao8wD8atYSlSqaurCSGzf9oz0GY+47QANCbmfD87LC4x8ehM9ygYVXE0THhKllBE/
hxITxtT1A+7VkgaMyt1OplQd4Ji7O8dH4OsdlEvgzQNyDYX638h/lwFKfp59GqdkVh14H76XjpJH
pfFxVR97QcyBaMxh6PqCPEhR67fBZO2I5p6dhAX1ooIE3Y2pQSNG1EY1DZm8N9M95q5/xMFQYr3r
XSrk7Kx2YoaZaW9FBlbakN3WQGjetOtGMB8+l8+obFat6r45x8YTxZ4g3VY5EULhodB5Eoyk6EmO
e72LfuxteScCd1s0X152nVwKwrJ4zVWWOfjoei36nBTZC/ZZaW5P1xiu2m35OTVJb7ZjXUNqXIJ6
DmKKge9BbKLVW76UglXwVIKJrhofSdwc2xTTjhjgKJvp4Viq8TDbS3VCAfDNGR1eFUJZoyYhI4St
iRB8l++A3KrknzAXzbJtGfWxIT23RpauAu2NpnQR0QVPYySKfg0dARdRzIunOY7etySZsDHVSp0L
YY4yrCPvvmIaPH1JQuJvFhcOiIt+/J0bojgQTL2o99l5tT/ooS1KBQEWhpIGRTf/Q06UVSuxZOkT
tMSPK1iJ2+nd/hg7Xx01hgK/27ruqV3mZtPSrr8DGPy0N2CemCRv6GbWIMbbKyGkCZ9jahIU1zFX
0fEuAEhe6ACppSElo5qpnOB0Qnwi+EEe1k28lA149siDaSw8N1IC+DAF400owQ9k8OvUyulS9C4x
WGzWpzUQrY7gWxxAKQJ8CKpucmM1oBQ3ozbLMhR1CxldQX21OVp+VZRCIfOPTeULliwxexSWOXmy
ihybfRrsMfjazElBHy+ZeBwzo8qsz7e2KNr2MIkIS84V6pT0F2MAyn6vY0JHMAysawLkgu8AiFys
KBIPczmEIDS+yeoYAc6rR14uIO+n9vnlimJh2TB1QVoCg/Mffo7vWkWAY4umLj78MUComJB8hqVz
iVh9s6BIXR8cyL/cYg7SwCG5VVBjSv/KYIG8eEjAA7ZwU26lrLxXxhwzwEQydlB9YyLtBGlhNzZt
KV5gy5rgX2Qk98qrKvmk/kdgFgQuFhHbd5ssPd+wJJdFchmyARU+d3gaUxnArhWaqWSavhLkbskN
5RePtqqYbZjz5isFBIxMebbJFcvns2UoFMCLREPQvz/tFU9wJ6QqbVsCKXC8t3YQS/IVIAYv0F1F
8h5S0XIy/my57U5wl8sAMhCa0BuJF9Prm1nGvw2ICwRbUcPxcWzOF38XLqpYanzyCzf5FoD3Ydpq
R4OhetmKKS8VT4tAo+YBY2GOao7veYvkSU8IRF/ZGUW5msM0ouxwR6e1o/TF0a0K5Kgl7yqG5/5z
AGa574N7BBgPkEnoPrnS2FPsvteOLgPiJWkI51tK0TXh7rk9hDAC2GQPVU4TQPxbbIFQXC+/72fq
IjFhuA+NrLrAu7jHSAujpfhlBcwlgCRjQ8QJdZ8uulMNxYI+ikw98nRUJMdi1C0Jx/HtoExXYPPW
kVmUrZGEHQwdJKymLnZOqehVN5FaIiHSie6hOmwlS6TBZKjLrR1s2/c2O0+u8Ymprnj2HLxCSQ3S
Zkj32qo29PIUfq0ZmO4ezR3jc/2ByxlesiO/rCTjKRGmGZJE2Y6SwBUpyjKcn0R7afktmr6L1DWk
janbnMCXapHt69Lpsdahq5LM2pgvYTqea7BnQm8D1RLCuUoxmMo33CHM53j6dVkvdhk/Mcy2fzfj
2A4Oc54nbxsHQuJ6ewMRRvAon4ARB6XYNx5swL1ImgZqOsTBUpWKaxNW/QN1jYFejDYM6dFOXLcN
CIyV4v43cEwzsc4TmEEEYih5H4X6tnLMxjjclzmUiSScIZleS6tqsaYaSHivmA+jPPZLGnXj+pwi
3eQv8wVApLHgP4ozzZB9ZE4a3Fd+mzgAWgRDZDynmhR0PBAnZqayo2o4RW4Q0075qncWDSRaHjhR
rmtHTzorGJyGuBgru77UTUfg222fvfGpHx9L2k08IMysyB7GXJeqbUQT58oJlbdw6U8n1M8YqlP9
gW66vfzMaT4S9knOe+Q0Y5tkPc8KoauH3c1BMGlDxIGpRCzvvgsHDhJlad57KaVv3YjZu4JLA83W
Jy3z+SJtAHc4lDeNfU5ClLkyROvfYBlWzC7vXDAvIvJc5kajqmR2JdMYy74jk1PUFRzmgcGoB+2B
x1R5ZnIfGYBEX/utGeclUPjksTzJ35mnLGx9dsYtE2hfpEXg6fQxWibMqlddCdLUuvjX6TuE1D7o
kzur+Bva1MfxndWJSExqF8bVNeHLxqpOmVimalhj9qJ2JAfUhgCwuLq2VaF8V81o6OwFydesgI8f
0bWOkJSOGyskAScDWHWOh3uiO/GQgUtaNcX4lqK2kPjNnq3ntss6adjbRPG1n+vDbZp3BUjac3GG
Jsj7+vAfiFvGkwK6xM1N4/uwoxE9g0yzOoW0RMtXk992LKDqFjtTxf2VseGLqI+FGL6b0gtAn+ou
m179AuX6EBuSGb5DcAlxNsXF5i8zdIgyErdGSBHFM9SNEDdvqmfNhjzqyaOzEH5Pzb/XpSB43SYE
N4qFGGAYweIMUe2k2Wwm0P6zZvapkpanY9uPPntZwQPWWtpdghu3JWN/SyKrCtvKQUovMJWO5TlR
JlDAOiujndHLc4sqmnH85vV0i18dD6udDfae1d03/3Gaoqb37bO+ETSf7Ejiy2Mxu22YGaObXKXB
7Ap+syUZcKHvtktK2FurQDg/vdHXDiG/d495CravjdRSNUNicl4LGGra8x1ISkbegvGY063666Ld
yWU3Vgldwa0oxkcrKs/lrztPbBIBAiclI9jaPG/BO/iZLSO1V/DB5RZJ+9bwERXTKyenj0MIVY3M
bXFOc6Rhq/zXPQunZS53OWHhgl6C61+4kCTepN+Es+LKdRWR1Lw7pr8o7CdPyEWxz2goI3H/uGSA
4PD04L3TcuDimvhthVhawmqmf4EB9yelDtYPpvAfYAR1ln/E6Ol4nY1kseISo7LXisAXYRJuztbg
zCjs4EJXlLxTQh/U6JTNkYsJQ+R9LBStk793A62i1QDopJnAh2UTN30DYbMxm2luqSCFTnCtExcJ
ybRZO7Iu+DMKZY4yEONtO2xoC8ehB4B4qoeqSeDcD0odOuAGJYTTSLBa4z+TlBuOwgNfcj/slnl5
hypeyXO2FKrH2QlVZPsv1gv4Yyfgc3GH+Nzlwyd8lf26FF7oJK3E5MsdXeLfNOLdkT9WiI6v5b9X
1CiM6kLr1ZM8BXnIYicSx/qjPWa5PtHrk/aU0ZHKX8wg5gOG/2XEeCgdFvsGMw8R0S+W3Us/c320
dzxOPoHwFWvkyQBpdE3DS1P02w0vGWj+YwIJJz6R7/P7+zqf8eg5rEKAq2k+w3u3eEqV+SR65qC4
a1hSkZToREtHacwqm/jXfYQqHrz/Da0YzEimLgPKUJX5jLVY0BEcu2b/8pbZZCwdJLNNZNBST/Ng
0o9Kbb2tyxPei6lRROTqt5h/pJNegkvs34rl4/7E4eNcWttT11SrepOd3XacaCQ4Enkk4zKGaUh1
hDbTU/OTnXcRDXwF/QQEJF3XgSyahpHZMQDp1vTLHV28yAxaghBVHhqytI5Nh6Q6UdIIYzNBYkwU
tFR78mEjAefiiKLQRvCJkM8l4cic0jQzvbYAumpyk/OVwbB5A4M0PEXKYg4Upq0Mufd1/R51panJ
NLejN9gRZQ7nu47/LQIiGmiADV11nyDHpXSHGno6SQtSmX2cUmNr5Mfz95JEYCfOm+5QL8qWQOeH
FotZA3YUMSQ8XNSpz/cj+LbDrYjDuEeIzAV4dJbkXm9DgAT673nMpADMwwmVhcVmT8dIp0P8gcQF
Vol4aNLUiqoYEX4Aws1rAyHB9uvrbj1GsOKvhwFTALLPxxaCj4jZv0Zo1oIvzq7p9SFtM115kld5
ibGkW9eN5bZU1pcVwF14TNHffaII/oj1QlLbia3l4WPcNJADwZK49ExmeZEpoQKfCq9QuA6IqiEE
IKZy2zqVsODvIOMT1Daj1NOmUFu9sH2Aa5jBnbCEAxfMqLBbV3GYVko+jcc0x7DINI3s8eVVdrqR
9ohwmcWs21olgwpszb26ATw2KYgcJPLIrD7dF01PIpSvl5vJAwr/QA2v+pJtxavOVAUttXO+7gpk
5iwJ/cTO1pGRF36LVy8PuxDynyGiQiihdtk1kXwd8IEgtV8y+AvXbq67GRBfYWxQZ3hVgbiMdTny
kgoetE4IX6T2Y/5l2KWYIjFA1h+RxApYBil2s6WEVBN6EpDLo1MqNNDQC7mt3bMScU7e8T12/vAr
gvR9r2+wLDH8m1Uu3v7y/LWPEWNL0afWsSeZdmqLFiOHuARDwA8wQKwLNoLYWnawhkdKqa63l64m
/yG9zhZjr1Tt8DTKX4HJgDuvWInFSyIxBXgLMZidCVIOWwzwYJi6G6o3J63NYd1I+Cu+xS2VNXQ3
xbKVpn6OYg/3BeQJWLZBmCh6OwdI7aTcMZX99wWXof64AfsgQ7OUkfuEZACJ3Wf9jEnnOp5ElJZP
h35ZoqRVbvSK9BvblmZx60jLBRGnLFNrGNe3pDmquTSdTUnAZQ2s4RRB7+E0WLgNjTLVAE9jIofY
dntGWu8GXoUniYFSYCSd2mxAnKNI1PbjjQutHvlElBBG221TWH9Up2NVGPfkfioOO9VX1XeUS9fd
MWG/SEKTjhca97R+ku5P1tix100ccT/atj7HzARW2HnzZ8/ZGLupyWh/DlCeElhzPZv0MIZqbCeJ
Ihg3UWjbtsPtBN0IdvCV1tj50/uSDRy79G69eA6wIWo8+jdGCZj/R716nhD4tklpm3lOSxFuzQbF
lAP5KN8ZO3zNJVQxUCKTANbiYg9CKzmgSmxPGfsB8Ydp1kaaVoGLRqqimpAbl5KXGHo6YlwY4zk+
4shIZZH73Fp6NBfrDtsU0NlFZBxNe+sHcnTaEbTlj76VMhM74J4gQgq/tRN5TLx0wmLK6icxrKvh
+mqmkKWKXvHleyXiOy641kpnHqVtcJ5vK4qkoefX/RbiX2tyipQ/ZruNj5IkXWnnvZvJ0UtsNsh3
G/m+3Cz5R/nB5skICOtZg5uDvR6kOyzKR44RHpt/VWCkh3DAH7eP3/WlXtJcS4Bf+L1DEa6HbI3m
u19xfchPn8pP+Ke9fjo3zd9Y+2nsLRxBDqiO4K3Z7GN+g8h6K97GVGww5np4gNILajrd0kmRltLr
1OlsYWafFNr+/C0R7d2CzLi/dSB+/YQMMGsRwa9PJ/n1Ipf3FDV4pvlu4C/MZ41b6Cag2iWG2Dr9
4uSsPr0fzgMpcXIpn6rxpTgIkLWWZEPFPtGc4NNu/QSlJdrApBIXlsNc/JP4lnC6eVm6WDz7HcxR
aFmzYbY9hns2vJkfHP9Urb8VwGqpUea62kjWOFobxsxZqmSwBnaWAilgvUp5I37etULUAY74CoKl
r2WSksxbUhvB2t4h/PLEvukDv/EnyfgsbQltsCVSKoX6FGLTtZ+LSDNEkIt4vubHE9NGMHWKGQNP
73F45vWnGfbHvvCtRPvnS8BGn8tsJM8MOUFRo+4IKM7j1Y1+je3pi8KezFLnSzx1F0/0e/681bX6
eKmR2ml5DjA022CU4Y4Cm4kg7JBN8KRppqMjK45UpBjCUfUlcZtWagnOfjvWbamsl5KgtFN2grJh
FAF1aFthCMve/JArDP2eNLUC/YkSsGa1Jv+Vu0fJGg9bXqBc5BsioSqN7xUSBErC+GQzbsxHKTKN
Uq+EgdxEDBJ4zSP4ibQfXh+VqX4oamz9HYWZrI4ri88oMY444njWXzv7sL/w8NP2FNDR/zqZzndi
fXyldnqkz43L8A46v+giQc+4aT76OtJOjoM2WY7I+WRhiLaRfRxdpBusQ2XsTuSmPl2wYXLGvtwF
eUXe8bLhU647GgytyKnSAorf6optQxVUUZrmRJ122Q92Yl5yHsLE2xzPQ/OUkDpC/CKCyVslXyfq
hVnDqFXBkoa6ghwSXduQEpY19wwgVJ3HvKKLseIhbB5VOHav+27iFpBUkUxz9/Drwg7VLv4tQ1t9
448KNGaXnzSg+oCBBdVYhbhAOpSnVJ7q8m6ZF/qtv2KWlsdxI4gC0acIjZXtmYSgBJV8B0LwcE4U
3qidBYbbAJpBkh36c9O/oUCWLO7+j8ly5vz4EHHkt3sXq6Io2Rbx950/8QLJIULYkcZ5nTvkWzL8
eyppZ9zpYYdtZh64hSK7U3cdZQQ81qtAVJVcsFefj3mMkOxDLMTThhLozC55+MauusT7ZIAxjcRE
9cK4SosTCACVPj5UvePDa9Ij9E+HI6VeLS1iIydyrbZ9HNEGsyqDH8x5I6AHM+iWNrVUEMnHNBdO
0pyw8SrpXPB2JPsnF2jJPAviVfKwudstTwq9xBEQd1Pp+4XwKRu3qTfJNlrfKXoLYRs+x+f6k3EW
hBhe6tXqWEoxCDm/7XTMlIRpiPDwJDMrqmeB0Y2lny9gOMXucMJg1jmzPQSNbVrmO1K4d2kfoeaC
jF1efP1zrHXtGQqXkdpej6Bu5wNDo10swO4VCt/Dzy8ZWZcOoOwyULx3k7P2650OyAyhLGdiRl5N
gpzMPHbmAW1LLFa7pCWChs/BNbvwBKDXm7DwEAPgn5WNhxa8aGYw3hWO5EEFJWC7fF1tOKr0/PEW
4Iu6vCimwtIC0Ly2Qh787DhgYHlUJJsMiP57Jq/TNsjoV6MU/PBH6mpukcWRkmvQPvh3kErElB/G
Mvuk6NxKMbMgw632UiKu8yJOG5AahYU5MJrHQDdTd+EHuJwz9hxIA8R07a/wf2Ju5V2oGe1cwLly
gBBmui1RVgTRxHaoVWTDt70nesg2OgG4a1T0epsf9VDiwEBth7fS/4/JGZdSFafUzBwb74v1heYP
D+yHg73ls6ueJxgMf6NtTIi9nFmAwOwAa/ueQoSM80BXM1w2b4vW8u7HGcn28mzlkRr7ltltHURS
o2wTm+AEEaLkMFTzIPAuVGBR5SuyMLWKhTghKC+Z200a5UsdwtDuvQ3L9IwaW0/4RtfSwUYfZ+4k
fhEXW6fvmN7MbWito/0zh30xCvk20a4n7clfPSoETD0xIm2FKFuh6z9O6HUc8PNI4YGIH6PpW1YT
sbvT6N9bJ93bh3vpGeqVII7Zl29mKNOZFTaF+Dop/CbTNlo1iz3yvmvEWQ5CkKww9Jc2HFf9YPbZ
Hf7vYlwXIKoDcHyJeLpGugzkRfSZZ+mPuZeMPFcaTLRUp3bnp20o95QBKaABDzY9ogjd7H3vVIyQ
sR/tkjtfouHNjmyBBuBtALN9jP4ADIFM8r7eWaq0OTb3Xh3W4f0aY99xQka9iZU7PFKuz7kgiNhj
K+X+G8ocR25u9JiLvx29UhF9zEiGu0/xhlvp5dNqOUpzLbAE+CXMp5qWDe3X/7mDd1xoFzbI4cjw
mm9aDMdUIyFMhrorxrVvf3tRddxKsOMY3f8JunoxpdaazAoa1Q3PIB3jYmhDHSumYDj6RMTj2WpK
MPPJWxa9eME4WBy9phT87lrh7fimqUnlh9it0mD5WHxvpKY3D2V9Z8+wWqOm37m4mmqSBpG/4Oyt
Cgkw04e+pgDIMUMuyagjqj98M8JR3eK64P9Kft+dQ4QogLdJI/LL+S3ViMldC+HvC1zEn5GrJIB5
1+E8gtwNHP2005hqjGBiiX32DywdwXg7Q4wlBTFQat7on36KyPeazbEIsz7M85u41segndh02eh1
2hD9WL+4AHKJQVoscy6I2W4LZmymmt+DYiPNoJ3czMde+xmUxnZs/qH11lJyCsu323aWxEb10Igp
Xh9RhO7SI/1GhpQ7Agy8hShd3bANMKIT8ubRnRre77wBJZmj5b5BPTm4cz/27JiU40PDwPXEYJnH
+3bw8/q6J77MNpJvEL51Px1rGkCvZQ/7cDPFrqPe/sKOO49Jn8uvluPf0kWDIaKOOLKUXTV8Hqys
asDx8MiOs1sQmm+0azmE1ULbw3M8c4l6cajELko/PvR/lnSuvRBNlHPlCnnfCCR8UxtXA72975ic
t/4lDZOTghbsQbCfPmI335Nt3i2RomvES9/MLc0OwAbvjuh86h4mNuzkNmLSGtHS8UhL+ChMc97G
poyruljArIdTPJzxlQWBWDRYKoj1FdP9kKq3hxJwkhFkhAQUGDJzbzO2PQfYczK9zIsFbDebBwej
V0+sM3qyp8zYZlRiDQL519WOiRhhlRERC1v7Ubl0cBcK98CSf+LeF3t9yTf50Ff0afmxfY/87wNL
3Kl/VpWew0hStCcXqI797lmWtX2k1tR+zio+LVcfEUBwcUwQeLPW0RiD5TiINzt7xuzUYytdn3F1
C/ey8KtrfPIbf68TWKhgdho2NVB4SXA/yHxDs4b244tfg9GCgPuhfagt2jljkfgvZPKrEyiSKceH
OKteoSh5Su7rEase6ByNZYosuY8IcWDneCA6z3rFNaqsjxWHTE9PfETNvSccX7++lSzbeaspxdmw
2BNAfexPwjaQDIaSVqLqcFA6jYXoUAsE11UAepgNTuuUQt+cmrUKtgT55LDtUU/ZDkHHK+j19sJG
/wrci3CGROrxpLUZGO2Xj8itNE0wFkF/7r/ZTogEQzslXlIV33ALF024SK39j2UJPDaRpduz5md4
CUaDH20sxyqU6S6qLZKf3ZZ/L0ilrpVcPgYzIyU/190g/3zaqVS44uWf9nVqQek1ObxtmZH7esH+
fLjKXrKl7gIgbzizCrQ5Efxyi2ztU5OJLIgLBqw156S+qfbRJ0//G2p+nPyZ1g6HwYcif7G+My/v
sY+2W5tVGhUBU/XwWZNf/nW0dnKnJGA3slWSmKG0M9hGWNGazra67iN5uVw8bCKNhdHhak3jAUx7
kaL9GGI0BIyHImTlIlR5LZ5pafJcOaMCne3IeImGbfBq3uLgE8Bds59BYIz1BbzUDIDwi+5GRl78
LKldGRuO4kMvIbYnAKIB47fhPUILqEyTu7U8XYZWv+IfLiD+1cw4dZljQqqUfEgf25ThJJIeZp39
GpyGsm5F4kGrKtS9eihmpiCx1rfTWUcHfAn76mIcBi99N2Hj6o5agNkrz0V2snhxh5aWRTL+ELia
I1MOOtjNNrjPnEfbcw2Uv1jyOo6K0gM/IonB/4Q5yCzg6FJUpSFj4H00CNUzU5UepNa0GlTWEXaq
y//lzp8rY/r14BxbJ9wnmKRBWtPBCpv6HLCK9GXPeXaqLu5IMEROW4YZaISyGZ6EaUYd2NG+ALLN
+axJ+TdGikgjLxW/qgQBXz8hhGcqB9hhOb6enf64GVotrTY/UuFIW9uS6vsQWs+3H6oXidYTeFPo
5d4Ca3XgqItIYt09/5tJZlvfl/w+1ryatNtHxKBxpl+OFkV9e8GbbJfwM2B+g3+UbBdTVHGo4kL1
Nv3PNs3glkq/DYNGXoWViibJdvklxCg14y6++2zYOjCrAFMbMkQFnzYGzPY4bh1O15gpn591YrxY
QhK9Cq2eeRydc/AI9FKsRGP/gizHBvHjqZesegATxE8FYDpT/5kHXIBwR6P07vCvQGiuSaiyCPz5
X/1yMj7Ogyky8tF9O8MNrpi/UR/jgrlcJy9feT6MBKW4qxidT2o9UiknFHg2pQ+RjOjvU6Pp3btO
VuuCEYX1WIVFOkbKmbpmTSWd1zJhKeuZQh8uf9rLWtggx3BOigVneNOYTk2RdyNMJ3U3X+USPWss
/ISoq1kBnQXjK96JNjiS3vqmml54kY4twTT0Sj30yW61cZV9zempF8UstFpf+1gKYMUf++o7Wm9q
knJayLthbgQZsH+IUpvPXk1DE9Tp25JO+vyfFsqPreLfbDjqdZkzEL384sZ4OoLmFsnbn6t66wH1
EnnEp2+yJyI2yyx3AkkJVPL/uGn33LIvoDGy0wlJuRMcPcrMTVwne6rpEZGI6NMR7J88DI6yLSO7
e4F60Dez1fp5Am4g+hnT6gUW6VOf1PR2kOb70+bj6aWtjtshjW2ngE+v/liyOiXp3/josWF53QCH
AGDqKXLpoPRVx3QlB8JsK9gpD7/ZSKAkY5HGnrQjwhOz0YPp+baKj+gHS719I9H/ypwdGA9QitT4
uv1ijEC6O1vRaimoTcgZfzc69BcczK+Dph/hX8cP+y8zYXbtxDfVsMU6n2Kbxblj0w/PifbXOeSo
BD59bMMSjshiILEOB2MK6mUtMyCzbRj6EJGOJkqH9Px8+d9IeWsGxzUXwcBY7gHEAkAZTdk8dQwG
xhYiciBHOuy9XyLJgQwOjmmqfQyTcLeOAqv6q3tOoSgNSwmojKARCDiexFxwkw1oRRUvztKeZzU2
kub5Wx5yc9Jvl0Ox2jriHLoCG9hMhZQsAJH8C3VETo7KbheY2x+bzvj/Py4khcslfJJKTpLhd1ow
6K+BKOmyRtD1ilY4Im7DuDdNJivxtG6Mnvcp7Ka6e+/VbsnmQG7v2/6dlFtyKVNG6nwfvjClGEzc
qbtdSg51dM+Qed1/qE8Ts+/rsQouX/ieUo3yLED97mxyZQJGfPqAoaFo8QCGSXE1GjAl+aN60YEN
1tcWNnyK888qG0aDT1Wq26a7PeYXraAJb/SCsp4Mn+zaUS+GkkM+djJR9UtdP2mNNm9Ca0lybpra
DYUejWG/hDxfybv1eWjZ95tuUv/mrhf33gCk4PBfQVgrJt1lhKXEingv6o2yEmaxVq/R7Y5m8BLm
3gVKC28tUmspuzSGG6z6qfS+EaSnY1ntIlgkTKcSageTC4ubCqQDruLAY0KLWroR9TRgc39nR7Dx
cac+lbisqJ6PeN8dbtQrn6SUViVqyzKm0fKi6eJVC/Cfjj+N54uWYXDiP43/22EVWyUjTX/gNUsS
wZbzmljy2DTjgEBuBj7NvKAP61QN6e6pTwuvKdAe4c4NyiozzaCIL+2yAo9BN6Z/3xbfJMo7SAY9
iveSNXDJ/uCAiB7/6WDSbC3cXzCbDiq/o/QxZRIVtUMe/R0wSHAL1ZDU3ZHOol/JMsKMchkO03S2
g4qlClx7MM815COc38bb+bU8hkx2szDYGRXCeHi0q9jTubGufWPZMEpdGc9ZFd4eeNxSrNyBLjfH
Z/T4ZgPqm3Kk74PvhPWA0jWw/ombEqkZ+UT4DvgGMxm6ajAFrKe0thPW2pA4GkwpNZHX5nMLOqvR
/0G5OrSmUj8PTZ6EUaGHa5EzETBnJBg4ow1KakW9iEW5ZIGm70vlayeoD3lOLu/57nlUDax9IFP3
m6rpAwHmTkYjzh2M0x0zj3yfL7dVh5SrnbtYfdNrUX7mYaKMG7//ueSYondYgm8lWnBWpmhuF7U2
GbrBTe+mtSG518Ps3kHgltoLS4t0nSW60Gav96mCv9u2KRb9+xTKudatlurDu9s1RJz+8fUIFL+t
lAQadONqu45S/0kQ07ks2ABHck71HgSEymI9mJYaFFdDOadfi5kYzjKetRAMd1NEYfbNIFB0w1tA
8gI4TkxuWVA3b54Ehm3l4wLvauF/CKW2kcnf1ogY3EuV+MEyuPrvAfJUII4dkmnUXBSQU+xVN7Ew
7KsXhBLRnw2aM/tsIYV7Qyo8Xq3Vj+XrWG/ilx5CyQbRi7sVIZabV6aHda0yBp32WzEV0FZbi78u
6z92A1wc0VPvhdEnAq20YhPB5Zjwo3kmU2Rt15p8YvSkziCkQ7TJbpXAcCIcnCLSotUCSZM+Le3f
tlzfqNMjiqAFuEl7tdh2aySow9lCNAcAkUy7hGJO+dktZ/4fmRSh9rcVjCyvM3epQB0PjP3tOP5a
TSzFDDg6Kg6nd60d4HyHS1NNuM3eNRMdlU3ueTtQ7ToE6E7LhtXxiYfdl3llAWOYw9tckpxk0mCL
gt1KFL8fG3faWtVBpw0yL7DoZdOayNDmwQ0naeGd2HrKBHFmgFGVFiHb96cS7uDhVP7W9qlZk1WE
2QzPZrYucaOSmpGGOmrAT65gPJWSxhWxVF8eORZVwL5cUfo+xPq+D8fnRvsV2LI5Q6aU42aXAV2d
OqiVom1cCZgSLGYe/MhM4+0/6xyp/plvMXH3BcQGH/YxGO00mtsKsN8+J2QXH4SdjcwR1Pg4QUWZ
eyNzB0H04SSzboHpfMgqTApBbk1ivTN1/I3VAjp/mtnbixZ91tbpjhr8qcWp2/zUsomTTv/pggAz
Bmw7cEnO9t8gYkn5vkIASee4Yw5J25Ju6oXtowUo7Kq2FzHXtnxGm3BaAPotbWQuz2lBghEWwysp
8kr6ZFcn0OcEuQng0BOUhTUt4qo5IfNVNzzgXpSwllgQ/hbr5QT1PRlegQNj+hmx1BVy5kZuMApa
rallt5Ml/rxY2fnkOE1gJyAvJhwMdLiHghZ3ligXIoWJi7hwuPvNi28hrDpoaQcw/ITjZoW7XC5q
pbwpCAnZ2/h+aGOHN/IKdOizDnFcntPyR4qG7Bq7LTwFWWrLg25usfpdeTilIeduOH/jEK2eBZXK
+DCWr4/Ala6Uu7NeUckC8cpkAQOdSaPdKuNSFQUSPzSxVosfz6vvUQKX3Q55pVUL7g54wAuN02ER
FDN8uQs017NRw1A6Bix3Shvf77jQHgyhl8FBfp9jITSXQPQVu9+CUiYzYafbXBkufgxB/XDXBtK1
hf93v2A5wNqk/I3xLttayaBIGnyyLIt7HXBhQ4uLgUdaIZAul+SysU1AmlE5m+5knDExmLAijB7G
n3iiPXJEViSz2uaxhoVIY+enx//LhUe4FBEP8xcd9Wrbgi/au0iBiJMUIYM0/AQ75bRsijxTcBiW
GbBBvfdB0GN8g1/kCQLkUxbxrt3bQyN+ViZadf5BMIGK7hDWMrq/nOgQeiabiJ4/y71sg9HKElXD
K97qZvZSJ1TVP1H/Bj7/2vUylKmlXZPBocU83jYhOTsmzTA9d/1JmK/3gBAyCRZl7PCYkbxBjGCj
OovgFVEta9nr1tmUQAs2WFFBm60XMvv7w05T/Ecd8LSSCJTYoCkGeSkZ+cJLCCW0ARsmpFjCDNDz
V6eHm6v2dBqpQP+QNd8EWi4RTZoC6igZQhl1U5B/qQQlAznU8MlqyoDU95f3T9p9FdvT5fFULDfv
bi2ISDhNqg2ZpqNhiSm/+YbK2zUqUc/lM/hpv3hQNbPd1QJDUUidSVX4kAbMB5o9HvOmfyZpm+X+
1OghmaLaBP2VXC0pKj4XU7hapBY5EHXHK8+V6Cjt/24iXjck4mRK7YvFsAHcClS4g+3jyh2WbOKh
o/o3Fx9twY1YT+MtIt/DZLqWbHz1yY27UlmQD+Bd+VuEwIezhjvmXrAElG3PnSFplICK7j790XZr
KiE5A8TAUwbfJUdLNK6cJvNZXPm/6nr9fT290Pg3iL3Y4r10RtxGtGeERnvG5213CsIIV19bpK1Y
/2sb4a3tonKN83sqXWdxts8dWzc+VXQE0htBJaqcmt5wUgA3vSuF418haDKOm8li7FoZRetUQ1rI
OgJxBr5fMHUiU7gPlKGWCdtZo0CxEce71Pt9kUJGQz+7EQKS23O3DH9zE/61CnNcNHXjfOzaUVRK
jOsYG4GkjvStZ2WoiJ84quTBF3Y1B9TYpxLNgYeHJCqarHldIVOLF1oa2mg1hP643yXPBVOIs2Bl
VNPWzfnedQDdoadrI6Adrb2Hy4u7G/Wy+4L7itmybW+ULOeIgiTvvCfvaiqIa0f3ibRtWjtgpso3
16lTHSZneWBpRWlOyi81e7mmoANkhdVYuB6yGUxdS8+83JgON2YIhsWylNhzrX5kpi3RRe/Elzqa
jIhwIPfL20xnofsBfA23W246H+IbN3fZ/4PDQaX327OuqyObEJkuSGR/f0UtiDtDIXRT7KW34bg4
YwSvXY4rTCKaLWSSOVQQMjsS/Y/+PzUtXhTsvlkcrPJrOb/2U6enDKbBK/fRUME3rm2v97aG1kEo
Zsj70OiT4fCbvH1SJZOgMJd3gBKLycImX0Zi/QouPPwuWhrsKJDNi/pOMjIGttkDvEGDz8ILLcNF
1E+sJB3Q674hsfdpuu6HIbedJV+NnoVjN5K6A2AXe/Ygj321wjIvmA04/i8D2u76I5STferfIzaN
qnU4PeGcRU/u5qs+W6pBNvaEnegtI/5YUw7ukG+BpMzhv33tuFmLGZKDXm1ZEEW3f16+nJj6pykx
Cr43PMtMXgBI40iSlEoP0ApUfjBq8Ho0lzCQH/AXpkZFnjdo4L2J8gdusZq8qekDpG77YOERGhoy
8U/oC6gBXksOiMJS6pXg3U7zjMc8KZjX1NlBOgbB+s4uIUGHzTrq+hGWKlWXfBjygQmmZBWHEx7U
UJCqCT5iGbyH43JCtksIO0I3bXVog36leUshDZmgkTv3m4TfNH0xbsF4sCVCQJEvHc883aZiNQYX
ciaYqu2sdbPwMvoasbjar3p8Se1W6APz3tpt+RTuMLzgkpvR4UVPQ8iGe/6a+Y6/SmuJogmIeNSL
38qHbkcwrNk13Wqd9lZbJpHxZs5u4hKYyUDhKBOcMH7+WduCPQ8gnGrq5u80OeKAN43LoX67bSJ9
t2f4MpdVDEEz96dc7016fQTMc+UYbJiWH6BmScyGGpoSlwCtF4rNbiYIl5EKLWAOKjTgWjwPawNg
xXU4JZK50s4aQ/MvNE5211QBrsifeYdZoXzAp8Qy16UG6yDU8EfYwJ+FpEja95Lxxk36IXNSjXPB
pDmuWViauFAbJXQbjpEsYQlt0zvW6exXR5MV2IOKwWi0jgJI+gXWs56z9mFG8gjOttKUzG6HBJed
7jeev+dHL9wCXYSRBNC6rOvF1oQZqZsHyNzyhiydd+901yX5MBdxnUs/qjqo0A0rxWeoi6P30uX2
5ogyairgLd4Ot7X62ZvBzvXg9fwcUpdfEH/wj7mRBzOW3VW9I6VQ8iUVWe8UyfukZunpflbciJdO
mwW2TWUFmkNSnUp3j5kIRm7aLpmA6hC01gSJXh8PVsb9UrAITcASGijnSUuDN7XTkc/P6kmWlJDk
ylarVnQAhVXzoG52V/TO3VCh5OXwr20NK0UxlwS7ywBRC5Cg6zsEhlEX6NKoNdqky60oIWs2C60U
3R5zIzMflp5nRDfyw/37/CHtX6I34KhFv9sHaiz2nz1iCJ7tAiFgQndcLZgXNfoncSDIOVyP6SS2
OeAV4EF7Dlp7SuBF1PIOid+tPexHbCjdXJ4nfIpXwWCaT3vpS4DaOEIadf7eXeRnqKTwNWGGqYUU
1Spf9m3MbseCSN21aZCW3TBBpGH8YAlEhh9L084Vjea/JISBmOT0nl6ooaGPj9N0SezNpyNdBqHe
WQawLyz0YVlSPH1kJ0usDOI9aosBGq6/jvl+uo/NSkwt+CJ+3QBlS+SKXWCIiQS0uuETQJKBWzBK
c5VAWCJYvejVpAuKr9SC1R9hcdhS+CPgzTtUQE99MWhMOCH66nxpYn8DfTuFSs9h6HdID4n3nGb1
KI+eqRZtDe/WtqNOBo+u4rFp81Os5Jpd6DYrMK2EyBdK+ayqGld4JQTw36omisUPoeBhz6P/5/by
VwMTgY9FO3wai+vCdLczt22L0xemtJ49CL8Oiq6/3ZLL7wxS9sx4vfJPkibTANi6ERpNo52ikgqV
lJTYPS1lXseoH5kahdkekg4A3jJzEUCDRfvX3/tD8sWe1YuhpMxz28VPz+UKxH7wy9V9j5e25A46
hDA1N9ruqtlmu0ZdseONpcE+gEkSPEul97CDw7r7rfI4ixn4qEJJ0vIvyrTxC/oUyHib7Ot7tRio
vg17wN8NQ3pd01e/QvxI2QxTaJHYe5T2trastsC/hvB/m7HPA+u471NV7XywXmXeJsPBtoZtTCKa
caHMWqNuKwM8PYuoNYTPy/L5GM/QgEQ9pjQLB5B52TlK6rJPn0b+0aKP4NQTdSshGlmSjH5soCXG
f8ZRv8I9FEE9BVsiz0MQDKSq1N/OmqZ1StmDRFohFldnCDQPrTY8AlivO4jkhXgwBAuqFB+L8X4t
pY621VDnh0hVfIt9dcUfsdlgC0GCBixDsBJHxS5/sp1A7qJLDZfH2ubwNSvwMXB59/4kLOnoDelI
P4znXwnXobPIsUVJdJvkZvZ94kE3IYB5M4slFKqLqxC0LFvJiW1LgCNoLn2G+MXvJOQjW1AS1KUs
LJeCoyTDBkzA0dbGWWQTZAfT1LS/I1dH8Zlqxx3+sG/3iXWZ0vgs9igtNowyA/SwIhLo8BU1j3aq
F6g0MDWQ/f7br/6Q92W+S5RMKZqyw8mOJx9IBjYev+NQnc4q6FOya9e8l223/+q0TF/mPhSPhvOg
g8yIXK0x5KUvZabHr8Orl+Mu9XVsgPpHbhs9sQ+nNK/BeGLgL/vGGQ1xLAaydWv7xsZ5WFO9E4Qb
ImUlo8a67gy3NUUHuP+HGIlsdqzxqiCrH6fdXOW96zHqVb5vQMBp1lKsQOpYwRiahl3/3pgnW7oH
QFJLWNYviM0sVCnnUF4BkzpiG1/bvBJxQIgNSSF4olDRDgXs8J17FXLFv4++o70xEjriA7U3M26b
4Jno6P/AecI9I7B6PHo+CEZhyPLL/85rmR66jDkKGNy+dVu9BGFtLcrwlBiXH+YW/13QYFF6ROTc
DRNIZhG1zeMeKNm13765cztHaBJVGrwSOiJaPLkIepgWTGbbR9DcYd+vi2R3KzMyq0JlY5750TYB
47PFzWC2NabTt94286D+2IRon8EaCSra9PTTkAvUb1GY4fQ8ZS7fNvSMFqeVIwQzje7HRRBT4YVK
LSzRBGBWvkJ5uVzIFpgHbaJ7ysJU+KLeDyA4JSHbwJ13ih+/4sd2NJ7TyDet9olD/7Ne8unYDWAd
erfyv7IVFjfqBbz/KYnsuGt5cHOHrpthBtBvX73A+yizpTvuNYaeRnyMTifFRdcsS0imcdOXquFq
WG8CpAGi4cfMzBYchUX2pVLUs3mp7r8PGsHrIIFCwSeWJL2m7rKVj2GkFABx8KiAlixVkIOlKhVM
1PNb3WKps4r88OnfSs/oIkK2OGYQA6F31i5Jh5REdaVi6PJ3bB07RQYWdxYTSHZcPjslEdG4H6Wt
DVgKcVSqaf6ltbZSsij9r6u9mSWYMisdbqdP3TOSL7To0O2jNnigd9ZqPGRtR8Qc2cxfQXbc6rB7
29iT9lQD0NcJ4V+JIGnRxu3gUtgz74fVJcaP7pFKeuFem0snGVGY9+nT/Woemav6CzCv6fQIq+Jo
RKAHJEuTZlTslls6hHu0U50v2qGmp5MV7l77W2k5d4cScoZ8dtiKL2etiQK1TFD62syTncba59Hw
3PTHOZ08e7/VOPypQVgV44Di0HvXn89MMwbgD1YnjoOu/l+X1Vu4fThxNiOOEJv63KbiPA5PWFt2
1zsXeNony/unkiGbCka278w5Rx0uSllWm6wct1LW6DE1FSYeuA1KBk1wzIkL0XKZwZSOWA0DXm12
fn/mXje1hMCbRMJ5uDKN5jmOglL3nE1PbqkugRiNo9JA3TYiSjT+yD+Jrj8D1ILJoOFj0l0vfFTq
TT0Pyfl00XZm1gTDDfWsDvo9qBQjo5S8lyJTDO9Y7BcrybkRUmYcxBAE9Kkl7AUDCM2crL298MZp
URo5YitkRRIQRMb6y7GfJ8Sn4LbbkZuJqKROZaagCMlCMZ316cG9xV/xsiwXPdkbFk5uCxdXi+Zd
WccrRASz+hhgDU4b7J9D8zDwbN7UjYm32+vPIMMUMuyYklAx80aJYFe/6AFRjCYL1OZ/+JPf2omy
JfhiwFV2HJoy2JKyBSVQBHZdHjuftfbV5YJkOZqb8qJI8Xmznv35RDo26Uq54rqOyJ2h929xHJ+o
bIupX/xHQdZ3ggFULVABuiCRlPVpUetH2COmU4KVlGBnXsq4A/wIikyHKz+xQqvoQfhw3SyAultg
2IBtgdvTQ5cfaXOMVLuyUXfFPiZS8P0U3PKx3wk6BqWB5Kw8HmAaAs9KRd6+bsZrPjej9kr1MJuy
jj5sUpNz2Wm9Vp2YiPRrUZGtMcTjwALVvGwr7VdpKhG0T/JYdnQN5F2ZaEwf6siQrtqky8qsYWSD
DSE08ADvcwD0Mt8GSmmvoriaLYC8WrlD1GXjAOo0OAwMzPFZ1o8PyzIaurCoQNRpjHvZ9QwEunmW
Ugwkfg3EsBhAnGBbf6CFlDUIBzKCtnHEuYSKFbOvp79cUWU9zNdGJYK+M+kXJOpxQa+gdXA8Pc6Q
wmE8rCYt1YNGt7dIJ0yTBMwwGblmFrN4fJbMtxRxOT8kL0Jx8mm5vMD5A4lHyUNgJEBecwJAuNCP
NGtYuAtIQ/WfxDQw2r7Gh6LI5Xz4dcV1AuCmXGxpY2szcUwxOpBkWqMmlgbbXMJwrmntXZDw+VwQ
jQxg2RQ1/gM3T3hte3xq8QQ3qtpA2RQragIHqB33ZlXDRL3UXMF3FavJrLYWDRr2m5v3B3anpVKT
S9kKoF8zgbZnuTs1N1F6hZMedbBOzCCqF624D/dh46QEpWEawuFc7MrFpbxDc4Ahc90iajonrYtI
rlH6Hlveu/bbaZnc8NGFzMeRXwEPgEYNqggedIrRfrOTKscx0hbNsi6Wtdp/4GsWPzWy7WyA8om5
wew7LvLkejkLPyJQeQF3Wy3ysZJnCYJCI0yeBiGUH/00ftG9gw84onI5Y7mmDYgtN9bT2s+dqy70
MxwqhuFzADtmp5Jmgrsbtj1/BJXobvSR5YCA24/Q7jqHFmPMFYDkL2tl5Ma/d35e4C+AS2XMRGyU
KoPhFU5o3fKg0z9QjZYaTycZR5zkRp7vL4W9ubek7d6/iQbtaXPOEzax3R2R33lGzk5cQaXttT9t
eOTc3/4h4bVxuv3YpC0G9s1MywOu+266KDT4CffJi4mcf7D/NXeyv3VPMLqEejyK3FFWq6r4KBP7
R3NQ5qQdeOfZTQIoN/ucFiKzUTvlTpAqLzHTq11ukvffDMD4u6ADKeWwbpGQMxhIGAzb/TKdyJu5
W/H/H1yz3QoDg6Y9UI4quh1m7b00l0zZ0QKKjm+qtwvmOHVe77WwEVSwonqtiXSHdK+aiw3fHkh+
RoogNIhXROUY/emwld799mIsuyVAASUdGsi1IvPDdBDbg5PCOFK7sETNRD9drBHmX8uibHzxe+8j
GTxjf7nlXVqtMY89PKzv+TNnDEJik7xYGRLNoFF1PVI1IWHpuL5Q/68sIwzkdzZDxsRiwgnYP8dd
XJ81jFHdj93yzCc1caraQUQuP+CgyGxHVgz9Fr8e0rQ8ViFbIbYXdfLutGtn3CAmVMO1ghfWs4xA
LnByHRn8qIh36hy7jS4cIYpb2Bk3UZlyN5du7l1gRAJn1b2usNB0J/DBNlKowLXWnHxu7jMoJivK
d12S7R8hmROVjuXDB4ltxeo0xTlYzdz53zTviRzpC9FlZm2g3+SB/Di0aGVqrT/a6KrNlQRL2JUF
hez5A+sb/1GWk6SXip2zMblXpkoSEGxCSkdQsNvSdHYHTnKt7j49BnGB5KNWpRYIzFwH/zyTPVaL
2AWsR20mxu/b/OvUkhyQD67Dkfibgyj/bzW0Uf0bY8KZkUI6wH6y3CKGUh5uQtPaHCuOdFeBPWSY
P51GdyyMK3uGXAXdEu8rosTmB9DqP2GHcr5w63KMl8gpAYWZLlMdSCzuZhvgPMeVtNfdxgmBeeoe
atAmUTPTw4YoEG3MwTlSpITSLk78fcteynijgSfS3PjJCfX8xynvQolRlXZHN4Ko6NHAjq5LLr9E
0hqbB1A/mmpO/v1V30WXZ8+yXBnyEHtrDcEehpT9THTrCJQBR/IBvaIHBgxbLTteEwdOnbdwIi/g
Kd46lE3HqrKjUDxKobxn4QgUuXpnaruj/kF2d/tcYgsMAqbPw8WPNDAVNcJI3b8R+7edUK+6fkvx
G1+IDnfx3a7zGgsb1DYUjDWbDwUYMzGUSZ7EZQ89rK269HLOlhtsziMCAQGXSFHx5XSw1wzKLN/Q
f2nZayhFucH+p58Gy5zgYpmuH+7DhklrUf+IZWYJocgFf+8OE6QdF5Ci7Bpc7FNnq9BcO0qV2V3d
wjOpMjdBAyCP83Np3qa1kSwbv5Lrzr8IJyoSeoDVQwRzEEc6NUGYaW/Ossitjj4/DeLlq72v+kUq
kwpjsXBeSuXfexblSKeFHsKYolOWPv7z46D4TlmbiQnleFZa+EXhFsrIY81xYPhK9QrtJOtyaeIG
yiAEN4nFIxjVzdc38UJfn3kpKYDDRL806qj5ungYGgOVaunTgxbk/3tImtcik8TSm4IcLPhdQWOi
fQouqnEl7l/qT1XZHJeEZqF2iKuRS44GI/c5NUh3e3ROLHDfFt1cfGS04wGavRrP1DwR9my3ZzRb
6SDAoV87a9JGjoGraph6yRjEHgBh2ocWtpYAYleKFFGM2xrNlgnOY89VZRgqi5yMnVAOIy1aC714
KbVlzkEHyA3R7Ab78k7OfoB2UCuHosdO90cgcTlu/cj9YNgbADe+WZSR72g2p0iwYFGqnr81Yatu
KMzRSksrnEzvW9JzxG5zdE1jKgEWvBQVqgBKpY6cJcaEvOOi2dcaK6yKYSndBemj2NBg6Xphytoi
FABcLtEPU03jeGVhm1Pw9RXwpg8hNUstOj/+aUgahGU5bQ9XhCQvDZJUn4ThiRS4JRkhs98mGTid
Pnvzbg2l5SEiJlqMdI6qQelfKfb/BB+d/qsT5byVBUjOHcqQCAhpuNVvqh6dCtVERj5pGz0g0ZUd
v7EfdqdBD2fHqMOLj9aZuVuxyH0WzX2irw/Lw3m+S1XXP+YYubid1kfG3CyJeM5VqItmyeMYPc1C
DM9auWfGJZAnlJEDjZhEdzwSEEWXVnDsI5C+DqGLkVOx5XAiSkv+JMB485mbwtzQz5zdUivOvbFj
cepReah5ZpmuIWjSR+7UJ6GmITgblTP3CYbKy22LyNTRWfm5gmfCoNBowIfMKxN0R/f2nFo1HBeX
mhEMPxNWw/P6gIB0HvAPHsGKRAyRuIM6rZ0n4uRXQqKZwRhxSkGD5cj3H2M+BPXdJU8lWDCpjaCP
K1ad41N5Ptg6tqztZjJ/86psTl7a8S59pZT3k5cYw/uxNUu1TSR01KRqF+vEYazZU2ehu9ggHa/b
I4YRCFvi1aEHUFPW0dT6zrkU5kSQwZBplaACy+qXdCAp7hJxL0ZlWLyzSgsemyDF1rlWZIHmqDso
Q8zXtnrgYu0gUR8TcMk78hZchXCjL5BhAzUpZFlC7s36C5mYVDrz/w3P30MxJs56f+lWFnm59oqd
lwNxR6yx+bbUu2TJjCLgZBM0PNyC0zF5tM8ldDM3LAmd+4zyDczYIuM115ZLwyOqkZXqyYIjLP3X
FNmq4F/1RbRratBVlNzGZzsQjZjLte+Nt+XxcI2DEfzjgx/xPuceRwEHfcEOpnembdu12yInqwGy
IQEPfgFACIKQTBu04c0gAFAUHiYn7DMn4bL4dMXE1Qs1DiIxNTYFOH8vQFDI39KYL/ShCXYaHrJJ
OBouCArtt+K4OwHd+JZPWOPc45yt9d14nOTEZWJhrTvBVOF+WEwxd1sEQ9+zaZjeWdcr7EfSV3iE
sLDRyzyHQUdplKpUdtFZWo+f4x6SVb8niFJMCgq0Q4kUNF9gY6d/4WOH27ZYJG6B1t14tBpTyUs1
oJin2q4bU3KyqPKhu26ru9qX530u3z7dd9M97lap2BUPkZ2HvT8C4xJSrty2DjGbREHlNdH4Xdp9
BidfJ0ZsiL/jnPHEDPS5peQ9PsxxC7hlfNUZIk7G4lHIXLMvRY77n2SfM53IBru4E8wMRpUzbau9
ylYyi4vMY4dNVtXrDlQyDh8IfXGWYnei/rBV6vWcivuFzJv3b25NBI6NZGqNUPL2hXWrGpWvv2Ed
Fwm7DvfHTabmAU6wKUJDos+JpMugGiy8pcsj8qcr4fZs8ojegzkeDKSv9p/J43X1nbZbCmjcpvkX
kG0yWDTqp6A40MoQfy5zjcNIMCY0gLgnB2mWkGasNyO+RofeRnIXUy2S1VU93Uq9IE4lf5PjL5sK
WJWciqW7WqGTn9yx6vRBYJDJho2iXfPxxbavf73lrfM4EZdxLx36MzNPHuAyFmS72gRM7qpMno3P
1Fb5nXBH7f6kfiIQhmY2Q5bkH6uPEKSXjFrZOf46MTy8g/fY2x3ubF7wLHa5+OWnVFQccv8PRGro
088PzXXBCXnrLO4G4JnSW5AH54DzBtNGOA5yzul2mVWNZeiPhgr83T5HaIpyX7fpPbvmrLrjyrRp
hKiYKccsiTrYSJNp+cebfrCE8s+InBbNDPtkjzXlG2pV0zXAfDxRkYR/0c0wgFvQU1nrOYAxBFlp
kjnPpEWC/CjjVL8zZlXBFsjWJGirYHirZM2uy1YgXAcR7r1DuKY5UIhTx+kWeKf0nHKj0cf2ynRR
sHwgNpkNaeMmuSq2s8aRRlia3TAKz4jRT8cnHJfN7+5rwFxW70hQJxT1sJ8FnBg2aeOVVKVrjL1r
1dlkEY6Npe3lscBxrmE5jFgEV6tmQVW5MIH+2WPtyElCPZ02PlK/mP3nU9rT9kjG5zcELML1NUJ6
R/QpfPwvYY2Z/PZM7icCOLjLONhsS5gwcHzv9aFbGIHEuDsrWWXXCeORCt6a4RMsxpPfZObhej8I
itvc6v/xr2WzVsw9btx1Rmuzswg1X4ZcSbdPA/McwuWjYtAsvy/qJneUUMJIBQe+pdg97+czuK+E
XBSydZDpzD8L//UnDdVOUyPlnjFUteT7hSj1nHahXeOZgv51WKOALAr2AbEGjr16zMp1OQLP3ZoI
7sgu8IcF7LBPRnu/GVTUFO/8ukn0azT/h8HGBsXHdV+gQ+0G9XC77+Yp/WLNjRPEvGJhNhapfnm9
VmdQmDzROewQZMmN6EqHftQGncNzKuT6mWZP4nrlCszRh02ILOcbF3GGS+PH9HmVckk62IBadsdH
t5BXeMhm+VkIqatHNnL2KXOQxR0x2t3Sge/0V0TugrRDVjQZfnTzaTz3ZdvpX7TMdTf3NW1mFoGz
uol5gGu3/8Y416kX08071HuCyhIkn8PuxNssiyeKPBIJJ7A4G+41UUConcjV3tXPNRbZjHEOm3Py
New4l2Q6u2Y4gqK2kd1SG1XKLuJF6HVHPKcRBpKGGUCCcptb7m1RiQorDpBSxgnaFWtTFzF9BKPU
Hlu2zchGf5/pXgHNSbwoZuTeMFAQ2T5L5uc1KqAV6A149Ei1zf1N6mqSL9MXyau4Z36npbHhwdqd
fguZYjYki+chZqQc8a8s3C90i7pOhx3yMpLVQeNRbQ66Jg11s+XwS6fxEOJbqovBmzToQ+ErR+lO
oWxqYCyqSLGBv21LMlzZLymdmTb2N3RjN9sliZrUDBCdF+Suf5n9cNKWyKVOGvytpWhKuO2QA10d
6Dez14X1RKr8vjtJ4PnzwnxspCVT7OVSoWRL514P+TR/wXVFMOwA8BfA2gqoBomTNXElToLjOdyO
rbLiRfxJjkuoMvsnbMCw9gZzSCvuvqluXixofShE0/PyAAjABXk44u6RomyJgHIKvTRiUzkYgBZY
E9i/qzjTtsCFx9NnHPs7fVWEgMAHXa/TjZQQcQbwSLy2PmcLUpCgsYFKduKCN8XmaOt+yXAZMvV9
/4GMCIpZwmZy1yMyUUhw4E/QaOZo6NGycqjxdqhS7/OzqXSSz7/x020kbaQYYikhIl1wqPw3gcJb
COXs1xVx0NAhwZ2cUIXNp/PaqIoaa3seKjrMsiuzC8v5Yn9+dAxFQmMJuYUegDTe8viXQlv0cpLS
QhZWbIB0r3Vy8OwWYq7x8SZSqfA/5qygp0YQAjM9aE49NW8S0kIbMD+E2597PiG4/4SoT71gv3IZ
8GZ7g75Tge9ADRlaSOEf+EdlAoMfniE3r9ZfiMBFZByh0WRYnXGz46Uz0/ID4bO4+BV2ErgRr51L
ggRwzcB4ubZOBSHRTsvhNJFtsxbyYUC2Xh++r0gwQqE0zsxHJqeHh7HricHIwLy03qSNXuHhVSp5
s27Z4AGWCXoAFETpOf8atSrkj2BXIA0nuFlanf6Ln6Zso+nMFbdOiTQAzJMKgayTK+NhhjOm1X7u
rvgxkCsiutgRf4zpFKvSiJ+7PFLMmdeNMdq1hmy7asiz6oA8uMyAbyRq9YW+uesg7187mDwQ6oSy
o3IwQn+2beQ0lmJZZGYT8ZjJvnmJRsV/PUNQ7YyZOc4sXvKmZtWUZyRSz/0YaJojvRpDlQOF4fUr
FwQdS5nIg5LFSwGbvFbRNdxIibZTrjV4EOZhT8wb7FkA7ih3567AU2JLb0DjDPhpL8BNRkJHQXzM
ZV+YPGzXKA5+Ewgyv/llYzYh8EIPSq57Fu3ufYX36ZnfWw0sM1w2vUwMuHPoCKPZFSm2zHwAtwgK
wVeQfVuQnFTdUT8A0V34A22jZOPxX5L8NIbUNm0Hg3LSOjUdcV31pCL9bIvcK25eoSce+9THvbGG
d8B6wBWKlPzK2c1Hyvm1q/eJyyuZiQ1OAQ84ruHiX4jhSnNGny7RDLqX8p5znn26JHL+W4GGR7SB
Ql3flRWztEzsRpNKmcCLaWe9kOQltCFBVmQNPZGufEa6+lUblDEBs/uK73FOEAL1rUXRlpQobGlu
xXez1KJxT1w/ppmnKdcnZkTgv1AwJjl6Tf4FU0EdZleovmJz88ciDNCVQZ/U1Ba7MFlL6+07Xeo+
qqtxyXwFWtjTw69pTRcIXLOKV2DD2zfzuiGZqAY925qfSeAy+bOX+6jhGqVaiLhWlc8Im0ubwwEA
n9pjgRrpyIn/5mecfeqK9Z5w3ZYwUMCSBqG1bfnqH8oeA4261TjceLUV2YjJbGOfd/Zc91ZPocoS
4YFPN48w96Y0q7GYtc5gCjRHWUZBvzARx+mAgtQ1bWiC2hpN6Oj0z3TLLrbGfSe1v30Xv7tPkohj
60MbN6xKKvKe0rMZnwDo97nWuWp0LUBm8y6UWdNN1iQVgaTVef1kU/OoyS7c1CAyJLtQ0NPt80qV
CcGj7yntDWRMmnqkWjiA1uVCLnij8+64qaC6lvlQFtzW9bn7A9+jFbe5BhXnGXOmmCch6iyqF010
T3ZPwRyLTBbBfAR1f9l/+5wajLvT2ljvEWNXmNrFpOh6wvPNc+WI7qY+fGrViqJ1RoPvNZb2Ko5F
g2vZ9I4C46GG0pz2lvIf5DPHAXlnFE4/eRlmvoDIOditzFrKOqopvI3oZ49VI5kBV+re+IyKJOD+
k6aK2FhMXB/PeTkjtApIfKYd/GizI+SYrNWvz5conqRvV9W9UJBs7Nh7hQXNX4eGsOIGC131NY+o
yR/w55uZmI+w8mTgoQNoUD7Rq3GP5P+QIqMzD49kyDConRHOU0kyLEJS9/r2PE/t5Wo//fMsgiFG
AAAFuMdsugitNbiptaN6EqhrAZAEvjVuFMxY3pHm4+EdUdQ7LfULwIxNfsY6kKMRnXNDyCecmmxl
hEwi4nNJQV5ZTdFjPrFySCjSHftvQ0XirgfoDeii5gXaWSgJ4Od1hYN6Um77BRGSgWiTvjIL324r
ccJlAXCi4yVVS2SYJQipeFbVgX3G243FgyNXB+/lUK3XdBH6MuSNmJZCUyllODbguGpBgijeNsKC
8nhgIzZPhC1t2qx2LQctzl4jwtuZQbH6kp0j7jGtez4ddODbbMA9R72CulUkdivpWGjgvorgP0Os
x1g0SFUZZoNmeVEQJzv/WYy4A0Ev7mszbi55uUalBTBKcY0GABAAAJp08rYe+aqSFnGYiaaF42GC
mmdXM7DAnzf5rofXNP62dYgoqJm/JGKWf8nYypE2ZBIKl9knd+6sHSInmMr/zvyVaaFwhwxyaU73
vEUlfXMN8fLnsbyJiwY5RTFXPrfelIPHuDx1DfK1++fqNjSbK2g2WN/7iU3iXZOumT/DcvY1czey
Tqa+Myzs4RWwoih/ISZrGqgiDrmRixbUyqVX9l+UtBtlpp3l5Dc5VWg/r8dWToskt0ktoQbn8p83
XR2w8HIE/r/u7bKOzYaG6EQBpQRdCAC3evNFKsSekS/sd27KXDoMMrii5gBOpQbwXa6EPwuIDBtt
1VJX7Hc0lcmphoQwbzbZy+aN0wuKq4J5BXsuQoAIpYOOT5uDE2TSBdoQTAP0Z/8tchQPX4y3ZJr9
f1fyAgZkQyUA+vj1/BzReDyHnDGfoLVBKE33pJ1dIVp/p6a4L/54DnXNkpCxfL+9PtMVwpRWq7hM
YJSLuPmru48Q7VsEbUu4At6AnqtjPSuZV60uzAXlY1uF3woWkk/1+MPKkNmYJ7cnLG10G/IW+07O
z/DGByJfbKaC0CPBfDSAJloMCrFNbufI5Wgp42OQwCbv2gaUgcEAgO29j9C/jenyACQIhgZ+8fCa
rsLdC7Ywiv0nZutLiPoM3XjMXzWqsh4qk/dXaVw9NFf1AuCH6ai1BsPvdabdfw933bNpatpBZubY
oEQ17kwH42tSXIo5z68IPNYOry/JLoiHcKVrp2rqGrNp3+03wXw4rJ4ppoKvCBa7JMWNz0XMhbfh
YeBbAUJCiyMlSVVWR74fNZpeQqU34IbgZty74/w9Fa2OXJNlCln3PuWHmjyhAHwlkuzqPqxwAfZV
0EexsdPJT9/NhRQwVr7CnfjAwU8LacYWjxK6B5OOnyF33zcwJM2WvanSt1MadmtPXCutkTlB9UAb
7+x2jhI4ryvkLQLVS2c6IhqGaWJ34JJ0Y/3iIlnMRhcKr9qWHo+Eb6BRE09yAqgZjasdBsU0HNJ4
o47wIpZVi3bxiHRVILSfxf3smJkMOlB9PGA1tFxqAG8xfA/clAhvq/N+NTxvp/9dSjjtR6XK7Pio
kCk4sqwpezw/o9PLlnPf03dxeq9Bmtn8J+/aArfwCBwcrTUpBitWX7igypDUvEFEtjfMMgOShAZI
FqNXr+GJSeIwmxf5eTnRMDwRWAul2lbiu46CFURYMQVWcHdCs/Fzrv2bJ8nUIwYKGgK7ZyCGR9EQ
t0OJLh+99vdcXVwibUYDsCwS0/Xyb6hiMg1iuCwrFpucvxfF8dY9N6y8psylP3IazttJ6gv4CTRN
3qyEE2FPvtuhi6XCTU1wSPP/di6K7JLM/3VkQ/A+PxsN5DKhyTkvgnc4XLTDY6LY63bGb0NfO6gL
qEluO3hRWZHAyo/mjRiFAIq4jSoHMKIfOITBkOvXZImOmdbShq/OeE6L61ZHJWKI0zTvt20l4l0g
+eAOmF787HGCz7HqLT+C1dE4wQKabRPS2PT59nqKC3uW55x8RYOsPYrvoI+Cv+00AEk0x0FhmcTU
GJTIjePKHplGnrJ11Xy4SMDhFf1JM/oZw3ZGtQPVGrcqs3Bbaka0VJJ1fempXZTngVLrEL0tkdV9
Ffco519b5POzsJ80qI/TJSjMqG2WRGnVamBx6w2CC9IOTcBDHbJETgUSUWLUsdzlOxYHIHtpmF5r
7e3D0p/aaBA5H0G2QTA6hvVVaSXwDRoalJOuFZWmQNIMUO1BsJZqRM/Ui6H2I55tRwM1gBeoGck1
2q6Dfu26hoVJ4nU2xkfnUcr3zh7lR5Y1pzBMw6d8pgdiBpPGJvKjVTEeak8h3Z5q1bgGCn50R5KI
0sWVym7Uv29lTaSBu5dBulD9utHiR9YrU0xLgOWfCH6vUgLoAmji15xeSSN1GGjlOnZsdBOwZ38D
GVy28UuGL+ce0IevIevs4eVAq2KrQqC1AidtgbRNuWWHm6vYDh6nr6X6louyrz0si1uOkTtnpNo4
gbYl+FXpfYDIH0Xaljibl1F9Ar0SVo3NdZ9AQCME6Dux0fjqqhhhPD4y/D8zTMkBfbHz6vE9CNQp
9r8LL6wMKuDD7CK6iLT723sPmOzYopOCZvQG2uVpYLOeL+4ISfmdafC3RJCuGJ6OJjkvPt3QviZM
t5JlDNTSZ5CEGMYBy+XmlKxNqdMnbG/i3aY+Xmq67MoBjJP2skpbd3EsUrqBWx0g6ldz/Xv7Va/i
AbZOoOx8qYOjuSOGECkGf1vMWdd+fz87+QSe4bGpPR8EGsdLp+xD4qhlgYgbWa6/UdrvnXjKYWRP
NWSRj2rCsSytCfnL6oB98MrRoWpIcJo8IRMiytzZi67LoggMfGY/xEiq7xSeoM/3jCiUgBBZYgWN
e4nW5ayIFcyykTZvrDl4TKQto0Ud2MFeofVqeS4k0b4ErP37xnB32P1M/HULanV72R9JWPGn0D3w
6xd2BvSOqDt8r24VBL8n6nqB1Ta00XjZQJL9oK0ah+qgYBFHrn1hPl4gquQINpVIEOR7MJQ7OJdN
NawMy6kLwQBRu/MwKRt052UbMESSokCmnj2XYG1aEbi4PLers+2f6C0qkkuJ7+GSeRnR2o7nzH4B
kAZ6xQpZPb2Tqg2DL7YZgYBW2KGwdri4gECC9sCVRcFlx9djF4PxHMutFkJCPbP+6PQDKg49IdAx
wXhZxMwXxyuHl/NDeHFIZHb/Spi0PDinBeBRjW2b/bDCs3y27K+zsk/tQGzK0X/4rl7L8Kle99ls
IEKSkAJTLtnsRLysljJym5rl27pN/hJ4+C7hMgK/erlOcKTyTjUMZN638GT2m5jEsOJStv1roDap
Hhl4U0PgnwEAyQ35SsEHnuiCXnPe0MNgYVtwxBOuAGDXLw46ZJVk6AUoKV22pORiF3aOYXMi6YGZ
lAR5dO3Rc+xtj/ogyFebRgw9Y+dnWew1cmI5FsUkYXmYtRAO3KwGdp5TQJ9a4SdTD3PczzOQPN6H
7krms91xib5enURYfX54IJAOcRcLABc5Qm5M6lioJfMyL+wJd+CI6fhHKXDbGx3afN3rMEagPjPV
eakNJifuH6cHKWfSKC3dfCppCqTmKk3ReSuj1gTkAKMpm9lCfCu2i2F8/cVfX7PV8oOny830lYPo
GYlnmw+iiVea3SVmxSrA+V9eGs80Qwl8YX16m9DBUryra4Fk0eh5oFHQiWYiR5oVtx7Sxx5uip6F
wVQZIkprwL1upNoHVroH8WeYtJrUCsUYCeEjWbLYOlGAMU0IXowHR2oOPRmB0RjMnLMY/EqTQNcr
TaJHvGw6apcEXThW+iRSSb7viWadGxLDBsAMlXu7QWDvO0mvTJRe6y7IYOBaQnJeogGqSJM1HV5s
bKwXxOvmWvna5NTWKNM9fijYFxLJMC17ZG8xxQ/rZOAB39Qvwlv7B2P0Kue9nXFsB9hGitZH7OoG
huzgeL1Mfs+hb2f4bvw1ChdLOWgKMCe2e8GP5XI9wkpJyCxh6HU4lsSuX5sJCCFfKVguHnN02qZI
y3Ib5yuaoIGyPiEr0EXiOjy1PI6qSweVquYpOvFXerthqzIJ4bapg+TN94VMNVrwZczYGRH/sT27
Jozb4YcAQzj/0KHh39S3Zbdgc5ZekBej9Jye8ah3/E8/Z+5eQTI/oOsw79YWe0fHp2jvZa6DEj+b
iUF0m+G0dR/rn8mhdLobN3aWrnjVCeiZVp1Tp5pjmICs75IO7axvq1ECtSXBG/8mrpPHEJwRHVXD
VLKRvmAQlLTBh/ea2ec0A83VbF2gA9nw/IKj4gl9xHsayPDfSLpztvpISiuBsS8DssHzKYn2in3p
gleRz0AB3o0Q3HozfROrV3jysW+dnN1GjEjZQOzXk5lpCTeOSoyfffTyI992CEPibscCI9cinn8X
4otNfbgn5/oL1aYZlnCU6gUIofkbxavq/Yfna1QXnmrH4eIXUzWJ40wJHebK4X5qzl3OU5naF33u
4vrg+6vqgQh2IaWMJHNF8icxjz5LMdREtBU/WdpoBpTFYCoAisbzBQLDCQpAGpHORHOYtlpDPdQZ
piXgeDbaSw8y5IVQGPpfJQiYP3fU8oFxV5KF1ASHzCTWqgEGWLjsGQ2RUTe7qtbqwKGpLaDPZOTd
2DzY0+l4UVgdXwW4BNJsVY4I/3vzQLfNKJh9X6atujXBlWPv+Db53piARbC61WFIFvI0uqOtpmHP
yyImWkehF/OOL8mLHP/6NsFe0omMDFbKT0aiKOTMqalof+YJkwSqnxk7I/kUpE/0QmGVlXArt3vh
1e1oHblA/mx80DU3RoXUlqozQ9F9ZzQpebxTeIjPltckwZ9K2bvT3LPE02VR4tN/rDoDp8IjoA1X
RsSs+ZiVkwy2Z2bdqUQSgLBX2+Bqv6U6sHNsErEznTSEQ5ioo7eAvw4toqu+QHVXZhgiHF5EKH8O
132liBSvLqZ/sgOzcWrUCs8RbSTyIcJF+5vJ/To/1w9T3qMrYaCiyPrIH7+D4ulJ2a9bS4tFxS8B
dR7//cF14c4KJgG1s6yXW55Fi/pJrwfEmNZVtqjJEr61PWZ1XUWRnytZrG1qi2v7p25m4svwYt27
MfHshr4IkGuMUPWIPqy91iBHldCvO/0SlrqevP2yDD4o4+aXr45hzRQn+j5f+WWZdCJLXzXnRJBS
1PiZQKGS9m5m5RFr647CR7AYLFXhjk24RdZ0LfRgr9p5yRdp76foon+6qXSF+XwJsrPaI7MF6bRQ
linyaTkpgjQABp8NNT5ez3EIbaJIXLOrqzQDjF9bvPPKN9gCmiLjOVAF0mFxgd01Zv/MZcLU/7Ma
UR6owIXgQdBMcaqlHxIXlYV0vw31xxrd3K399X1IbEdhfnq6LhJKSd4pbfmWWbK9e7B8sW2Ue7KS
D02J8lHantFH9O0mSnGwyb5OCuhmYy3hg3QxH9jMNakpa3i54xuuwZDEihEbyrR1wBy5weqI5VJK
C57jxpgFX8NDPMa+K4IKIF+W3SC413Zgjn8rrRbl8MgQnWpEzJEIdYiKIPoCq9K8jtUinsl6uo+o
ERAUxYLaThliMdRtMoMooqFA0LRxfk53Ky5wXmYPuqDT8pywCDdzypmYhGdnB9CHV8w+Dnm9Xt1G
h1ytOSiHOfHeHRSuoq3GirbMGRjQffvjXIea2q00+AK8k8vHWDvCVo+jxeuMUxGNBkO7q8rKcoJr
Ro9ZIGd7om2q6PhaLF5TTqMfperSQiBcisadtrl7KphhZHR9g7OjW2YtG2HAbG1e1fzPxLfgOU49
h9CH/AyJqKb2fCHeysDu97PmDG6TaHivHvB1gwHtSLURf0anz7VBUVTcnhuGb0+Elg6wWgJLWQpj
zzxti9l7KhQUvYGGaaQIlVAaWcdPftRKfCF33tCQvru7eZlDFr9Hy1oBH2oFsQ9ldlY14jGa7gOd
0/QPfICB8U8F9jvWtVVs1uCZ9sBV3bj8ts0eVC9+g4uXUJpO47LV+fkuKDXH5XbdraUZeDIxsmcH
pnaHC41684h8zr3QkJt37dpmF06vSWZBZRPYf1dKOnqhTNVaxkU2/Dt61pAUMDwvtzqeG7gnwV6P
Y7o34xZCnE8uVOMri8PbR3TjjtnnFx40ACPJnYCGz5BJB5/jlwpkpypw0z0BD0YqQ2KfVeY8riA+
wfFyQ4qdh17VeA9UVSq5umWyLrK8QRunuO3tqpcz4EXff4ELXBbAKcepMNAtAulpHdE70CiaCuJ/
Ioiql+DXgJqHHy1UugkRnCU4yQKTUH4dQS12FvPg0GHyI2EDFPxpeO6oKFx9FvktvNj7WsI02N9D
4PcA6YnkvZzcPmq50axsgSzpn8aOAUbQdUt3fZa4YnmSXbJAbYGHoN+kWKJ6nvYlUHCy04LA/MLa
hMv13Ph5iddzHnobax44LgJiRikAMnTyksR/CSS9ZrxfVvBrPnnpWlwf3tJ5AjVGt4apxsCYMV/f
oWOATfcdEmCk4z9Tue+o5Di/zmZA8UoGDxImkeZdiGv1tAl+yOAMsPzztv3JNg4v6HIv1+B1D2SL
ernq6t4PkEYDRuj9uRkjBrd4AHCS5KMEUpq2DK8pwdi+8Wd1Z1qwmtt1UJJ0QPcogzejHTQhu+Sj
f24tXp16ux2SViTpH2f1MyoABlpjRM/f36ZTL6E3sei8yfc8Vxuc4DTYLVLibMck8csMkRw597jR
pKzJlPmRxxoANgo5mb2qEPAqU19/fnBd5cKIPIynOW+h3aqJIXo1sR3cLVM4VEHQjACVdTq0Vrg/
+nm2YnYgVWBVwB5IacE4uLIGLSNUxFfEfTKH1eK82gdL/a0pecjuK8OXGKKis1wWcdA+Tq1+lGtr
CjkeQQx48FLNsrCmn0s/gfyeF2Kj4FBCPgGVdOR0jbmErRzZp4zidSE/Z0jlrRe+THKvOo6JS7mR
raFTn1ljkL7LuKl0YPOhde2G/pQeWM8jJw5u7fcGAo4VCP8ik7jGFcFzX0oXUnvvSxH7k4r/Aaka
jMZvNk3oyPd4Uen1UEMaVkM4Us2l2kxxmjRAn+cSem1a45AiGJpNNtk+A0SMSyuVj4uCpTenGMK/
yerL1um/MTm7kBsquovDjZFUKZ8dsExNR6h7VgIJ6VkPPZUXkOdcG4TZZ8yJkCMfZccgCzmmHhNU
ff9KlI+IhtQZV2mUSowsDysqNXI1UVUV3tubL8dWg0MRYrNKp25l9US2xueqDQa2JCokKg2ClzlQ
xbRwd8zqigbFsKsV2L8xQYKtiuOWtp3/xxBTd5cgw7z+DWuKgfj4yROyFauKCBj2lPBRx2JAuuYJ
XusQ+4kl5ZU6Hy4PfV7l76WjUnDQ+SlE2T6lXqCRT1eFrLU/LmWmEm9cCdrRFjMEH3fno2Gl0qI+
w9Dr4DS9et4GfLG1KM6SDnkeLEGti7zWYL4TOAQahO5kdeVk6v5pvHKk+mWsaVh+zZXb5X9s9+PQ
jXxC0pBLMvzo/y98cZy5ChXjjBwHpEeu+ZHmJTUAqbWWL+ZQIWsUfn6DpgdrdpTm2JjegVRxMoTk
gxskNQCh26HlBV6Z+qo71AaePCQ+J2D/2eiStrX/JZoZDVVix3FeQrDg4flvbBEC3L8QTSRKxvbO
vx16tXGCChycLsFWWrrFMx46dn7ixJB3p/vGeZhtVaeqm6M7U6tYiogVf22P+8MkNLAd1RNQcX2T
wFmpW0Z+QeLY3dmsGR/DXVC0hEG5zXMESFYrEtq5FdFaQgJAQ8TGJZIaPJ1Dncapkksl3xwhq9Dz
6dFnrjN0vgILDR7i3If4I3Wy1wmzm3k+6srhAB/I6f+m1VWKTKD4LEmgTKpr46Z1km5xPX/pt3X5
IeP+E5HTYNmal2ej5tdbWVc9U42DwbXYv1uwEDzVPNQJeo6UR+UpaQWusSWKxLWymvvoEGVMTzOv
98jyr7aiSq+NsF1eKFfbhtX8cEgubcX+WLwXLHhMD/RNVf3RkFMSAIL/AcKCQKCaiF9NHsY1YI3d
CQggEi9ZbbVGMl1OWQWGXMC34AEXeOlyCj0SD9JOK5XAX6IZxO/EHhVNSwg+1pZSfxrh/c34x5Fj
u7Hv1N1/VlTPhRzwxQ+/ORF1O3Ru9jSwaOvA4CPpaKSFMBGHaEbjqUtfskMC288ygaExNYIfWUh9
i2mpwHnu/60zEqmYKdapEx4PaPSQa2YVBt9FKKqexhJtEJYTuMZyPSvchwvDTmUT/QbaYLNghzEZ
G1sFOI+C72TqoMwLyhf1hkrA6IXBNHR6uOHv8hzl2lZKpNAu1ZpNo3wrBu7lrhZUUJYxO+NPg22h
/w2s/kppKCJicyVZurTt/baxf8yGAykYkPhci3Lew4KBInIIbct1/2kdUOajy0I9i/l+UhtEq0LI
OsinKG3uN9pb0yu1FVtaaePxRM43xaQgR3LcLE+mn4MeMO/CQxgpvUrf52LJijltmSH/ioB7YewF
QeUNx+UYDKLbp+KhbfB5z/colOa9dub5BtOJsmyMn7jad4cGrOKTQPNXYtjYjlUFuZb+yFTxIoaF
/ieJuk1YeZVXPwnCHwLq4whAaAKGRLpzwS9lFaulUwbijtDY+OvMQE0E/yzpasbqx5loj0jP8syb
0RYSA5bKfy79bXh3IINVwQOzB4I53R/cqf0yyMPaw4PQbejqEHbo+yxuoiJpdWUX5aVuoTqcz8an
bwtqrRr6BqnZ9hzco9bAPbAgbiD4e1e5O0KovIl+Q2k9UEv7jzaMfKGnGv1cEQBMLl1baCksRYj8
CvSWo7Id0PkUkjq++DiJ6I9IMcQqzlTBCFmcyeJTpz56JsVH8aQcOLIIuzaM/r1i7v7w6MBIk9u0
ZTFzSX4ODbW7gR6j7kHdV/id2UUIsT9MzxS2mwEKcL7xi80SIyaO/LP8Mt0TrxJ4QlbNYSRT4LIG
S/wGbHEBHKy4M9JxFNceSNsY+eInkGqBhnqJv+7aM2SRto9as89xA+EZkhuO53iIt5D3SV/8n8gG
Mh7ZVrS6td87FK+1jj/Yhm47Dqd2TwUDS2awKsQdNM+sLPWqgN4YmqE3mxuKnVrX8OxDptr0iaxn
e1Y8/ylFZpojjjMAEE+p3yORDseIESeYuZCZ9/InGz1KQCJGBAkdQBbXub2Rg050jeMKurGgWBI2
aRb//pYy56Ko0wHGWA4ueAqQmZKwSXe0CNTfz6jfgHjL2hR9hz874sBKr5yFF7VRKGm+IFM0lVQR
/FDeA2u0BuDNpbGEPFbE88mXMj+nlOY1zD+MhNdnJqkjlZh7B3aSUpbBUi5TZywoeeGyKtlFUutV
oOC77bpYxtjj+Z97Q4vCSrMlIumOhEXJoSI4juflX0sy2ZDAuHZcCebfogyhxPxe1mcz557Yu+ed
3Bopsvu8WSy56hs8OpnYHKX98hzhwOSImyOpbsH9fdTjFrBIAbjlKvvYnR8B+Sq8Pe8v2Wwegs0K
HGs7707KmfANrNIkU47VU3TOLv4u1eS/8u/HaDi1CzurbSdlNxM3UgGMGLOEVaQuzg766rAvL1ui
nCaIwIQppKQxNJB6IpTCJo+6ctrWCdvLeDeC3D2Par/UMFSF57lDa0ZfyfSf5XXlPHDHbvjQ+Me6
CdI4WFxK7QLs5u1iRxAy9FXJg1vE7hhEwm7TRrtxPjHeQbvWfpfyOOSvGiYyEFwchfVNZYoiOIs2
BV1IRB1dtdKZ8oN0M0Jz2HSJkTkNy37V/Bk0r/pPsbWd63GXRx5tZbiSL52U3Jniv+wBRa1oCdkr
elUkf/ZPvPbudNiVnLdYs5+1Wbk8PvTzGEjiBRouTqlxXaaF4+RpO+f2CJQ8trLnSlPWSeMIFPjC
p8/u0Q49W5/0+P9SX1cjkm6pUaF0rG27U3XasEQFS/Ghz7w6m99JwfTAQuqyWtssh+/cU1GV+gfi
tm3XEcWczOUgw+Hk7JZrC6ONzMCljQJnm67y77hK3WeKAz5SxutT+qeyj0/jtjH1wVz7hFMmmBVE
hRcitMndR4foYdq+uvIGe698z+cT5K9Zq1lWZAOxsIRMonGza/9W8dQQeJTo+KkVv0f4X2tKb2wI
eRtBULZJq+uFWYV4yJUe+azuw1P6Yo6iVevr97O4prqahtTYFgrGYNX39QugbumUI5MqLBK2gQCu
3UgwjC8KDclHW8qtShkEoK7MgypwYcvgGBpp2Jrf3sqc8cFIx40B5ByeixHZRfQ+cK6a6+P10wq0
S0TXqzoSDDnsdueeh/S4IijzYKfXSD1FP8751WOHLgSAZSx1giJaYGNfHRER71/DiuXHqHAHhahj
l1go1yAZGdsNuSrlFzyh+cjMfTIFVZHEf/n2MzXwxP5MYSmdeNVYGxYQNHfMmij2k6zPdC7Fdg0a
L+Mj9REwoDWklhU3kcGIj1dHEpVLhdDbK9htXoOGdpcavkmOFILWk3c0Ts3rNpEIaZsP0uQM6t2R
rvsXT+hLgWV6gDxxrqVZXYNbVqUXrXLws9ZZ756Up7iRoCgz6HvFH4uhS4QR3R1wSyJdvCaeZAx5
tuGwXaMrd9SoXvAP0/yqZJbDPf1548+B8OF2C1twOO5yp96K8UyiDkkjqe/VkRTDF1JWIXLmNjIe
G2TVXd0jyMMdDIxFlbAaPM9iena6WKDMElFkBMYPaw/HqkN9/1TDM164ih2Zkw+eL/WcLq1NW1Gy
mDOeEIe+Za1ADdP+8y9UdLuqOxcP0UKgoDtvZDWLssjkcYNkLMuMP5PowJMLgPt0X3HM+fWXD5Ks
dvfpXdtvt39OJmhodqy7xt3M6zsrueijyz3U1XkPgXnp7oYkRkCwLrSv9witsW4C4XYHw+Z7iV5E
DJ67Lg/MjnyQVYVQ2Lmq0P/5WUzxhWRllYwpooUPJen6rDfx8HvKRtQ4dcVdsMbrSWlJQWhdL+c1
cb348cT/rSy9Jw7qImCLuMMCiRrnSJMekdPOxytZ3rEtmndtKCx1GkXbsYeMwX0MH8qzTWhQFYmR
kz9+guFnHm7dk2Nao5kr+G37rPOOwmoQNAqp5AIoh4ZH3Ryo8A1m/YSTJ8RPxeqUom58lMkX0UDQ
ODAqq5qv5Zo1Gulg9RgV1ByEXGxr+f5OBMAwx5Ws8ZKuUt/VsA1xpjSXNQRzmGBM7PByEDNEZeQ2
JqoCRxqmk0gJwDCVxQwyT0tkfGEzw2btJKKOviV2mZutYlVs3/hnqeMRCkstgR1wtHWT4c/9sDjj
hiHfkZFAvw6c/eH+paIe/gzlpwD6PYva1aBoJ6/eXFUD67vSWkAnrusOJcArHEb6HNvajyujm84s
UXRqnJubkZlGB6o1f5TJBtyLp7n+YhdvQdbKCbP8zvJSebi+K0HScoQYMEuHWDf5udo+PIZmVeHJ
igN+b1hcLA9Lmgph0648hh/vBCeoPxTo9VD/1xMPbRu/FXFlfmWOi31gkIj96GMqp02mAAY4RtJz
iP095Wb1FMBY/isM7XYL++p40udePgqUd9dFvrpyKiFSLv7pTROna5Q5PMQu4hmagHHNm+lnnUpO
gKlWnQgX3XxDd4Yzpk8lrb0S+KK7zNeVm/XeyRcZtUJ38KlycG0qc9EA7Igh3cax+LV0R2iUBApo
5wyvny3E6+aLqI42qX7qAziMINnSYLr1GpSWxLAvAImS0FwYg76CdmrOna7pqC41Vgo/8QIyXIkB
bBzR1j+pGzNlkeoJSe+1Kq7NdPp0iWNA4fSTHJO2KbRoES8IUSDfLTXgriHHtozLhw+nSU/TO/Hu
/1/T5ZHoVo5/Nx5ptupBvrx8sBP4Xf/BTvea3mHx3SN8A8vGXpuTUfsRxnIQbsL0RqeKgE1PD0MR
ejUinba0qHJswsNpyuDQEjskjK3mnGz8h38myUDh/w4a29IjNSdAiHA5FK/nIX6nfMCFSOq6xgbV
fC1VQjZ4uZEA21+E6TvFB3TB04etV5XMCde5UPudAT8CPg0nExFM0ceSRAt7HGGQ3wI0JuIP5ZTJ
6QLEZafpLHq/bps57mhbG8vkO4U2seHRQeB0lXY4/oE/sLwavLf3ulS+6PkvnpHyTypTkqKB/mTY
HwNbK42IjLsFantypaJTKLW45u1jx9O0oUmSNp/o+xF408zlBtnDYpQ6bEpZpaOUugakSvIutjQQ
Vu0EjX7JDbddEh7C6p4avc1j2wWREYjQTAYFzuoby/uEr7nOXsYXNuDH48RbLhPwEuhXWZKoSSBh
bnf1F6f0tuHzNkedqgxxvs4Hlh69Kx59zaooSybHXiPJZMERHvzzUFnM9fbBRPkss4YzQIC/SPBa
A6hkQn2SlIF6rzFPxZAprGb4JKORUkVnXsItinX31oqwnzk7+TqjIHGWprjVNLQts6pZOHDzmlQS
muDq+GguGLpQQCsvILCrgAnqy76voTzqLY3uXWE0RbLoOvocEqWenUYs5ByhzjNCtAJnVAN8cXBl
Lbikzt3Hagn3SU3XlhBJMMJFgPEOVuKdBcaruWdgZM1IESHwmmrq7X2FyXNdcUQ5iNKuN1n4PPa3
pwR4QwjkhUk2pHm9Sf3DHR0pzqKp3GK1SsfJ/gOtEKrwicbwKBJYYqGU0a9oob183yOBb8gpFQkN
dLUeVGNTCmEggYvspjMG3EU2HKjBqFI2ESM/KhotES2TMK/yhkn9WWzInioM45CAORQEOuBcvrjc
edACFWgjRoKPKC6ZwrZAnepb3qTRtXkb+yeOL+X/oiwxgDmCnp4JYl/86H5tHshhx0fqsSWI6FXr
NVLabfhR7Gm3UbKdglqQZHhusn1akM6DiHRKI6hZmE5BVNrF4yRc+ZmfF1fgAlKzlHreVu7KjF4O
agELvepNl/xQC93gqSG8WSIwHHZQG+cKpMqlOSzsdFjU/5q2YONmsiVKlxcnP+4KuAyoHlzOvYDS
zys4d0aVBRRSLt2iDAszBEh1OGsg8bFzay5+tbBaUj4YiVW89mXWd1cd5aTZgSjUMFZ8z327PdEt
aouJJL99Z3JzCMLhK85Bb04lhYMe5mRduWxjBgQ7IYDYqZti5ptLZCTMTE5cZBv6LoBNlyaqjaiD
+P4U5akefh/7OLv98rva2dCmGxdzM3sD9rBfDb6HKwhirkppP0rdEv5H0A2frfbw6z9ArM8YrHVD
MG1tkzzMI1MHidQV2E/llFGLdQQaDiIJEnF3N7nMxZoY719cRKK5SfeGOE1IU7Lo7Xs87tX6iVUB
q0zW0ArFY5KR2fq3qwuwbE+1x5LzAudguLUUkCQ3HKoJ/XcAa0gvDohgQZ0iIHkucafKGtmdtIto
RYDgrfbG3HE8BfvN2iQBRjEWhe3Yy+DbMPqLg8A/JDmz8/H/OGE8UuWqLDBjmqIYCCLg7h1eYv0I
OpCza0Wkncqhxlq9fYwWGZdyPSVdFuUpEpxY4Gf45UELYZOsQB1jsJ/CIpaMH2XJcYe2/3l4Sxob
CeP4k1AS79HkGDdTRSg55QWNI8PwgEmZcL1oWzpxFoiy7OLjr8a/cfBdGEYKlXgNeHBUQMAkVjmE
PmIr5RnE104dtJ0kQJVvrojHhXAiIM8Lm8ozjHZOEHyCRERvbo56nLhUP0Vi3LIZwQUzmbE8kLWU
DTYF4FW7r7qLyMo9XQ7NAY705SP4DCx/LehoI6/RPTOtCgBSczlp8GQA00h+zP6f5Vap4CmEbbFw
i2y1HJiugvMYpYcK6/qFoW+w1FHowjPJY7A0tTrhbKORBpGIxrPpD+kKHMYDBlLJS9/lMq86alkK
b2Ieu4Hr9qeJ690ms1t5Nr4SZJk3qrxCe2sYhJ5ahRt/ZpoHq2ZGTl2mtiwEQwnLPrIv24dw53Gx
1DV+eJV05zOC92Oy85nt2tFyCFoi2ALg5oXslfOya2QMOjkQBd3IdVMrsPstuK73nzNXSNcsMEBR
e6Kg4gxQ9RedC9+tMCpWMyiIP4S7yiOdZB/jR5ATqDS3OH45t4nBqz5ro/t+5ayIpTQx2EowRGJA
r6SnyBEN4HQMJxCngszWuJNdz69Xw7DTKGVOWdzzcvj9BsmSzTCBLPYSENHSTDA+Pfvaa9Ma2D9a
ddbGdbLIG+RoSThZLuYe5OFEePWz7/MHoErxiFlLGMyCnvE8IGTO9M/Ux9aJQkQERtFI5wbG7yUZ
gKWgpF2M+xTrGQXV8lCSktaI/5ylxcZHfhIatDUc5j718HJlezlpfJMYUNfojJdZ1jqUOiZvWqbm
r2O/O5ViADJJ3eH2ew4YYNwJluS2fZcn0pXZCGEaTfSvwUqMrF7+9akR9Td921jjRO6q03uGRJAo
VPo85PAkF9RrUeUKvcJKuewwIKCaLT2CNVYgYiMdJ1aMjcFSKK1ouwdzEhnYAGXQPA6dgpiPXvox
L/jCUK6S+BGQ70s9NS/bMgBY5neL9pP1PcdyvrTWDcV2erGYZDR96DmMx936WxdPMcGoXCOhfv7Q
KycBHHabmi4fiV8DW4oNC19LmmHdmvj4TVmS7R2PamcwgPlY3UeNiup+XFPwlr+caQ6tVcYpe6YA
Z+Gz/vU+g4paI4DQb79zH54IOjfT0OCfu0K6WQq747IstMDfjKtFjGnHSjYuq2W/4d8+jd65xn2k
TbFNudHPk4b/CAmk3aGB6FdgGN52b0GW6A9kH8hWuEYpU7wuNNjIkG8X3ftAGinLpERbCrsHVDAJ
ly3i5/fd3htIzTTGt707iPHb0H85XLB6ZYoapQ4Fy7djvZL+gZcpvwahh4XmNGYQ76i/hODHKPr2
+/Hz3myDFe5zG+kvve+sa3JOQZlE47+YedCF/G0Tqi1pWmp7ewYHmydmbImzanBBs0IVaTghZM0E
/vRzz1pE7ZaTXZMG1TuVbp02smDuWlhrZMHqQXu8b0jjTFqCXHHHmPhiFGcUfB90RerYjl7T3MLK
7o4l8ppBY0dsUmJBoJN3z/EFIw6vDchoBdRZBKC1H657+cnuw3RhgtzLDjiJHlb5oSRBBBk73kgt
KkaIOXbOPqGVodng7G8fggtEJQoR4aC6NgrobBaq19jGMqJvjbgOwpEComvl+Lc4inUm0R6y8Rw1
Kipr2tlCLVtgpyz0qFQIAPcEeBHjibU6TgWA2drQPJfBkN28cDvks7n1p7d+4J7zN5xAAUDm0xa8
vk+aNaZOMNQjPs+FpjE8AJymTdzZiyOWAfqsmZ19lHteLbHy4SXuj9BUWvL3P6a8rBN96gkqS7xR
TtuQet8BQqtQE69FY2gvjWJnwv1OW0NkKTXO3nk9cLKZmwZQI10h3DYwZ7jVaC01KH5pAXpEzpUZ
pIf95tXVh6fMbMzEVMV4QkH1cdF1Jtewr5utM1khBc8ol7gz/jO/gn71q41k6ipo8B7lzHfEHj2x
S0XzcWBVFACJ3DC8MTUydYEaccImwP5KIb3agKbIpjWCrkQ5hSKciYHhACOmJ1pvXfCO5LlZGAb2
MH416lPIIDeS8Y22dlwAEI6pq8G1KnTS+UYxBfEovSUdqF0BmWmKC41++H6znVF9OXPkQqEl17OP
jSlD8a95ONSemY1lcePGuevhw+QnBPJ+ZrUfpuOkVqwXl1Ne5ZVK+LpGvOwQz+beFUUrnkJFuNiC
OsodaXnWkKH1lXlkM6fQdLXuPqjcNoqYeKsuZdXiTT+So8Fye6GOGjSyq9J7znwQt8KYTI39THJl
Xf0dypT6VpDDvXGuaXj087zn9WreUgqaeE1PS4iLxG3O80wM6lqOpV7ddrHJvz44ndARmbluxwiW
EB49kk6lmei9NZwaPbcFsS6vjeXsz+PzS1qZ59s5g6xnO+4inolQSDL+AvlCugqoUUVk0kF9MP/A
PqsQCm3nMzfNy/jqRaZFLQZwBpsKaCG5xM7V9pTYLOmYmEx8gzImtlxVxWxSj0FC1BcFvxCXvCY3
e4EPlDdnAEkcvwxKetI+Sp2dw2MxGKPyIuwr3hW2FNjUgR3Vk76qMK1c7oTSJjVFThjgrjc/n9MJ
Yol4Cz6QlP4AyQ47KL6D5pniWQN297Io/MnE9olsTEz/mVbj5eKnxazmv/bL+/Ku+PdPgk1ctz+7
VvCf5eR+dQDW+JgWejArK2FHoCn93juhZ5WCtGYax8oEJChosxVZdzmmhvQnAzDRd4dPZrlWIc6s
RzeAxuhxJ0u0j5XlFbG/yxDQgKsd/MgIT5+pLRVYB0YSq/Eat1+ssI4aUyZE30Qli155LZ9ctG/Y
0oLq9LXnRn3EcuT430LmwEVDW4K6sLFSGOzj3ifv+ktm4552tXMJEEsJ8y7a6yrJtyPsb3QPSnZW
dSTbNuwjPcBLPZdkodjjAsjlpYM8pPKd6+XtCtHLjFD0pke8VGOLeDgsrtkNIrcDmBUKBJHViVXR
8KaxIgCpy+CuRxKfEeX4DrLklDx6SRO9def8c8LQPgDck93lt6qdzGI5HTcv0k9Ql0jX4KvxXHr8
tD2SM274PAP4IhHND65jP3mubhIbDBSY0A72lZhA8H4/4L6XH2ROlrIpMxfxfG5dgsO/q0C2esTU
VeTKGn6TaZqnzROPNuDHgxrq+Wm3NBSju+glZ4VAE2Jo3gaqzWUvzGUca9/u7vuLid/BuNG7+P+I
fUBOuSS05d+xevJNE+VzogFjharV2WWl09Dif9iNfidbGYEiMOaPwDraIDStf5crZTcUgvgvH7zo
iiwX3nvPSz7e+ny7Ua8pvxQ0dxMaqYDULyJ7trH7aYpUEi9d5IFUDKNoQEzPI2McL0TgEU6dgTEY
eeNBddeO22ejlvjg8ZkBQxs64JvwtgvptXMAf/kEK+HWtsZvHbwU26bpH1w+nIZwcqODZYek5Ob7
XNGg3PIPumOIjtAB+XsvWM1qkHM6H9mfWQUb5rSKFZt4hnzHn+NziZplAqtD7LhDWTX7YlZqjwnS
DqsnsXrlSB84UWmMDFL6IBeOygGUFvLaKO2gXcL6DECw04H0cuYUdZ5MYsdXmJPxOR0xgG2paktM
IIJ30vyN9fmx7r9GKfXU1MNtE+/jw6ITl1zXt+PIifm2VIIAxOnfLaiqLd6EcDu4/P/BGuDN0ge+
HborixeEvPdv42rQrvvn9YCH9/KTVjKpSXBsi1fZXzEHNWy0IzR8fsdutxz7IRQ8qVn+kzOrOJ+2
Tl7KwW/7zT2dsl+bN8HATyA/Kowk/FffujEjW8fcdO5pNFRE4pZ3aIv4fo2fhBgMv6NktdL/9ewY
vp3YJOq2xs3CQkqDmyaWCw4onDITSrGI11zkU50qXruHftTX7O+2RGp1h4jYQDrv1aSCUjJ8mhmq
+XZldF8qZZ6NyHSv2AgvGexOsn/ATL1lQ9GM21yqH/2i+mjRgjHUGLcfwxCqPiYG921bt6LWnj1m
cTVpvTUkMELA5tx8Qzh8u607LtQc/ICd/7baWUpGoLEMvVoUJc0r0Y1Cx452d7WknAT9Xl7e5HR6
fI46ehEKsIWu/Ql3I8JGvV0me2i1nbyQ86ZltnY1ASX3vs9t4L0A5kJPjTZxtGnoXPQR9i5jyKVF
71m4OBWX0tyj1IRXdJoqjhWLQLB5xofN/nUVEcj78qQnsf0/xPyQvUGG9pZZzQEdAMQyivtL9ws3
ufY2KOHavRSHl/k5r2sVEA15VxayyyLFZhdwhi5+mUrkzsfT3lbNLHK8FVmgS/JYBTAhnVU7h6Gn
LEyLUc52YOOJ4oo8OYBsFcsysmbX+grjGWL22beXPr+qRlwri2uV0Tacje+Htehub4zeafoIMbq9
OBCs3k9CLYSmieGN/R+5jUUGtVKYcEAbsbBetiOeasVi4jdmUrAZTs79HKPQ3O1hH0Rk8s8kJnuB
BwUs8IenyhftL1JBWvxvg8uGRWFMIU7iPNOr9pAqW3H9HSczFEqLZl6rR0vNPjDnfuQ6i3YSkKeP
UKUHeorLCqyDHDA/MHdo3SWn3pVLl5r2Ate5S1VvTRyYyh7Lvtu7JW0pQbC0xnTE5AVl6ZS5CVai
plJ1Kgt08k0Ne9SMVXSYu2wxcfA3twhv3VhHtFLAh+3gnnvx73BxNjri2Bz+26EH8XFu6Gj1G+Kr
V6KxW/iF1uv8WwzenF8JCVyZSRzRkEet8Ob4wpEiKG3N79kBXt5P/WJPmjXa1LXTOBVFNnsI2HTq
++ciCPbwpvSp+lUb1qGjrcfqHe5Q8kJxfVVBfNWyibMj+9mKpZOPOkoo85opyRMC5to19RZVBNCD
1dDLdLHHW+/GnedFtbFT+TsuqoxDczTAJZIb3sX7VUea/yZD7+F2amMC+cOIDD/BbIdyup3sgqqu
zLyq34apCpX5j1s2aubzLoHo1vlbkJA+4Fnkd4r+UnqGcoao/szlAWtgrZxdfXBFFQ0sySDQrvfx
k80244Rq/uwTmkE9GgIaUS8ulVI8XDrKwPBCBrZ6zCzYje47FvH0kDTNjJOK70p94gxnnD8s3I0e
rDq0XJX+wEVVIGRJ3139DSE6K4h3vPAfLs9HlmqJ6F8pLsGVbPpm8N/gRlQJN4G+AdvmYVKOySR7
0gabgEkWayHqRoidSKrReJcjvz4PQGfhVezmcn3uebNHUllH/Dnz0IF5ifLdGOr6LhZGgvnxDAhA
XwxTAmiSLe6oBJBacJND/hKSYX0zLNkDfx5aN4WXUvA9oo2RENoCbmabdoMWva9XMgQ6sc9BDDo4
ObzdBB1aece5Q1nuDTqmMAJ13qqWrOM+SWf6ehq29W2miFsLAx3zUBuGvmlFwEvf8JxEWuFZIYAG
QkZvvsez/2IR1c9VbDq03dSq/V+hcYwAJkw+KgklQaxWMC6+XopWErs6Tl3L5Q1jtvDwXrlci/gG
jzqy6MlN3fot+lHA4zdJounjPggvuhSz+vLuWbdTGkzU1zy3QVe3xgfpYVyL7TfixI5ObqEaujfh
LE2TmhDHThdh++SLiJjZ2ZXPcPyK9GXaCaqq+TKL0Pm9al9brldKQZGr+gWq4ZUcB4YFoOZVPE2s
o4YBbQsHWOLm8hHojUMywoVA9/rC1V6gszhUkGFnNaGnAVibkxxQGsv2/THUbZntAOklj+e/WiCx
yKus0vDocQfN5QBCwowL59qwaEgDQeMo0WS8Y0PReQXTctTs39e8UtntdgQXYe9CznVqEUxCD2S6
kB/aKZ6crPAeDwoMkkn4ebgi644qDwgmotsuWuDcNLlSat/gw5yWabHNMbp3NX0KgpzX94Up66qX
apzRWojQl8xhXjcFGNBp8sTp8yiiSNwHsfFIMYsTpprAhYBk106NzD4Nbt/qn8bkghxcvbYBMaH/
JmxOFHglUQCwYSBn7Aa64TlU+7EJ3V+gqbvjLCOQpN2ySrtWVGhYxCvwq+j/Khp61uzq12XN6tGD
BVIlC0uxl7BEFoooQbL7gT1+HFy8vRUiRuzKVv9XaYLfYWuzBHiWgRes1okffrTpAuh+eFxKbs2+
eyY/eXWzrFKc8Q0jWLTk8nbuBp8zNR/MlKiNTCxMYgT+tQJV1Kbe5MgaH3OeVs+/fIUTNcc+S8c6
HLKJfaNK+ES52/ieLFqdq1PD5Lr5vUfj+/mu4NnugjBmX6rgciP7/dwPNM0S9fx9Qhh6oLAHxfwi
Eu9hqDIeOV64F0TmCqAdNT30DbuTtRKF8yXMQvBGJ3V3pu8jiqfh87DLw9oxHEOlcxnc6flfzvXY
EIXSSzp5JAH7B0AB7M2ZBp9Dvd3+ydxfvfJECfDwcAHHVFvc9tIUM9UcrddeehbWbk/dR4es+o4A
mXFcvUr+WXs2P9itC33Wj6q1V1EZIY8re44SkpRlEdt1wTlqrffy6YS19cUAssBpJKKjMfTWn3+t
uXjOLpUN6GzxdmFYSkweI4coCE5E6Kz3tOOVcXuELlpda0uiAGZ3lWHgToedV7EDbhHiARXr5xry
DOsU69TFuwFbx7TK3TsB7/kgVpGo6eEEoY70KB4Ml/oL2UxoEJ7mv8vpLKH94ajc+Q6ss4x7R0Mq
n6gj4ZlsI/GcTB/pRg/haQwYmgOO0HN8ASwS8OxC3+YSg+iyfX+WqtjaOh6aT+fkNriBL5tBC7VU
VtOuh9nEd6Ct/qLBEBpL2ype9GUV5YvDeE8OT2SSNH69tXKbs6FTZPKhaBMrUpshY2iQpgE7kn8f
foERtlea9oE/CF9oXDF8CZCodjsO1MdJ7D2al/jO9h7hUaG2lHPXQqeLj2KrnLVfB2KS15BUw85t
J7goQJ0YYwpmYFy+ZDYTCuGD35mVlOoBwzj+tequkDD9Syv+ZNJlIrSmRTk7jjT7uwHQ8Ke5RRJR
97dN0SYbQ1vbaj3sPpwCpeIo9qBhrOb5soZB0UOZNlt4EQz/2Eil2XyEWB3fZpomkmpM70XNdBBd
6kmnZjBNmIA61TfgoS2PfXCnqe6HzozuUeB8Gp8ZO1jFAtluAnATW92ZecEi66h8PNUujsO6Q1sH
kSV0eTdJvgkxC66d7PK5vO4tWEDwAZeSXrzeCtoIqzJ1GiwTb5B48ni3A6dt6evVVTZPovvMRoAe
HUiJF1dKApcctkNI4fbpyBCEQHSVcZdiv+/bfyQzt309H9cpiN6KKiJUPeyGzqGjJCfkvHOUZ/0f
d0rZu6xSQjqhrRVsizSM+5isAHVo96GVDpyobc/lxC7CSxyIeiSYL4ialybpaEXeGyc/wy40LD5m
4SbXLtN6J0nHM6yEMBlITvXNWXwwNu+3OXUoAil8bHA8iiISIlN6pCYuQFRlw+F8iBwFUP0McS6R
wjVfd/ntjl/6ObooDzOaO9p4GuTkNYbfY346C18efx4HEqBYO88PX97/F1oesyaQJRscsbX3cBWT
rjrT6S6wDdYvtvTLQCfrvtSXqOZjS+JGdlqlY6+ll9oue51+Wp4JbR/hSGO62xnuoSbNnbKDhTP/
U8SVsZjf1Hzi6VRPSaf5KOXstAAOmQsKd8FHGzMJ3+I3B/chaMLnSb3HAYICiLqfGgzbCYzGyyxg
Fd4SMdbdWTjgmUz5xx3kOuQovQB439oWgBLrQckJ8gKC+sHmk+Wz7F9pGPTvuGkT+nm899JYNOE8
woEyvHGZXiiVKWiIO9z1KA2YucxpLxjaUl1JDnJb/454xfKil4Ga7lNNsb9n3PQTty47+J/j/1MR
awfMLfk5L83Waqt/r05rMNMS00oi9RaPdy8WD13hREYWXGPXZPWu1G7UuJ7+JnhWc3MOAw/joFB9
QHLTugLuiSFAUPWvOFbejPn+ej2W+imCTYd2FGBo26PlsdspDcTruKffVSYaMR47jZTmvNLSw0EZ
vMHQMe7oMBh6LdsGkuAcC96jB1CLwIzPd1XJHukqkvSVG1wSzUdu07M7kqDNGFxzx1Jwlar80+v8
OW8L1k07qkqbZqqvFM44HWREu9SblRtcYfqZSGBtuNe72v7SlTeAtn3qeC2JyZxaMeO/X6vfWt6S
SkmxPAVqNCl6WR61ITF8vzJUz/A9VWdiprfIUJ03QfUM/5dcgBQfYxX+zvU91YkQFou/uhK2MlMD
S4aujD3pHU4sZcObbY5+y+Fg7UW9cmtOpDPXQjAYkgCvb7Zsrg0yqDMP+CYkxiC2JMSEH/QImvpz
mthEq/n5CfiX2qQXkr7aE+96Oy8WTmTtWiskDov0ShH/Qe91WIDOzbD/tBjGMQW4v/G2+3QfxSuG
A5/ryvKb7gnMtV+kussPLWkQcFs97hmOkSxxerB1SFvQrtQ3ELUCW12qvkzlvGAr60ncnawaZDEQ
24piL2CYoE5L6aLgKQH4Z2fh3VWFassQS0yijZE53TsR3aLe10GcBmFVLapwr9+AweJVL0QI1TQK
6RsyBizKZBghTB02ThCLbWNyeW5YEExIQQRnYalAkXArg2yPvczaMUCKzPFRrnEmx5Rjyed/3yb8
/chJi7rf0ZhoO177t2K44HGO7bx80jGmoardxnLJUyXwHdFX/gdg0Lqm0lTFD+tjTaDyG7tVAJW1
gWiyO7vhL33PZMdn9Uax50575IaVdMPt/OQ34hv+utU40HB115J8cFHSg8d9eSHxDlnw3HfKEerr
2ntlSeooEkLmOz+NCqO3VMyfEsSIr7ZhsJOQjkhXKz+bEZOzUaoE6BL6hHiEqhdkMxMr3c/wEn41
5KahzslMrYdF/UVS83rkFYM2RJJ66kcljFjWSJ9KWghXtjdbeE6hSVKrQB6/G0S06ixfxdp9TMW6
Ddb9A6dJhdEwhWDBtNU8b0pXidUzKm9us3jJWYZv/ACkL1Imlcvxa/qm18Q/5ZoRllP3Gwg/tDKZ
Kt6UORQTWE2VTuU5WzFyzPtrOJ4L4yu1JaJXKS1VW9WI9MCLCZHylwWecPIGY4n0Mo4JQ9A5pvSo
QFw3/5cC90+TugUairubtqxo7ylX9KO6Bf8AeHT+mz74yJPQLX7kgtOT1b/o4vVoMqaUlAvwZCJl
KXEvWHq5FXszEihJjSF3T2yk+DWR7gtz3Ue9iY0MN0uxm//oOKSJmTsMrW3MFyv5lS90SkcXm5jC
srzbVFQ92yJcKDC2OPeXzR77Vod2ylvh7/fdkTMJ+mEMpYXf7IzCllF/H9cY0qJecsuVmv7IoMGx
s6qkp79N1Fzz+5QP57po8K5jNLAjPoqmQi42fVqwPp3CWtC5LLiTzWlnWMsj7CIO+4/PpSy6XVyu
Se8SBf4ubPV7osIXkVH9uL5WT3yznjodZRrORz0A3bO9CKxJNsWu1c5oBIC56TLclUjayYuJZjut
yxuLhJy6uYTjxbHJ+8HJQCBEuvof2+ggMh+FCWH1xlbq9sv6gLdILkn9fWpQekP5AxDWPTkM3JYq
4BzLK9hMT4Sxo1yonQhUTz0GsROUglHeB/FwIfEWsjuW34X+JC9BAnunqemug/naC89xDH6r1xyh
NKZE5zhwwjB/JVi+M3vbUoo+gFbPZm+yY/l/Gwgz4A5JpNE37DU1FAWFdlgQvSsTXJwfKSDLt/SG
IcFTlfWJTvd6QMjnaLo2AZtqPJF2P31MtcxKnQtYEg2hYMdd4hoyKi5AsJo1cmwJSTPbU0C+a1h8
6ejL78DLuAMypww0kyYGF17BfyDH6hWKUJeJgqsp/T3PHt6FyGztbj9afHtcQzdPkex1SznGDdgg
1rri5XnIG0uxqCsrxP8mrqd4CRlBWLHsGENsO/zSxTc8TtsKYWHzrV/zYvES57hupWg6ZfaVS2UR
FRBCzO1tmKQ7m0S4xOKVuIMXyFd5GdKgZc0WP2cYXjtpz3n/2W7M+lIQ1oILlWJX27khCICmNYYo
EBV7mZiGnLu/pw0qOksalPJVv+Tz0h1NhqZMIt7xpogRQ0b1CNvtw7LRi1ot21hHi7DIsQKq5Nfe
WoflmswBztV59MfJQtlbFiWMISDYem4l3BPk0BhoJXfAgQePo2yWud93StfAF389efmJLcjVbRYB
6ysDaripLOLPxRQaIW79KZX+dJtSbhpT6yAZ3c17mEoFY8s9lniCwLixHR9vKJr0Y7FlwOukf4ew
TjGaNNEsh6fmbGTzqEnAkVusvD3BfOX7ldAO6a3yyuoVemnLQm5snbWt5l4oHyDizN06dYLaWtRU
41m143j/sxeYpRN19GNW9poH6l6UDdz5KcGoS8MMMKCzuK2ADv67b709+1KgrA+Jlho0T65WLNTX
B+xR8gKYTwPLPPB/KE0kLVI+IEu2+SXxalxt9T1gMrQ7NcpDCIkp/LP6VrRIMXLnkzGfmxZm5Vod
SWUQYKx6Fo+nOtHfMnckWh4HYUg2o8E1D8R4fQR+jITNH9UxDUlWZ9ozJw8ojBFRYO9EzixlPiwz
iScDUc7LIIZc7I+KXtCEnf05Va8wOwIpolNxFBM8E30JNOR54GZg5cVTQWouGp1xkwQa2ZJ6TdQx
X280Na7H5fmSGV4sf2+7ACLqsH9dJ+c2Pa0DcbF7cINc+xNHNtdNHtkJaFcEghpTu3DMyiTFvqf1
nOwfnd/Q3vFO19OsgxXt511RRf5lJ0DJh2NkqAwopppYKndhFVuP1BJesFrvJi9I2B4OBMUivi+X
00gZFKVMzFtJ1lVLEqWrU7uAHLVXQlbMeQtqeg5Rt9z6cKgQgur3Kd+qltECd95t8awEUikYUcZL
HkcXT/V/q/4L1YEdC4CpFIJYDnnazAsVbTbArF36lXRw+d//Bp/Au31nA9/bU1PN9uayf/lxh+jS
pULzm45MYpn+8nZqeZIgoFuQAalTpMWpsNHh/Cg6bMs6TA3E8Ni5hNUmLwiZ/WpfjhMn8uk0FIUM
KcwgSD3Zrgisq2ldGjelCnhT7kfG+7gETTOAd8jbhyRNIyu9mZYc5Cht6/vygg8IVVz6C8qaEVTX
7ywURlmU/CvZgFVdoq0bJrXIiMll07v5dGj+7ET73YOo3eZ3qLHy1WP6hwzhnw+Hh/evP4DmuoZ4
ltDWH1p8WnmbHjv7unvTJHuieZhrMBRTTXawcOB4g0/QtQ9eCRU/wejEug+Vir+8bLxwIuONCP0I
MwLWr7fPufCzu4vebAKFJqDNz8IVg34RuN+TX8pui/sN77B1cW71ZCC6ohuC95tzJYqrb9RSZk+b
5RwBnzPCKkw682k7jYRapoKZs06FXfsl2G5IfPpA6lhbgoRrj2+9s6gMdCxvyjKq1frDHfT/0oLg
ZmlK8EodPfYFnBhGKmg2QpaxJCpO/FOLEMF2dg9uAbkcuSU26GRL2Knf9vbIr+7e6hsQEy9VJN6G
BNS/tuJ1pc6/xCNAxvHiDWxbd+F9teBgEQByJfVDEzpxitAJRoLA5Cc4Oc4/iHC+A0+bn+fO3Usq
V2cihbdfjwRJi6YCrXdPzNRa3hrjLt6jNi7TCbYtq/3eurX9CDpvyDk0axPH/emqj394ON/9EVeu
/CYVnNaqoNtEiIB7PBYfMkD4zp8PZO+walkCps0FCYyesQKRo3KN0hTqXqb6aiaX/Y+UUb922VCT
6vqgmRApeJI8JL2Sfi2M3PjHh1tC9R38RWW82VG99PgUdtnvs84J/XsloBf6cF0ShiK3Ki+RDaB6
xKss6FUoNJeLUolbebQrM1TOqT7TGcLQAqyXWwoOHRhyAT+CQXPha0M9nvx/tOjWhF2THx/LFqa/
uAxMNcTzDA+Olz5E+o7LsDoQOeSrbrdihaj9GRipO/JxA7MpGGlEGI41pNlcZ5NHd7VyY3xGmeBs
uf7nCwPdXNmHnM7hVmpxnsA35e8dp7DZaSBCSwhJW6XL/mnWxFa/ArSOg93KNT+G9vQWJ0DQeLf9
eiFtIlNeEwB4HCA/nSeIN2SvL533sFixrg0+Q9E010aEL2xzJOZ90zJ0TaAiOr9aHjx2kkzSAUq8
FGEiKaxtmyk96KLsQ6yqBMpyz5S7FJKoeusqRQzCuD9CpHGmUlVbXM4SDjKPy+WON6ehENBWlWJA
VS978erAbepiGQp0n2EHsDvMm+fauLggUL111DeQs085jagn9ioxkMvqxor6Kb8NaNXPMXoOL2ND
SyB/geX0Zq7+ga39RV8Cppd4HiulrRIBdR3J27GZ5v+qQR5Vk6LwzDQfkVQ0MgCH3xT5v1V+D9aa
FUOSaICihlKgWQhuAtVghypzMt6CUNVodKH8r98gJfmLBB5whiW1qur4OWsrZw0eGmidCM9uzJI5
wSXSgPCraPrZYDdW1O+ccHCSZyZE8rnLlX8qn5BawK42C/Ls3VI/9ReSlUWDGLbS8Ia7Yk/b9677
zUZiFHSvNG6xwMiAKTatN+tFxmj7hc2jR63q7qW4DDuTiI3rSb/FUkyLTtf6EhUhqjULi2WD0f20
RUXSqtFeswHdPxMXXXJ32i0eBsnHEmkAaLOj1jLm21khLA6Nw8Qvr9gqqAbgIezL+TAbm53F061G
6l+H8QkSpDOA51j16L1LZiHMzBpzu7uyX4s/kr3L/Jd3xxLmxBKclEojmtXv4nP3shmZSl6tNt6x
qri7icPmwSs64yzKSSCNanpPbbBiZrZEbv9L/wWK82Dxk7XwYtoL42U66hNkDh1hfzv5+QLFua4V
n2WY5o3sgsoyOOLhSzxJ/SML4i8zsHYI6duh6TIqMYAqlpYb9trJNPzKAzGJ+CfZNvc6FXET19DT
r1Qa8hiAPatPE/icL4l9fHLLplDEMbpSs7N4DEIss5eEMb0ORkslzNxbJefuCefORnF9aICGWEhy
iC8IR+fs7g1gSrbPihnuoQVkHX6YgJOOErTSbDO3mORCxdwqYOQsGLsOwPLF2osxXoLd7fmnWcKz
adgbKF7QHqIiGasy+iypyw7Pb/71Ssw/DnTFNCnddsm5z1mGTlXJJRKSMk12q5FQiNSUDb+KMwO3
aVBN0qCoY2X07nrIl/h+As9y6Tb/u3FKjb+oY+A2fLhbHh/kMIyZcBv6eScJArantdkivmNJhDRV
9GNkkubXT1uAdPl7+z4OhyKJVR9VjDFwr607YjOiFEfu1BayA0H713EPyjDudst9WAw7KwMgW082
WGUIOnwvuPAIxYxxC+rwR+bIviFyK/3uo9RaAf9AWVILgIF2XXrLJ5hJMD+FW9JaRg/E3s9xGaIf
2SvzjndQbW9g+HSgaZR34lDCm/mN70uww4/0Q2bWgBBJFVfsQQ1LRbbjuPe6ci8AEvIeI23T+fZn
pDzDT5mh8KpEvnVpmv/u/qm59Od3UKsg0ffOD7/6mdPn8SuMGMk1HWApb3VkBMrLDtAyfh4rjry6
PvrztqLUHQwge3XXah02kg2VWi+f5zd34qAVtD0Rw7Im/USTwO8b5iLyGtqbZJbjFhNsRIB9tAXA
n4QjYLmZk3FUjFdaZQ4y9cvCQ68xVy/8WJB7upilvRsiKdxNfAjB56bSAzE4tBSnVreopOwcQvI2
ItRrpVX88xJL8sIjHk60vZ66SpvIfC1vLwxwrfXUeqDqJOYgqVz0ZbQlnbt5ozEzxv0mjRHGGtmC
zxCAclfYlVDKT/WnEKqh9gsjA8yzfPHrxG/IpJj0UbPDgXCqJiMu3FIdAnJPJ+DIXpcO+Z30Q1ZX
ZPe9aN71IFknOvBzERAMn10jlHTtX9Hcd3wj2e3j7j/o/R/+us2d5SXY8dru9AvXmVqMBX/ukr9v
19qvcg4mr8MZkS/IMBNvuMa11Un0fDAJLt/mlVgxWcyBslGLwe8LSDchDJ0tPly095VTLgefjrmH
Tzl04mDZlcFBDPs6MS48Olz0qNWH4vP9c3lCgYtc87hCeh2EYnx40XM++Kw8CidUP+RxO9r6wKnM
nF+uvCMfW+QFmlgHYd+nWcOrcKV1HkB0xYbbGtehzY3L5rPUP+luaucsrG7R4qB4ZlJ72UV4ezsE
HRwZvJ/JMC52Vm7Lsybjo6M1prDL46cb7UgCAIUk6z9GpUzTxa00Wypcjt2tCwzMm2G/9kn2wNAc
BvJIsR3eCyqMQs0FnsAiOFW0H7uR3zmBXUdu0pGKg1u6ebsC2bJ2ErOm6tpQSxNMiRN5iiHaYuIQ
5afSkzxfCApY14+1f3YQq1ynmQDOp+9wA4gERGftKynq6g1UIzut3UCG7TabsydVWEURxe679yBY
4ws2lI2FPeDcU3qQeavcPfixYCQzl97uA/56QNb5zAGgCgWEInS3DcDxPux+zwALYs9EC5MoRl3P
t/wqgUqW++mKA21oFNFFbWxuTVlfnlm9w2Hed7M1EoRGv4iCFQ5MWmx81Svb8c4vksCULpSwT0ok
Sp/Vi+gGl25Aui1PX2hxW72ZBd3EAivJH9RnUVM3vEQHFUh4ycwXr9hYP1Djj8Q7iVN0KcGqMTg6
ZtKfSevPm9TdtjIAdORhWtL28ClwQlCZefRuwRm9KxZDQl1qs9hDQx4nC4vZ2ACnVb2VD2mvxUWi
+t3CY1/qusarafLeGpqOgvOyEKl88CorBoArKE6zVuC2SqzxvCZI9NVxdqw/2P1J5pZmXCEqy85W
b/njW1aq7pmRy895A4XPQG2aH7cenbrkOWVviLivkGZQcrH02zAF1DE7gzi9egIfAZ8UyDgUuxbL
dwKHpjMrT9k2KfZGtCGGbcIIjsrpmmx/bU1P7pPb63pKOIjeEhON0L92F5r0YsG/rQJDxLt63NKk
4JkYqw5KKZ6+OaU9K41j2MEkrJG+rbBnusN4xxy6d5PK3hoE6i4eu9DtBVND1yFXvTSCLeZvM9MG
1+N65lVb4/P7H5q0VkC6ImKgiA3bnjyaP3+KJ1B8tnFdFnxWWZaFU2GEtSbBWm4SjiYbOBKAxKwP
jXsjDof1uUsu9EvK5n5msE5j0ez7hIoVcjB49QBJ/z0ym2OTPyVTtCY0dXdXYISryYGB4TgO5nXW
AIJsMlbbW+Gtf+zVQ9FUlsj7wnEqzEx90p11joJyUfUGGtsENrqBa7t3y0o2bRIfUF23efC1iEC9
KzjB/kmv+5JIbCHXzohT9nSHAOSTwseZ1z9nWrwF9JoPn2Ot4Qvb4XfIrVGUHH7J412+aezXpY2t
CGQ2HmV9QBMubml/jkVOJ7beFgs8auB+6H/c48duEZnIHuHZGNsLrJITae923LXOjRMo4JNxqGfc
1ZM+DuG8zuei1hTdOEs/71Y9d0mowz4ixyS98C9K/zKOiCqF2r4HjiNY0pKSrKw0tAr00BQQY+ES
jm/TUlVQ6/Sw1GgvIX0K7OYb35Ozj08nIu3fo2R8csfczUg66fPIfZRJM6gjCc4wERlqfsJjxT3S
fqT6r4RI/BERAwaB8tt13+ibTpOCzOk5UawAP66xIhp77j0+rMzFNoCiCPOJlPJzki1ahZSKjB/e
uOwISD7zQZ4wXQL4kJF0dj+O3Mu9+1ExDaRAj3LcYm4M7oegKS16EJ7pP04ZQxr8VmOYvhn8PnIZ
JGTaUGrf9Ngkp5EI3qawEQMmpn0EdEH1SQxh1y2s2ERNOoSWVlE4ObJr0Ssmg85ZOUyAERvRZIrs
UnKil5yYXgsB1Cv54GFYItmkWs6SPx3J7L2pNN584a67WPNuoinP0jzmdSWkFii4gl3BtqD20B6i
JcWEjIzyYjBi9Mh/YbXKsqPPcV4lrvFpOhtasz+J1513CUxdN6il4aeSV/bTTGdlmDcMsu7ZvkGs
TEFd9i4Xmfc14muqSb05TMvJG8EBFMkqS3z0VGnY4XLaPLW1LA4HLyalHzV3TrxvNljF+bqrRdNq
F17HutWt2jrIN4MvU87J47gi9ALJZRPrk0yJ1JNe0frYJNnApkh1shPyOKNqzg91GLgC4/rR0wdi
5+Sx/liPumLfw0xHr8z7WQfcFVVNkLQT3VArGsTqKlYqxowVZNo8yJJEyafiFfan9M9ozL2jQrFg
Ez5jmPm78u/2YcX/wNTbRqlBAQxg5+VSPCTYsexu/geyzSFjohM+Z9jJEO+aKAsqJnfQXvXLXR8s
7fjpfBH0HrpDJowWDgprWaurootSI1rfzldJ7z1/nfe2NiGzXty1rj6Z6404SqqW7gwantaNnL08
3jVw8Opb1o44NE/JXV6pjB3CWn+2s10w5PT3MLHoDUflvfVY1nRAM8+XtDUjrUIc45B44M5nLH3g
EEJP6lZO9LCN4ETchMC8nCG1PbY0w0wXBnTlJONp0C2y/q0nF+ZlAYH+W8/BvHB7LefxYPalM50k
F+V55eUPECWJgz8q42fZwb/4wrpq52kkvaDylnIWS9PbmMNWy2nwF4f7bcWkVp3/W1nnN6rcjGND
uzCt+06U99tu07MAe71KulOg7J7F7SXSH3GjdEBMok0IzifbWbkulKkXaJYAH7Ds4CQTZ9QyBlEP
c6OOB6lEWxpy24nzAz+VJM5eK968s0aTLxWxiuTDN/r6gNX0k2PXxvnyNpYwI4VLwFLQJMoXZu5a
bDZesofzW0Lf4yY2O8+K04SZ6D6y5tYB0D7JvsreaL22fiSn1X+tL8AwSiMnSl5ryVwdtF6cD0kY
6vURewuOZEyxnd5K9AkxCBjAqa12PR0fsBope2D6xq/4oWD0p7+bxnKTHvmx4ERR9VrbLcVolPFv
KrTufBdmlLccHtQFypD4kyEJwAW6t/qAdi+whyjf8XWkgwDD7veEVMIKDPBRrcSQoJoV5Hi+PQF3
zoV4Bbu7ymnvhot6Oub3RNNq+i9/FsL+x7ccAvd+H16kvQzsMYtbW0wIhZeO5ixxE21DDv3B6jZv
yvUzvcCGMH9p9pH7EfUbf23YI4kRGlYrnFFqXYBhy/rJKya4G56zUrIei/rhqJFycd0Z6BfK2B7F
LVfm6QuLhsTZBFlmkjIxp9tf2VN7/PYcnGN6j6zBF/UGG56YQGabkAwUOJEhYWPe/293tUCEOX5n
re7v/AorP8+YXVnS1g1T9SF1ySAYMmymkfi6XZQ3OrxFBICYmJJKlzogGnwdXn7wJJahlo1yX036
P1JdQb/q6NWXjdZwZ2hHA11zIidIe7mMOSw33ZSujoIQt8rBy9CpIDTGa4Cn1d8/nj/7VZFtOvqQ
05OeN80mSmH3B61zhtlIp26lT+VCDxMAmdKbkfnUHZ5EJUOuQQGOoei64ECQgRmu97aor7A7icL5
RfvuheJd5xnOclALyqbth9pMPzA2kU3hwu+dsJCDvxsx/WVMS7UpFv4cPtcJpGYi1l9Y/djuzHVl
U0teymp9gkZua8p5DMYemfSYA8XFUmLCtu6HjLenZmqRpB+Q4JJkLlToay+Bra5zNkDhMLwsk4FT
vQ17iHeO2hXl4cnY/f3dUY5VDMC6IZ4fyZJCwzLedwb2VzFDygguZyHv3WZMDU0FSuz1zinZqyKG
0EStbYviB/Y2R10R4AHSQBtablnlGqXwXlPy2ZjsJrL3ClbXrowKp9WlziZi5Hh5yt4Mb0aWL7F9
Sw/l2688Gc4NzhUfBhkuneTjF7sOIEmypWI+AwapJhQtde+gZ1jr91/wsFWw0H4j0d35RgVeEoCx
whPkydviqB7r2f8IvhBcR678PiETPqCfV2pQpvx9mGSmhzYWkLth+JKVdbMMDb5cc69Hfep0MM1Z
LKeFxYUJQY0TMMvUn7jp2dqlYbe3rJbbfQ00UJ/S0q1kq1fCcXGn9hDG0IAhtwUhxNr72SbdsNJ7
6HYSGZ0vfDp8SDoPMtbnecT0rWWxMa3BMUJfy2j2wa84O61TBdHHkSRSLYlLis3lzA8C6ujBJRSH
ITK7wErMLx45URl/mQl8lTPIguXZKLfpwcrqLeiHJGIv5JlL2e1xRb3OQ0Jl0GROdagtFcU9BrkG
nXTvS0HiHst5MxXCp8+oV4CTTIDfjLLDbOd3vKMMiui1Ndl+YQPLKkQdFMTbuug21O1GQC2c1JSM
9MVzKM2ZAetcTC+gXnt5T+7ZiiCOgOmnonY+HcrDPU4deX0grEyK20ffOtNpcsHJ6cYNap16X1/R
FzWtp0FZPoyLSyeV2Fe4FwRvRt/UOXPJhTYijvo6Csp8XCYYViroW4PP7qDqJY80wnPIyDXJ+4Kr
0AWi+wtbttW4Ha5Cdp7vNbqUN46Rf/MtJRD+CccBbzA202C24VtG2DVmCv12JhmSiQhHuF0MiHxQ
8AG5iIHAprV6aGG+6vpH5ifB2vfj7EXjfbdpmNSFP0QMIrgdUS5UPKf1HZBJIMa8tbCQzWS/CJwu
dzO407qy5Zo4Iv2sxDyaN/NSpz/3+dHq6Np0WXFARSsTP+rIYivt8TXkRZVorZJTyQopo8sA7COQ
P4qWlKvmsCswyhHTXAUBLY2Hhk+DnISi5bVszXxrzyqVMpPK8Qy0D3yOwIOSV8rU40pSAHRYJ2Ub
xQTKVdIPYOMLnhLs9RqTuG7wF/Q5kczzdmUZ4urGeM0YjwWXcbtX/HGSNThcSLOwZyk8FATn6bRz
eftC26iFn8dH4LIMeKFlv3aJApaKI79/+osFFjq++XJGJvvOLZBdJPWkKm4dAj8o7aI3gbSNvwVe
Rl4ScDrRvyE5a9OCdBxB1j3kUv+8NV/pHnfK+ck49qonCdpRNtBi4Fo8LjM6Nb6e1KIo1+mjDbZe
98LnO5cF8A4qp2SMe6WQVaog8HsiyuA5phXeGQm8CPcN+hCAjSSNPsvsOTxVDstjk6nq+V+yI07q
7a67TLZ88daCajEySg0/4+addKCLMdcGLzwiHqx8LCPkfIACRF22BAn9CAZDEbVK0cnO+C257KAB
mzLPrMSiqSKG8SNbJg/2b7oA7ImDKucvLXQO1D5DRJVyVOQYE2MH80uevenAuNKoCPxC0CxFrOwi
AG3uJS0v7oo4TfPNWh/hBQ+kfVcv+Dxg2Op1Ou1rll77PtqhFW5ngDS5qhpNV3Gcsp5JcsU8E5Jk
8cxbdFkfM1ufjyHJL+4Ct8K+faI3llUF1q5oU4YAJm5r3dNxhYgJ3/GJj0jJHNCE+m0f0RzKVhvO
DMMjmCNiA5YIDMTKr/PTf3TDYnqRMQq5TSzHNXDRqNxMDor9sxhWF2c/yHkDAnyikXRogSv4UwIC
5L8gXBoyk87EdgBYDJWYMKtQDup2JMgJWw6Gnvh4t1GFFZj9rUfhHMKUYirvYGTpOWS1KUupE6jL
lPzW57umgMjSjjqI/aVB2pawkzoDhSlIWwryEejI8hVr1HldQRk31giumVZUrT1/sKtp9iv5O1Hs
9kChXsWBPD6gVQNPtzyfQOD0l9aOYNoWbLU3Yr6rDjDrFyuqay0MqnvfMQVyQeVngEfRCwdP2AcY
LF1Hx4tRZWkPCCJ0Ie0SPvbtjg/BGcd39Gk5XrXLMGn1UuPGpt/pPjdd/jPcBpnRY6fvIXx6xhDJ
bjRKf1qxZOQrTtokiBRx1g70FXIVi5VN3dSsFpWVuNYoUXj49RVIAIBXqaDN1vWv/k/hoOgYc17J
E2p5vhg5bJQ9n9i8AC2seOFYPZZAlF72FSW6Lto61r2HkNHGS1oCkbssuBCP0pNtNA81hcrdc0cg
miWIQg7B/keOpUI75ydA8uPApPbtj26HfEAzPwChE/plBObdFzDFxr2oltK6jLR4+1QNvEAKoJPm
Pe+RzcotYNCCBJJrAfGe+fFuc5CpeIYWsQF2G27GmIwjAsm9PAyQ1xjDXOOHeNMu6ZmqBzUnfv+Z
VUcA35x8e1JJQX8MYoWcZOhf0rtVN0MRyK+dSi3fD2ch3Q2EVTtL0CETorYM8Bma0vF4SKhUz83H
ZXSh/6WfL1P4+eQTkTcWIbf4Bhv+/WHgddo52k2ErjDlWYDswKz+8i2T1LQ8UUdFfJ+/eqfkpAgJ
34q8sOu6zJwRVlXCSU5H0WoXcYypwyQAtw4zL1hefixT+a/0Y/LE1VqnUMMulxXpkS4KCGCR2Mte
e6fx9JbBIXErRQ6YxlnjvSsWxM2prONSO3w9B6ZFcWnllyCNpQdt4z1zbsmhZzSzL19nIaLHxu3w
AkMp6BZt/pcqjHc3ezOu1HMWvyKAbOt1JiyrXpfn9Y/YyfVb6rwrcmztCtAHL5P83yv92h0t/lYL
E73qqH9/XjGG/RSpuLx+SxkCR1DrdAEb1z7xuVYiSuPMb60zzK7vwbE7YL85/j8pk4AL6UaO7Pch
TKMDNN4wVfq+4uksWBrie6s4TLitp5FM7lNAZey69iW5JyaXjhHj/NT81siCn00+GRJupDvfULDE
I5GDskl15NOWDNwiOsV6uFc7MiSEFOYihq2Y814kww0GyqqesTVlJBsp0Ga0xXzDVbMobIjnFuoN
xRmk2AOq5qKo1L82g+n3zSBfEK6m6Iw9f8xeJgWHXfIsNuTVt6D3JDQYafyM+yZXZaw/GZNv7AUr
XzCJuUEY4QY4DJIHYNZoM5kpqF8j+cUuMfQ43qUwluHnpy4ItjbBCpRPwGxkrrI8mBBcXsgWSIsi
C3gR7hokmFpX3qgoEhs6zTUJGHVE7Kb3UKV0SW7eD8KTPsDdTVTr6AMmvey2zShCPeNs5v1xXmDK
QfDkc1ukZvemZibdVZIT23YhTBbT8GmIXG7vUXMJzmGe4vaO950q0ifmZaqdsenLXmG2z7TCdtxC
K/Y8T/wQz5TFV7WcUW8fZQwfNYgB5EX4xOQAW/smSNy8TBl75FUYq8XNf7JOkjsumkBhUd1wj4p4
6hWNHVGwkIeBmzkMgxaZwdmGIYN/qTnlnyvR6A0OnPE3N8Mng3uiZHxEeSAYENe2ayrsEfC3LHok
quiVIXxoqEGQTDz81xbaIW/0qg5cOMvOB7ZaA5gI8L6yr+oWbH7WxMruwZTaxY1UP9l7ZUgMzzeW
CBlNxXZpyMT0drxsqO2w21MSEPVcCnJFMvdcAlGtvyfydEuzNmGf2yn9KeOj55Wj77KFNvpWpN5V
hPl9NzTTv2mMI6QkXW+5noJ6W8LwjL2LZuBRSi6zqMsQAuT9U0/Tqra4gPQh6qZXoqlYrH4HX4Rz
Tb5joruRe/qH1n3a3+VVMxw1HSvE9s0HuzX/71aX92QeF/yjQYbzL6XeIcen6FFqfgpu+jQiccAa
5dC3Sj9NMofJJhilk05qJzqnr1733svN40A4RDactRMFNeWWOhYokX8AByBHVNErr8G6afn8FKRx
Qc2CFpw0Ojj7UQFF3zIjyNP+RvhF693O8ojdiv9/9GQ9Mww6bmYlUSZoXs6Nt8vijwHVof8FeyTF
c4AcnPOOW0yafoqaD8wb8Pln5tfDYtLyXWqn+I1IGU3k8OweZxh1yBejsm9k+PI28T6FfYtu3UDQ
dxcevCnFNCo9qU0IRl30TnSpPRxLyifRxQXeM8agFLP/2SqKf6OC6WLyodLEAp0kb40+JMZlSdRx
ZIrpr1HZKLDHW1Z8Ny2cQ163trN8spqqSSwHheLVvVXsiU16GQOLc1SGw8CVtKzjdbbv1nHEVDne
YvXIDtC1NuW2R2PbvcUWTAcxsT0cTAtQWSoWYLwgltcV+pvJHNrqi+CkKcVx1eXiZqhu7GG04RQF
oEDVudYLaQGewsqz6YUFRwe0G2tjDgPELdIr1KftlZAEjFqose+UKp9BMN+hZeh4JEwd8z5zP61O
OeITdHJyK9Rio3OnitBnPUikxC6d9hcxt3VSVdmTjj6o8mtLEfi6Z84Gajv1AxG8y2DtJ13oqYYa
qiSTcgO+/afBIKxW9eixfLsPyQlOGepuu35rBDm4tx7LOqTuhm3CG2k+QU6xxLTeJO84dfx0ZA6Q
E1Ew2SR5ud+x4vaoM2N8NRNjk3rTmAAG36+hSpO1vz0txnmp4MfBNmIezSjLLGJJQfJKS2SBCENC
arp+HfWuDw9oOObGonHmK3iViUZ5aoJDnnPlthHR1oOMSfryspV+xfXdJ3Srwp21pbf8ZZy43Af+
Fb2YsBtoIMKO5I4UK6ufdeGCkcnwDU1M1iR4KtflbgVKepmM9mo2uQTL0nYckVT5DsCSBF3NS60q
YFG+YPmdjkDKkq7V40KJJHx2onmkzYJnw4R9DaWjUm6LHVy6OfLFox/U/Z8MiNz8AeEt+W0FX1be
OqpFPN7RLtPblpIjCIU4Rv8LJz5QNWFCt/veSMyN+6XHqP02ytCIVAZG7+7rpr63W6gifEcvcswu
Ew1tNF1RksVIMisQ4ofeJVtiav5zvRr3EKagLnDGSVrI1NNeN7Qh60py6Y72Q5qD1GFDSHy3tn1Y
TyjvrWd8FgYD1hTgjnoMVV2Gpm4JceQc5SNx7y4K42sDNJaA76SHj6RUJ2geG93vg2Jli9iEYR6A
bQO02AaIdJsEClt/cm5qZAdgCLxmwycmcGDWkD6c3x1Mpcgo9oyaFkc/PzXOcmYylGeJXbu42+wf
tpyc5Zs09Vk6lYbPS9LjcV7G+jfhA+BercS3gnSEemzNNJ+yIqbRhTTw0igbYviEtEgUTNQxo81i
O+T7Cchg5UECCBuNUGyPfj9G5yTL0T4BeR2e/68VV6XkAM+MYLvBR/rBRDlBnleZH6hDDy0WgXnD
Lpm7PJuS0AnnO3OYMOZoZsmkCGWnmd/GI1IRk9Z3KhWTlodT4XYE0W6WeeVN7r0jhatrrOV1zV9U
1XYq5Ij7dBbJvhQ13JDtRdQ/QtziPm8Ilt0Hc2TTT5sck7EFppR0sgeWb9ZGVsgN9xwefgnH0eEA
RWNBAMEigtwfBTykNhSp71pWHpqEi1ec8ylPt6TU52+aICX5wGzxmEY+eUv65TnczLGpqOffs0C2
amHBPVWBDlvmlwQY92JT1K7++FqZkSIraPE8CaHB3ovneQGySOPUXupVxCipOMkKi8PFuXLVZGtW
D+r8IIjidP1bBbNTdaY91ylQX9iywqT8iTMRyqB6Z3GGZD7A9RYgL15q1HcWzd86bxJOSuqt+zCA
vZo8xu/sRi2mbkGmd2v8JCJJ9UxCUGE7dJVN7v8KqJ9VEkBy+YMfj5FZtrJST/vxfl9y7ljwjqB7
PZbPMXJi5D7kjuixYEotu4tCqZhQfpnvf1n5i9iCLLbMsO+80MBwhsu+Cqcxv/vYfZa4J5NFll09
Ti3VDSyv27CuCuJrkB5LJk2l5RcrX1gg80W/HVUCHDDJC287k7435hnXDpmixFKCjQhArRejwHlw
MdkWHuxPyfb9wJcCckdCNCMqapQ2U1RosAcGCx7/J3BmEntttECJg+ChljuNpM5q9k//9YrFxD77
2fWOTZi1eAm/DlfPbyhV4/2ID65kUJAJNZkN/OOGcnE3HUpWPrWEpKRH5KsQMqLw7ueiymfq23dJ
MjX1a/mpZ7C5lum8EqRF1IYZUq1icC78CivOmchSzi4La2iplN7ybEk8TY+CD23lQ5fzikYs8gWy
Yv/djrZRLDHi2XDOnPkSgTn+AuKHpWdD/tJf3qNVgkbduLlklOC1tvagr1RHOAh+jErCS06AhKjS
5w/fjbC9Ii4xg8y8zBQQ8VR1QVwrPkyPABdGSibmObyNB8QIu/0bqY1BJB2q4FX5dVAP4ELXqyZC
CXdeFoc0kq/Yv1d1XbyfsokwsNkZh3cdUyKiO+k7GCXwv2b2fgjvWMGj96qiJTKUM5/ekS8bwjCx
6TSuUn0qEBrNWv3u6iXZduTp3amnkKZ3Ry22oaMWoKva9WAy+0TRSkc2020JC+WmMfFIPI2Ayjqe
TRiijORmaYsHH8fBwGDlCVK0eChPGXPyFDL2aehLi6q2ITBzsgcmgIuTZt0NCYp5abP9nsBVBWR5
ANwqtdHEQErMM6TG/4DkTn1/YdVR7nuqG7AXS7cLZNt4OfQA/nY3Sdj8pVjPP0bgTjuNyEeMAHI0
uH7WSgJ3fkS/zqwB3x4/lR4PnTObCvl7Jdw8akelGwn7kGAlhCfAfG5QTbt2b1EGalUmlGZKClpY
EBUTFAS2GDP4xtqklpesMpQnzjqa8K6OMhkKDP0Tjf1Rmz3daGRKPGInXpfO+w3GeT50S7wyEei5
nH11/SMS7t7iB/IGQerqm+toputCCy0GfHqb+TaVv5G3gwKR9hgAP+fYHFoWvXUOWxlGVBNdGLFy
zyoGUfkmXVw5cbG1384FE6N2M7QnfVeoEGj/07hVmdLOxKzxQT23wz1WiopMlYrk4LVvl4lTkLF9
rf+rXwlaNeq4xJuKucHsolSbNIAq2eG8lCbLsoWjEzF58bUqK5PPY+mwPmdAzhrJj4GBoqh75TMj
R/OE6JLOGIsMPam6UV0L9t1XNf1fAYfkYOggvghYliEvYr+BQJFN8ZLW/lQ6Pt/kJr19UHX7Hqs/
5D7EYYv/v9ARI2FHEEvHXGtWSuw31LiHFLBz0p8o1pjOgpoUvCGC0h2OraTb92h/LiGX8cNsbTo3
2D6GGJzamlmu4gF0cDsN93BtgXmWe7S96EGv5FvLqVYkQgdaG+vVyK7E97VtVvCDF9LXQf0N1u2Z
l5cyqE5GPuZtiJ1BhPKOCNd/ipH7Pef7AbUjD0/NngHvny62E0Vv6kBnUmd52eKW2crsV2Rc+5jM
a+Www0+530k1lUX6u+o0uMQVIscLRzNbg9z9T0guIR7Ug1OZTHYb97DotjztFXMdSrOjI/Ku1gqX
H9d7nGA9TAYhhN/3CYJ0VHdHyO+x7Re0mMpv9bTRfOFw4EO/oDUfc4Wo+Z/U3AiN1wZzyoh9tNKj
n0ra53R7X9hoDbnr4UvbodIClcqblcpTXdhCsxTgcIv4PfS3N1zc9lb+ufsj27XDUOxsKZaNhDr5
JEBqc0Z+XM1FuQwVNizovR6kqxanL9EqikL9fDsUa1GgZrS/PUyY4NLrRYJevJQp0/NjqfkS9vMp
YTDQ1+0389dcdw95GihNiCILwXY0awT7HurnA/jDorwkjgFYIZjk6IZwGKU4s9qQ9h8vOSLKTHlM
SenBO0q2t1JrDfWWbvybt/Angid91j0YmFaw41nc44nw89X21KjS6ndvQvH9m6RGo45djFRP7y4j
may5QRfVPja+17cluZ6eRsqKzFp+dwtkhLeObv/Dki1ml6EVbY45WYq2R3K0tpllQ7VRGiqeF0tt
ajxkTGhZ1CFtmwu6yvyAE+GaCU/xalsxdNKNVgMA4Ozia2TvDVvd5QSGLm7b4Z/DYFHwjW5DMJv+
3ueb5VhSqPMAukUEhSNljC2UlM0DMX1CsWfTtDrqE7NPNje/yJy7XD7pwsxUxViSmQ7EK9u2mgL5
uRDdX2RPwbH8MnrEvomZUxCAeLeT4RdS1+BL2JvJAxD8OqOHyjWACglhOxPcZk+nrLNviHrEkyQl
vXiCo8abIFMFdJpFwc6NK47+tkUUZF6WnrOKoJDJF7pByOkfU/fP66Gdv32aSJtBM6WfprucQn1u
wh0r8ZGc4RKTXiDqhDUnnuW1lyxk9XBvnkPRaIB7G5AuOUjtBjjFSw/mX0Z1yILxep0rReAj2pTj
w/7cY7l9GeLqMI8gZNn6UhK9kxl/WzXxEqcYNw+AJcnN834w9fp4OqJA/296ZtSViX31rH9tWBZt
PWZhT5wuPqGwOd2I4fsQAjtAsNkFZF1bYYuouDEz/GJl5gfrVPhgxaXQyt6ko8jRoLni35medQ2X
FANO+Eq5Rp/YGxV0Kkllny1xaie0VvMJFCQvewpQl+PDbjyu9NzWoJ3QHDDZaIno3D+0dgZ7htsF
Le0gfuGSFGCAGOGWObjJuxi9nBwNVG/WPjL0lQE8KEmW/tquuJLTrP54fXnEDQ55KrnohYdv9kn8
1535CmgF0NbKhJ2rk66ImaRekQ45dZAXbeyb4hZRZW1nysP1lyxx2rVtsncLbaDnCWrFl5J/QC5A
ewzwM5bS9m8xsEhXWIlMRCFVwu+iSV/FOfN2ru9ckO1ZfXoWwROczFauO6V/PupSsb+uQhpD/VQ4
m+Ta4dreyY+ttoUAGBO+1NAI4rjtx9nOOYgNLccgPPtmFhPSBNFgBzXwis6Gsv+UsfsXzM+TsYzW
wp8lORICTxemxNbQWqAYGXZWvhU/vKsTPLXRFNkAdFSDBqI4EljzPlgBmfcViQgaZweWW6A4SerZ
Q1zNSsB+unpiJ8p/HEl08LPpDHmywtDoD6sCM053cVbnu9zvg1FO582a9+C4L1bwfoCS22LNhMao
xeQtMvF7OaDWdub3bnO6lUK/u5wm7ZEax03EeSlG1/NPa2PaAWEK7alK1xSUAhjGNlbt+9/PfL6g
ghqK7bowl9IbUweob3IEAdCEFRLUCGN3CAIHyEgR6pYAFVYUdScKaCaa40pZNK2LitHeHm7Tq7G0
Tk7yrOSZ/kB0isaB9TUmc7/HXHj40TGqRJEAKbuwhETHGGZbw6H1zsmPDHk2vPXYupRwRg89vnbM
aRNJVfURDxem63sAjL3+XfP6u9QFXRJEe3J9rlf7Fw1CPdtpKV58rFFoD7Xpi0InYqWnUPJJfa6t
U1d15cQ8C2wAMxhJL8zj9N48yaX9/eHuja8n2W6VLH2GQRi4LwtKoqasyy/k6p0+PaVWchxgv+3M
C2fCkbDAe/BjMU/FhAGWp+XqNfi63y/Sj3uStRp8uZKxJXAATgTOBc4XrdzFNc0YxjvhbZKwE6+E
cb/GrBriwkl3HcBvS13gIJyqO08tdsTKe6bqnOruNtiM2L1ibS3KI0l21aS0V3417H2zC2ys5yKv
6w/IArNQ+WrVqw36AYqUfxd1SDzEm/6RKWJ27sVu1OamaZ18Db1IS0noos8yzAzL93DouQ96Jo7s
B7ZJy4XbZam6XINLXNJ0VCK6sfts7pdyEyfGCwT0s2mC8Zoh7sN/kkMdRHH7bCD1TTppkDKpCo42
slmC9BK57e6Q4MPL2j9LsXV1Hj02/fj8GBfrzwNXjSzBwaRkQCAmbM4cewdaQajo2AfqW6UrRF4S
2ILc0q7gkGrDbyOy8wR3FbGV00fC6SXPa45uGcD9L/VtyQHLl75UqQ94y0vTxTegBgEJ9WuXkBLV
Aj2ViLy0MT7k6URQoZ/8xbnfsVl5tQISkN2pdPmPIEVaw8QPD3YsDZ9YGzoz5rbEAIVK0/7SlriK
21O1SypjpO4P2bCUztrruLmbHayKK3zKxd0qUbxJEZ2wlj+pRlTYT+E37yTLfgavED0+D4uILP/2
vfRqvQAUWT1U0eQBiDDVy/3242xP8FUSMy5YiKeRdi7+GrTEe+7vEbsWaqFlhyX4yevFbtL2e9Jr
KFZCjHui/oY5pf1JjzVYIoH2bXJyt3ONeTyrtDSj15qC9S8+FrMGZuG88f2nGddwR9FGjxjGtU1q
refOKjxPi/otzzaGqIlkpdh3+NS1+cJQpqmn9HVpvR3HK8kDlwt/I5qQmYLUICje5WJ5DNGoZ8Wp
5uS3YVnEDARN5tVZbuqPySfS7NAunwaHJAoDpAfN/VgIuXXTqEtFRd3LNtfqzk+Z2dFP5QiscAVk
ypDQ9jEETcJCIQ3X+gImF8dWPkP2f3/xvqgpJUGzQ69C84WSVRgJNxz3q3GEFXci+I+oODB+LVp7
U6OZhEr77sSqwUhUsF6ReGhghWE6/+nRrWhQMtIGdgx/4AOjUzxhA/M8rmrSCXXZAEKoKDIO1LiV
Ua4hDJgW+jJIqLRWwHr/0CnYhfPh+PnklRFtR+Bs3E75pvt+QGNmcDxJEzKSf7dR5KeFlTqxcs2L
/1LB06L+xJF51pNScnHTIi2pz1cEl982QnZ0exNJZKn35M5djZ3q3Y9S2cMh54AMJv++SL52Pa8s
qSYDnzG/rtK5hgiGNi7+qbQs92gCMe+oBkYlMjUZ0oqeUTkCVM0TIXUNWWs3OPM3xqMtHv4MPxdo
ovKjcYVmrOubn2hEJjzNTjyvUth7dYjhK3llLkQiMnXmZjMMFD5xyhwoZo+ZsFGV8BXECvf92p4c
TdQgfWIGT0y/x2vWoKi6XXbMds1so2G9N4D3IbTXHsUsemVdFlg57yXbZfN5SpxpKgfrjJTHAVR3
2NjW7d/msY7lHtWNeFoN2foyN8vf4dsoHbGVPY7YuVIqa4IdqM64i6y7rafWc+KZwqDqgF5YhU6q
1apaK8v6r6g/dga56RG2B4YcF9AJ0MfKsiLZBCP82EnTHGUIxyXLFCiGjW6eP3NG2zcMyU/laLCJ
Ry4N+JgRhxYq9uCCnsQVR7Dx+6yIri4Tj0qxuUj5P7pb/ITOAfS9X9+ijk+S1qLliejWdg3PbRc1
jcW3ccvsjniaTzQGQ5TzTIAx8QbSeSUMmYBLrzwYu3YMCEVM9XPxMtRWZMzH7AAy7dRGqDlQcUsl
jqzA2P2gZCHHxUXba1XSe8cPwTfk1s8VeND2E353nSsNRglDGgSiIyNwME1D/hw6bKdHUf6TVCsY
GTyC06yQzzt4fc9MccItJcG1PoZoafzSjd74QfbuNhfv1fEvbyJN/elnXdsCxTbRlaQnCmwn4g/+
tN3IIbMdP1pHyfO9d9sJVp+nwiYADMzQw4WcdbTRd2GA9Y23Cxlb7USHpEUdaTQU9wAESjs4KfG0
Mq5BhHRhRm0i9WpLo+9NPhsR6IMCw7UCPzv1yG01yH7+qk7AQ2lcWfVFrMty9FNr1uoWjSwScgKG
WTCYN/XilMZcDwW2i2O/kFNdrRlCP12k6cuI6cGH+3Cqpg9F/fz+Hul3gW1eQwioDt//3CWjxeoO
q9BGugPgqKP/LVVT9ci2sdsaqgwFNq4+MghGk1HZItGoDHTKpKWHCmoUX4pUIXYu/ap7AC/gj5pM
6TrunG3jz/lH7v4n6UWJHKDWWCdaSGAspJZVDDWCGOo2mkBIM6pZM8BpoWNeLB3IXYVulQbQv5Lw
ZlTqp0F6nwhm/b9jqWMZ75D3R4QtLo9PDBBnpE4zb9pznEA/OUVtviXosbxyrH7JU79/ZTE4lwpl
dblqI3hv6GloBma+mEBYYTgC20lRa4hmoYlEWrrMo0hvLitHW10GJyx9djSnCbQuM5Tb2CgTLjN3
HIgmK0JdKnuxn0ae0IEi3ijDs8zgIu9GDmLkLH+zhTyFykdZmACsrOsnQdbQpYowhxjvPJi8hRm8
2lDPhi5rpQgm/B7l/pqJt7VBQAK2JNUDD2jmxlMnHh7I1IgF9+xyF7ZznTxtvlvGiOHtueTlip68
yxeZM8qH7HFS1XSPO75IaSvc/mc0akMQkf2QiJl4TAFqMExZQKa/D1csJCRH3EdFd1nuPQVCKCyY
tTAonOqaWo3uzvf5PhJdOzOluBK+0Tf0Ncx4+PwHc9dVWu1WhtzOepqnbGzDp/wCtI6VCPbOwhqQ
he8YGsGd6QM2z+UBc2Aw+mZpt+YfFqb4PKdSRuPr3ZrP6qmHwOUR943IkfetWD55MZBmkzVM1BbV
aXDc2qMx42jshMGfD6TjLHDwGJPqzNNz5ES/y7VvtilP7dfEOpwyDKuO+9qq1LcJ+CZ6bf9yWNrr
NbnCbDPjr/skQCBuM8HrhxmOQKW9JWJ9hPZTyHd8KMaKLGpL+EK2qgKmMhlyGKdxY0tSWw9B5/8e
aTJkSffbqJog/IoRnz3KWH31LgqWlpQfD7GoKoF3z/jz+m1RjVwDJgcZ79FeRzwSh7Kxt1Cun0l+
ro/lTTYtGiCKL/JXShsQZFEEvRBKdawbYCog0uQwDASRsriYlrmi2Qt/lK+QcXmzWUCAx/awkJJf
71zB0V+onQBjJdW7sjc6n/nQ5zB04TaNJLg5u9pRQvPko/bN8HdTTim0QO1fttPXlT+NdlJQrCGt
GCu4mGJNgJQO5paRBMmcuwOKr77URs+cZzkVPo1ZORuOUUuHUmPnbzQGlyW7BX+MTEB5+CsQyJRh
r61385SRl0gIS+i7ATAZMuMfWRbQ8UQl65c9ICNhMwkayBkZ7L5+us5gfHSowJ6Mu5yaXF4AsEYq
/TGWzctll2B+H1//cN7+hnThzZqZeX+1kpc9wzUw8bKXBf6hGTUIry82KMkNVXR2fCpXiobWRb1f
GoKqTfj5XVnvynwgrtzcml7byMfYWPsuO4k74YsDvnwOdJbdy839Pk+aVfIJqKdEJU3x6USPNqIT
Ur8QOhypmVah/tfiYV7VKtciqbrFfw87WpezyVRLbB2sb1yOz5qeb/zfARL7lTT4IIapqAuNIPGd
Yc9ZGE9gypMWqklaDfSYghrg/MuG3O7sJnh4xt9VbuEChE+4QHp0Dsb/C/VOpVdQaV2ioJjAF+za
Gs79+tWmtioO3ovw9QI9XZTPTNGO9WFojdj8zNIuChWmtrj//dP55Q2opXmW0hgmZZGTYy15SMkz
4ehx2335qOO30lcsDhSWwzHiR6lMstw/gvYvo/ODY689zCBEwBaQGh0+5aaOKKmED3WKpCRcMxK/
a3TAfTEvlfxpc8A/WLO63WpaQrJOxM5xFsRivq3QhsCbX3R1Sq9ny9BEOfJ5oZjXAhe24srZDSWN
12sFN0BrPpUHxqOR9sK2NBR4r4qvo7UsNlrTCrSYoonB+wqhli82DCRXF1MgMCCafwvqvnthxyE9
plmk6ogn7LN/ZzNxQNYnTw+73b10YyhS+VMMF7LyU5z8Dd95EpA5uArEdQt3B/D9VaPyvtuEuU9l
Z5e76r6/sWx8t6OVH97OBuXiS1p2Pp6UWbofwzjwAbBFKEJK+WCzdgDWospPB8ldpGJsL+WwAQ5Y
7iiGglhOQsrxw62Fd7pgZ90VhlIcRDlPvyKTTNjKjABe2nEWTIfaK/AQvyELNvha603btWuYzGI2
M3TEbXOrqTprQ7HmVAMBeAiAu6oB1Eb2tUgtEavNdfo8zAuEkcX3DG6VbPkgPTrRun6Dmirs7IWd
wHbE+8PEzwEpel317bbDK+Q2WAPWyODpaSVkrbbG484vtojlJbJ1Ynzajci8EP+wU2upd5IC3HJh
uqvnD+Pzyy9m9tGyt7pHRLzUeieZA6z63W8dYGRewFo+lQUPN1K1SHxBZeeNo+ajPUHIB2hpXsxF
YosZNt3FsnEZY1R2BO2lpn6Nd0yJuxu7G6S29fqymNL2+yemyBgWxzfoon6r+i2Di6i8RxXlYofe
XzZ5Zmp6yF88FTN5Tg0hVVf1TdSU/X9JDVHlPViCIf5mIbBdQF4i5Ap9nM8v1ymM+W33lpvj40eW
KgtJ6YMhLokmdKaPDbO/HC0tc14HDCVaqwmRdJd7Md6j1FkxWaq6tcqKPiB3ekOSQ+lQJOERbv6I
fUBDr42X58N47vlGKV6OiNAQgNt/KJsR2VWqsD5a7jzKh26oG7xEQZQ3aN65BoqrmdSyAlviE/vu
6tlre7BHmTRIzX/+MMJpx8y9JPYW3hY+y72PCfpcBx3Oad6ygSK8guMz1sjWuA3b38swjeOClaac
wU0WrZQ3AIufM7aL+WFzy7fbAE500xevBgrjkcIARJKVzsVP58v2f6A24kh/tNJtt8S9UAYBXUoO
THSKmUOzKlRhD0hZYuKEL4AnoEUPp+Fp2AmRxtOebSM0EL+qfxl54cnzf0H7IXvvJY0Bz9m1Ch0V
Lmrk1gUmuXV2HzcOA7HydthzYdldpGqiLmPX7MhT2R4ur6//a2PBRrGqOgMyrenXEaTVXAW046Xe
FvtGxHAgbrGOgB9noJxGEA5+R5CyT+ezLg92TRTOuWMnrMf5zXe3KEDvLWKMAetrxAoY+8wfG1tc
uI8BXjc+MWygPesSEBJv22H3Ef9BllDjG/vasZKTTaybaEJ1c6xXurdVm9qUmBdI6B/DINkembui
PN7IPOqlVunYqWFvVTw60sH1K3z1z2W7xfeJpB9w5XqgNp02XrtE+2PJdcGhuhurP/3dbKn0gCJf
fiTT4k2qaDRenmmCS/xx3zFI6qebuZ4jkLmK8UzzArlrP3YhKb6ECfFrEwr7oISiEPSmcTINr3rx
LqR+5GTzX31gtRnEXdUHItPAtuj/UoxS0JZ2YdMqhrLvMxuFNuGAc25Qgbh71/GcZeiLkVCivSfY
jEHobRHcJejoPmuxveK3VFiyi+eq69noJvLqfpokPoS01x4s2R5NsZTVRysU6r+7a1yxq78nDFzl
tY7I8v5Cjmzm5gD2eWVNwwWQnvvkRSr5weDylDM80msjPCbqPGXmKX1J6WexvWSfUSO7sFuKmoBr
uXMXyM1nDLax3JlFmaNxbNbqKjkgHAJjnBqtklGCVb46/q0Xwd1R5IWCtr2ajCHsU/4Cl7mTIq+x
L2bQB4Z3s8qoA9N/fuUpYlAw+vY+q/DYnbjrFpfCtEqmTL2G6uSsYhrgHul/f+QeDI1hsIrj3hCl
+9C2UuploLvYD0sB31laQzr52j81ccZRJyaJZHBcT+9oq7AufphuwGOFdAVSPAAIm7+uY/qgUaP8
fnUWCiVkKvflkF88WfAkFEaECSGyyuMrLcKt6tIN6GVj4zhG2QS1ZqTAdkKDrPCyQMHMRpRKMRev
q/jcP6ImAdO9cJ3Yyy/tLI5hp9KpIb31ZyN7O01Am2zHEQ42MLsS4UaS48B70cTcvNQh6dCxLqL6
8F8X3yXidw2raHure+xt6nhQu9HaZzzpVYf0Chun19cX3cXlLIVIlCRu1tL2uVRHHMTG9KZN08lY
D+pGlJdjHbF/3TY5s3nvbvmvRFIFAusEpcnufSckCkDMEpaWYJ+irr77Jn6gDeGD8SwW3IDN+awk
aKtuH97oI0/Q76alqKWBZLGu/80SiQ5O8gVHiskQ/+ATktN6COUYw/ak9VWO2Tl3ux2rBlfd+JrB
sZQqSKWvdTGqyMLy9QqnUQe5aT5yzad4yVm2MX0swikZxWDhLXvsoDUv/KilI0j4EuvGrYLidSMG
xfc75UfgdQ2NkQ9YWtFKI9rJrG6eXnQEch8LV25n5SzANiXlcJimzxWw5Xw6Mzz18Mj87iyzEW39
tH+VudZCfFrNtcTrUGgkBgt1YiSaFb6dhq8nhFGZ+bf7vh28khLIamTXc7VHAVmI0h/Xj8GWeoVJ
tNZ6TBtc1D3bWAQPdNr/UsGZXfuBdMdbAe3pHrDFcquGwi9yG1rbTkxoJmHyr5gUeRj8jtjAZiV0
sBiy3Qg5AUK/EMhqZ656o58r9f/7SBQLNVx0ApvRRvYAmcZYg5JV4GUxUJJjmQVapzsf4et9L7OX
sIbqhkd0XeOuypFM2sr6diw0SHbtVn0XjE3jzrZ3Z2rFVw7jNrwrFSxw8J1kZ0xzA6h1JKyWgabM
gVgVnjYg6hkNYlCXbNYX4ELSWu1pI3WWly9Ua1S4ksloxZDxzsTKhMiBGaiJ9WkmpAY6Sy4+0KXy
oosJwF32mKmyyivJfn8W9g+wtC/Pe6IVaYarwzzU/NvpupWexu7MgXOLUpFZ4JNnNFn3FY+TX5ve
1Dgs58tpmjUXPah9Xo9HOcfvtq5YlrEEjzfFEFfqVw3mNKYFEOhhXCwm+wPkSBx60JClNK2T78ul
DNJHRDAmXIXUpNRer0EGvJR4ynQGISDw0z63UG77oPVmu+iBQwcwku+oM/T4i+wQGCC4cu3f3cOn
bxDpQReQ0DzpExWdDLeY+0W4laSELEh6L31/zmoGzGXUUe0tGvGX78Qcs1tlxrjV+APD+lJQ4Oan
bMx3aM5om7vkQZWjs1LhrmoEMKbNja1PLNK8i6LgwUcwgjBqOf0a8r0QdSNfpBUAro85aXlFhFo3
BKgaeMamh5kzO53zDOeILtDvrW1MAxi/4uszMpPv5cQKqvOJAzrNu6xf0eHxkOp2frnzRPag6k1P
S6uoKesBr8FaDe92HwTjsMQlaX3FQc4+oVWcr+8Z4CeqiJ+u8+VIAAYYIRLJwaRE0Gzx39OGl4w6
4Igz3/TQzvmN7N5mhMQK03CdI602S1317w1OhbENNTUKMJpzlcF9uFBsAYzxfHLcwiMjifOHPp7y
CH1IMzC8p2YZIf3W1yhYiIZv2gCPaZoujBwD1xKTL8O52hamhamcPQZ+ot5CQff0UmmYdSyX2+2u
oNb7SM7zUcd2eVhuoULdjqCztKJWjrbKL1iVcp1W+Ld2Wc9HoJdCiE4u3nQT/XBai6SoxrLnAgLT
sr6gaJmLnjxDYjXmq7lQtyRDtKRE5oRqZ+yydIRq5d3SkQ3RHGn5lNDEjwliD0eGxikPaATLI5KG
lcJBjWEXQHFJvPfBQEdJwGElQoB5oAUD8rKASlOyti9Xah1qv3ySo2qlu8kcaG+hVx4HR28FwHLm
yUzV7LqKwCwmY0ZVonyeO+jhQn3pa+QZphYAO4iCdV6MUJnj9kNjLyiMDi288AH417kLTDIAKSfp
Jvhq2TdpfMiE+3nR4ZgXooepxBj2UJ4mIh7bMXDWfcqMSX25dH9jcExV4CEzDkvwWjrr4TfC6uZX
SdCq51WkG/Zbo/nlqKzPqSSFNVoJtniz6oiZlYfyLbOazGRuyz8lnLngAzI8RI0hgpTNtgoc0C6G
OQbLHWAlPQcuOQhGDP/P01Tk84tjden1pK9xo1AG8o2Oz/DhncCU2cP1W+CzsYD+crQLeqr7qiEj
7Ry6My2qIiIwYhtNjX1Z/aAXe4lSi1rVnLOeC9NJQJ8/crmlKoi44XYZ2fOHs7BOe/0SX8zSRoMV
JcxZGIY3fVEyzIJI6RA3pamMm4E2R4EU57fSJtMqAD7bsqGeKI4u+jHWrDb6XcVqM3scD2ylOIa/
7EV3LqUeHHf7MOYr/IyETvE1p9v1mXJTCwxTtxCbDRU2yhd3o61mFSwhEKPAaz2Zi/KcG8dOm3fG
Ac0Vvk2fd8AJ00FIwqIvgtWT6h3irsfX2fSGSXFMmuvrKaYnUdX0fbJd3sYjUXrB2e5thcQOTLCm
ub7wXzbMij+gKgt+xy9LfF0Mo9aQ5Wdp6H9KEtUZO1gaVBRExrlQYHDs3WXlWXimarIeFSiPcE/n
2QqCDqNKVUX7sMR7BrzlgkVBJ3us3rQyR60nMBzh9cQRCSrBSF4fzKvh6frJOrWO0ELxsOV94can
t68HP+yI2On3SZe+k/QCEm8+JOIsv0QhMt9wMPi6h8/mSCXkLK3nUJJ4kjvFc95Wd3e952RK6Xcp
3rrbB2vpyRcW7FOhOg0OawCZIXBPNkoKFAEEIMBGfXJWSF0R4NDxFN2dkYdaO8wqZE7sA4MW6i5o
TsNHrU4bmosn8/sZ68tDfOj8Vf1Sd1Bu8chW6EmlyoZ7IdTbZ7TPA7sUUwPO5BMEVFw/IlFNEvJZ
Pi5oc61UB8mWEYNfrT8/tc8kRErBq0A9rRlN/bqh6UEjeZJN7pxO7wbTWrQVY7+uw2eNaP6DjeYY
wOLad/jUydHlXf9vK3jEzk5QFlUmMkOa0LDWCb+RxTKwBuUSPHrgCb/rlaBb8r4sRWcVmX2C/StN
5oRrSTNw+J88jgHRbexCLAL14JyIRQMypIakqsShOTstNkB7w5UM12HV7WCyg7wEGuF1zAU145Fr
he8PM+bY7eX/7Bpv9EVkzKbz6ExIUyfEtt+BX7fIBZ2MB1GDpcBL72+P69h8ppQXxONAJN196ouy
0aHtaCagNixwHQxrD5ZwXvQtywWoT/SW3z3AwVQxWZcDWvO79uGX2HANh2wrUroqC9hmu3F1m0Jp
9XBvAvi4XOSaWPr3jyWWhwpqANQjNuPyzQzFwg5/kQ6bO8riu1GjiI5QYYn9TahCMPV/m2sfxINc
VMO7WfDeFInZ78MZfBTOnr6nrOImuBwX4jetindb3WSP3WUwL2EAJp2NeeIXO16CkD8U/HaDQAOz
ogCdfYA/vb1oliX1qdA6f9xzlRaNwo5AC9g/kfEHHvDSluYw8NnBAAkqk2bU+ivCINVAFYeVPzbP
o4rcdTzX4DiW/AsG02yFYbpiP45RuljDrTVpZdM2ljFoSa94lRvQCT7d0+2tMZ2PGsLuOdAgXQiQ
L8x8cBMqg+ZEJ1MbwnzJvBm7jYsgkMHHUnvHuQcOEypc5aD8MGnqhaWpO1xahS1qwq14yfBeHGYZ
d7qV8xy1BWhV2LforVP3kUavO9YTLxcKqhxyWGSgGjNcvUeUVnwzReuK/W6HNaAqroytuHk4mpzj
YJkfiv3wV1gjN0m4u97xtwZcl4EcKorRZ/Dhvl+UyHqD4plor1Hoo8yu9HFz6gnXw8AidzhV9dj2
4MriwtDrzq8iY8q1kxeHpr4tR3i0lYtAWLPFJF0e0GU1rpIT/XwCvz7NTLcH0cVmNb1ofEulFYZT
yCTLErqTNo3OVAukaXkV2ZkWeI3gFzCwhZ4fxp3wM8Rz9hUi+qNnS4EnJMf3kcphQQfN4WlSauId
UXpwaWMYmmFyW5ontFrQKs7GI2yBZ7in/o0vvrnB1yFnxuSeSv9oCrd1ezQas3cegIhT6MdSzHwY
pquZ11+yNFP0ws+8DCzkOX9W59hoUFBRFLe/L4wUKlJTvpCqROZVFgm9H/eqCChFM7UJ1z94nnEb
353JTKbU2bC6dG1b9hulQHEpbfU0wa0cqxqteMgFgTsQ03uBGoJinejhTvH7LH6XejUsNsKzg13m
tZ1pytRKIwaGUn0mSvTgXgi1LJVSzVB/QmUuWJ3UyersUKcXM6u1uwmb+yBffvtJMD4XVgKkfald
FktTsN29LzPpmW/Z2eTTUAbyaRA7QlQkl3J+lPx+MDwigcptij7jNkSEpJgE8Zwvp8l5+cBbF8RV
nBiWlogvl//VQoPhkpDBVvrlxd/P71jxQ1UqT2zjWEgKpmGxi1m6jiTUG6BZmS77e4/vuQzH2WWE
RVlDk3kq+ra9HEGT4Co78WUt9s7zlOu5jBsB3T1O7h1LKn/2gSftGT4hfAvjxkPWC+92LOS8idNL
unfNfgmiUz5bqRzgch5N/5HLUL5tENGg+QijAPv+KqXozi9hV29f638rVG42ZCQh5i0E7sXUz0AB
XbeW3u+W9ERQMIrW+FzywrdEL75ZQlsysByhKvbwyit1Yf1OZzWzDBHvPxw6SfUgICXnn/7u9puQ
aOIZE7lRTrqpiAAZXqc7kI++SFVGb42k0Fgknbh/AoUNE8prfiodB58tqFxRV9Dj+UO3kOHbTf3b
ZQK07JGqWdWoZpMBjMFrYlPq5YRZF5Nhsu1i08c/3CyjsmFOET1ls11BqdjwAjp3m/P5P/neWiI7
MHWJQiQuipI8mrst+LyL9ch2fV1j0QBCeBzTD8YVSJcZ1niXuEfwOGlyDamyFk9kxql1SYBTrxlT
QqWzMqEirIyiS3NpC4VGOG2YeZdEUw84x91xWvxN/X8RJQmhPqqpEuXHJPLT8QRvI/X1TcnVdFeK
g70WVVUnL9Qg5yEQZB64KX76QOglIkBDlcTLbCPcy/fLxA3zwjFBl+0qyFi4ukEsObVbfiofYVZz
a5ROpexwCAkGmoy5F8iLfhtjlT9dS+uKR91JoYIq2mJwrvvcldibTg2N8IBg4hwAj6O/9E7W55si
N/KRZF9jtYiRHgT/da1/OAqz8e08RhYqPOyYeZjfG47DJ57X/ze+C/KKNO1wlsL1pZL88quEp3HI
no0XTuLqCSYKfNjDtTFdeDWTdo6looEAfQXidRdp2GN4c0uJPQg0+KToEsHVmDChq1GTdPdyfb3W
yl+6Ua4+lCvlEp30zy23iUzYnkJLPbpAKwebg1rkxgHnf937CUFxVZxzSZfvDQiIYmPmJ2IxMCqs
ys0rHf0gbZ/G7cI4lxOBybLHi8tStw6GR9B9Yg21Ly9evUhp9WihBjKtOVb2uGr9PYP6WYzrtZoa
cgAvQ76NKL58iCnzBtFB1aEWvat0/ekCwXZBcPUWj1mmwAnEhl2ytfml9oJk7WaaGnrCr7Lq0PPK
4SmI7P+NRXn2yVHzYXjBWFRpmG3JdedIiBj3TTrlPx8ayAZICcGzFoZdT8PPyZkudKpohYRj/1Ey
jFH9BZExQ6J/wdWumKUy0y46Mr3xk/L7IUwPcYwTWkXd0YdHVNOMcfCZerYApYGuytVgYeXrKopA
9ARRFePECZtkStB7nJaJUQhos/FcRo+C8RelM5TwlkG2WmyCMifSvNs6LBXkm2D1a1NobEDgHsp4
jaeEx+Em0DiT+qMXg2ye/qsek4OQp99ecFxyxGd1h7Q+4sIhAJ86BHpYflqukkLgnwYbr+hipb8s
1dFjWEvCXYDO+HUgfJqX/mUMF7a9eH95iWdxHdJQTHuQ8G8nqMuuI8pVLQkzadaIqfXZvKQyZhUr
ORVVc40oNi2Z5y5QJyk5eXQyrL3/J7JR+V5ca3S1dwOZy8o44KefDCZgHkSJg24g2ywtgv71kZFu
Ok9HqWcWiixr7iTh89u5cWNhPFyDKhfJUgPUsNdOGQRey9Mook/cfmx+AsLMRGQ4/7xCXqMs+erW
QdBjiXFggMgvSFfp0kO7ri8TWqAbN74FcV1MUCZKr7WADztoDEdVFYsJeX/35IVx2tOQKu52pVXe
i6o+uH/cI05cfxRjIWj+w9ugkI5kdhWNLIgYNjHfqdoZl/Z4mqEa0dfHJWJGR8J4bWRw9nLhg7RO
fMFLh+4MTC/R5ck3lfAUk1KvlDohKXjWWS2CFAu1zN7fR7RAM3IFmuPQvOWn5FutDNiqwd3RTDsS
hfx5uunp2vlnWf1KXH3Pazs+tyMbsiju8hb3yqhMnf/4hhjdpdx1ySAdRX/vAI6lG8TjjuvtQixJ
vE18TEtBrig8M2k1/M1n9jOWWSKtzlThcT+BTsqyrIyUNrVVPiBSqc0l2zSIutCQekfwhKQC40gq
dPMsU8yZ7KoakRKLvwKU2W69xRg2AeVkRX8G6L4HrrNgNDlgDzRj06qEk1JcyOgfGxybP99Zzfba
xR0QB26c3xPcSwVfHLtGf6ioWuCORIRk6nP39IOLFI7DhFRqJwierM+4T/dyom9UZLUlzT0f45kZ
QZfQGQpZx/rmWH3Htx4fsa/VBceWg7qSAZ1lGQinitJWRP/Z1/P8jxCXmnB/p03ScZ14TXhTmMpb
qtt7nrlKaK/CJsiYcClBXV89eV+ZZXeLSRB0ixaIQOb6W8CFoOUQ9M3/Wk+hZdQsUCZ/2xCb9jGw
ld8AXmyyqXP5DbvEYi+C7y5MUt74zM+uIRFW0q2ltqV2z7nggMYOAKsDvZe4qYElI2c1DWLUXaxr
7upOuwZDy6KJtBJUMTE8HPpV6VGbANTNkTKh1W1zrpjdn/X5bmLlKSkqE/PGuZK+qr7cUzoBrDMo
1b9cpfR15uKTiZwsbSWinc4xvh7CYQ214v6zh0hoOhkb581UIg1/QsvGK2+XGiezZ07cA2MOFQvG
TvxR3iyiCmWsv2t5ArKjg2IqQH5Ngs8mIpXRa3fjBAWuWKo0sv25xaCIncjP1p00bNPgPV+MgIiP
2ilstbKF0QcLQFSjP9Uk6GudKqo3slw7kfpqqlg6PZPSk2cfIhvxS+z8BrAmSSO9pn3VN9CwVIX5
ttcYKksBzccyL31FN51jL9DvRYifowazdD7L/KCvOdDnlwLDdnbNGG8mJnBxO+gUhqDPebN6Rssq
NA184KN3iqGgec1cYj2XTXgbuq9RrGMB2jfJ8ekZpFhhdXFUapyXWiUtM9xJv63zO4OjDkR1+GVZ
p+//8DOdSzNPZpQk+gGqA8xQ7+ZUkUieEBmUwfupOIdpd7dOd8KmjxPYYZqnl2lNU86RX6wtlREl
++GmGH7kWZdzDyKXJGJNsaHuO7EtEuJfjATIfbeUX2qlcPBHY2fA06jo1n9t613XSrQAUqtHmMT6
XYDzx9ywuXcXEYPlMJOfQ3IRBAa5/rLBFVfQ+l/00WcBHTS72+tzg5TAb+nzibNsQP7CJKX0Efih
gu5n1usJ4wulGG99VRmBJVK9RVz/cTIAJhrPM7vNUGAOu10Xn+3QcUpyvgvp6wXw10L0ivyfFNL2
ALTspltB/lqgGmEWeoMOYpK6BQLJcLRhfa6/WRLZvjI0QnW/8C6v16OKPZNN8RjD5LZXgk6bUW2n
GNc+nXL8njQwGp0CX7z/LgvxRHIZlZ7wocMeBvk9obrm/DcgUVQhuJ2UOP4ZeNCwYYEBdzthedjH
aYUQpXKjoe4AbYNGA4UnumB97wAYFAgdvupANQNQk3YSyUBkk1GBD97bVUp7c+SXmFaA84VBuFGT
3HY9x0l67MWEnwO3dY0xtw3cdjV+WEge29R54jHFjMf8lbx4vokagzkbEz+Uv1z0/xaSP8Q00dT0
i7bKnHgtRhdoJk939MSfJVdie75cPSDF2d9fT9UO16WKKhtF959kf2oi8vsornAFTjgov5cQ4MgJ
vmge6iQNC6wsAyMQDcQ90FdCSpgq4qDTcs6PUHh3kgs5fQg+nelKyi3DfOcExqUSwlh5kXTwWfYF
I4sgDEIoEEk9TZNMpidKdWP093DFMqtAkgRF9Sve/uJNfbUa95MPgCPberIrberabUtabnDw2tdK
vkiM0wditZjuCdzR9Is1JmooLSqYJZpN/ucrh/Ez9hoHI4amymnY1DklW7N4d7JwuPCeLzkKGZs1
eHMUE3bmiGgJAKJf7Z4ctSIYBZbZQq2UaRcv1RKLP35nscQ9jt05m1ErSn8303Umz5xjXFcVnPpv
lrjBLaUKGNgH/pGQtn1OXkLXxv4yXCLp3XQ8JqEAlg5y6pfXIAgbEFl38FYsWNwQYA737Wr6PHQ/
7GfjmWmHEyh5KoI9iFSHcy7dJ/hysnCgBM/59Cr4y4uE4zFhkNgrKMfBGHUkpu2BORmJR56DLbWB
C+4JrL5KndSIThWMuebftUH4LR/g1CkAHDJ1ZgF5jKOQOKYgqXb3ompjSacNPa038TTANEDPuJ6J
r8U3VDtOoUpbqkkt6fUFcl++Dx5jn4zxAxFxyVj0J1oQ6SnVip8JMYZnzXp08Ju7p6jjt+i12fdw
tN9ArIxDlhcuy/aNVlqEpvS7QEA5oo3Zi9UjG2PPdg4xplfmZ5vAswzF6RBbop7xFbZgGKoyt25l
5LLTZDN5ZPyd2eohQ8uiy/vkHToZ0QScBMv5chcuiCCosi1pP6ARHASnKCY3kU0e75rLeRguv4UW
JSFCudJGj7PP2FGA89EXB2X+t1olur+P4lLwxomShAR2QQWJdUAA8qKRmuTHpaANzSOYcancAbo8
Mrn9r/PFT4E73xQthOzNwlPZ2KegwwmnWbkDFpKW4l2TJCqEChjIkKBXTaKVV39aVjgbwKBClr3D
ccY776oF3M8QSLLqg9q3TGLuTP9Qg/XyJhmCFjmYm7KI1r29Xin9Ndio8RTH2o6Jw9SYaHhVkmYB
z/tDWVvpd0+9hwN2S7OsxjYihkibpsLHW9rveFUuIAg72akiRcvgEuOg3//y+OoqICnZO8rvcwdX
6XsT/e1xqsp1OngaE+N+VaYRTBIxuaHbjk8EI1RoDdZ0s7z84Chj1mN5pcpTCalifxwnDhJp7Hgh
N3ISwM95TqNZnRLw9YE/KHqMxHTh7VMpEbB109KYbfAIr7Gr4AbBgFO8b42l8RAVEgnzVKksj585
m1Te+XtfR98nzCsaAJlPdn5Qyir5Y0QKo2cYkH1ecDvqbyVNLM3Wnxct8wOF1WStp9t0wiyAtHWH
XdEclaNc3p0+t0LqvhlLH805XpNuExmjx1VfidI0JfX02iJ7D753JJKr67lazYtuZOIlhDgn7msF
v93EfzSsyz2Yw+GwNSaqaX8OuRxrRT9wMctd97z0s7l4a4yocgqz6MoBc8hOVUmRYLw6dfN/MrY3
Qh/KXOPWWZu8NXnyNTQ0fc/x7fHT/9ZXIRYqZHccHLyE+JPKyrHViXq4HUaMD7cY1+e2J7/NO4a+
qCauF+agOb04ueZgaJZ5HdmbRREk1axWe4cJHCLFLZVI5N2CdC5dNHLafGytJhvMGKZeoEtuDbRR
N6Up5G3N8RHBNP2dqtmDxZIJtkM3eTPOwylbpfQuWBVBjjJGkCQgacQbe4iK0DbJEJ9oQHbligwL
USx8x7jMQg9+NU4MTMQ7ZPNL7Rgsii30J0antYewieiDRm8VkuyXnqJPMHCpZ7asfTzjcz6mbjc9
qC97SDX65UxDmrkqhMAtIAkUZw1pbQgPEX1kzoidysLcNs3Cd0ErY4b12gYeKsPMZKhxc4DRNYqg
EvJTZWtphM8iD5AzYgAcHdR/gqqKn0o5dcxyt51bbfDLD58j7e9tWRrws7AhYyo2CJSpAk/svE+t
7SgE9IVyuGD/usfDjm/paWrW2mFmy2oifWSD/ywmUS/jGBjUSgDxdjqGmzoqz4vMTuJ7zccpEPsI
Op4BB3BlsTywyFURmERAZlKXY4jMZ42czt6jmVRDnW9i43GSUnswVlltkv4WYAzu1g5Khpl2cViD
nSrEz1Ch5Et6yHWmiI7CU4oUPTvxQp1yVyAGxIh2L9HgldtHgtglus5aumM9eW76k5I4Aa77XRCq
ueFvwHILdqgjytGMVCc1oPPkr+ovTIBTuvb6/ZVryfFxzfM9rm2y6KaksY/c71Qi4nKW3+ZTk7X5
4PEVCTCHcz0fOTEpc1qwohY7NfmiSRoToO4O1YTHKUrhpGqlJZnXg1tPCCawF1GhRGkwHbZ7dA80
DQkNKl4d84FW59CwoRASg571CNtuJnH/Sr7dUvVMcvGboI+xt7DQjP5+P3zIlkToPVogJVaKTVQm
UxE4kQGn05KIjG375BqyLzXjUSlwgLpTMDUmmnkAb7RDI0aByJ/BghqLUNrSt5GZ3Ah4u9nkKhCw
avwYDombJujNvZky06Zdh+TbfC1x+Rr1+IDteVIO3q2XjQskRQDAoUImyjAdaAcZgPnAyRkopEim
TwsOc65IQKugpotwNGK/UDC+c5sDbXZj7RnXGNr+2iNSvlgFJwPnhU9XlTnvW27gWNV2NIacLO7b
n4hoNwevy2dUdi864fiQ8yCOW7Uo+my2qobou13r0MpWZJc+Sg5ZYAcrwry01rqF7x4WYLgwijEY
zyGLbpWqwHDfu1quTQAF8rCtShDJp1LiL/X26Gv3b9KPvep/RSxkibflmsnhAWSQdJLw3wElpKgl
m8agOhdqOHd7+bjWgymaDbRfWLRgy8ykcLqVddcRexwCBxrk6hWWae1HY9g9T8VQ5xrXouIAGYCM
9D1HDF2tXa8Ioa1pUKOwsQ6zAvQ/68F+Ni0hPMgcvKAospR6YfnbVIb8HmFadwolSUZDtsu4mkS8
C/RRGFHsGvLLl/ojOwK8+ON92THdZTyEaDagx+qmcKcOEM0RHD4IJx7owkuKhZ3mzFN9Va3KUm+d
Nbl+M7HinUZTeVDjR0mo10V/Bq471hA+cWmKlXhhgEKmOfVSZ4KlHcKyqXwpDAYjqBFo0V3a7uZF
ie6Vk6lnsSUSo+tDIPHYQx3ClGO4wJBvEdr2HSQR16CGcPZIX+On30Tg/8soTWA/dLdO1x/KH1jq
TyOQ85vdGt4CPIXR4vDR/NO9S23265tTN8dUO6R7d16+xJUfv5Uz7fQMHpod+sVXyoHPUFVkR+NW
expFITjWO1nsrWIa/FLakYtnGZseT2X74X+FcE36X3T5yx3w2tivf4iLkxpb0g3iFxphWUom10tw
y1/gIVdUEqaZZjJVIkFR4jSFXNghQJ0XwRerBOxdtwk7xMIG7qS3jTLtJJBtPKXgBsZtm/WtJlWr
AYuCOxpkiXqZKdUv2Xzjy9AOZSM2jCjFJMmR4/P75jGz1mwITfGFbpbpsvwlyV58vuo20iRj0sdy
+B/hINCvp01/KOds9Aq4ZqLV5NJNlJmmTzoWKwvBg+o647J2Gp+Drt5urgR6dPVdRdfSQJHo1SC1
kjO0STx3JEIBraQW3kmsQqLmkP1bV2p78cBMCan9kk4Yb/t+KCspqZy3QOoYLTnaY4/sXNMfobR9
BoYHXiQAhT8PJT3aWuwmafEFLuXRwcQixI39krlOp70OLprC5/H1469k9ODy/2E2eUQ4O5kxESFZ
3C1NWCus7rndVxfdvePvUB/AXHtB6jNU5wt0ccamyyZEKPU3MswC3S2KzqG1nqW7uHHhuNbQK3Bb
DYVwqmb+USKls0s5fnBwTdCawhokV6uKdxqPmdf84GtCWgdi4zXSgazUO07HgjmW7FCFuOLh+vUA
QWxmxNU9mbwxBS18zXQye1wpJGXrkZy8LDJnwC7JsPMgxVaTOL/ruEFc/ZkRUE00sJZ9D/Pbp1F3
t9V6HE7TLv0Gswf8xIA+am5hyKHgSZOLBrWfES5WouH7EUJvM/UPnHFQwDy1K7SNe8qiSSGKETCa
c/oeh/hkO7019YXaRjZIXG9bPzgZg3OFwsUzooMFwKZHnHn3ZjVB2cGXJ+aEF+5NOozSFxcLoJ/N
mb8vwSOQqzFam2iUsm96n/GLaEQTQjEy7YyMIayj2CsNYVOrPYqJSGlGntCl7mNAWQt+vE5sFCzi
JzALuTv2mj3wQpLahRhQ/bxHtXBSgCkmZPafSxld9krNPkXnzyjvDVzgVA+ClZ/1klNru2P8EcZI
HuvdPt9aqTt2xq3kw82A5ePJPNihvn2TemRZbe0uZvcIWFt+GdGzYCJVHRIz9M0P+IAH8mQk0Vlb
wWmFeqz5CoFBS3cGl4QKXqDEli8idKQDT5ml06wsaa9PInDkZZJC3K/jwqU8+RbEgPx/2ERmvFuM
Gsi/S3duETt8TQWdfaRRT2wekq3YTl9bXGH3THsCpFzJ11cHWvYQPu4wpkrXavJN9OzTMaDvPCvx
rvm7ZTXpmJ79Q8QjGqhG9cJ+f8H17L7UzrrTZ1d/6Q6oymSf6NtBb2vEezgpVPOVAc5Nn7JtRWf7
YfRxPKuOHh5rncNH7iOkzTspncjtYHAjrYXoVfu7wW2OKuPQVmXytKCS2cdSVjNjhKQkvcDE0zlx
eu/LiM4/8VwuljwA0OcsGHfa3lt1XSaGoQzvaFwoPZIpCnCrbP6d8klX7lM5fLdnxD94YwLqRbtX
6+t18ykJO79jXkc+5H8BNFdU/w9Hzdp5X3V08KREQqjvqDev2CWGx+vZfM90KBITvP8d+RiyF/kG
d6X3HsUPZa2P2EiDZecGQrPQkTmEQiCrkpFgRrtyTBQaOO5BiWKAlV0QMMbDGB2cvogonVzSoc/A
w2ioo7D+GDC+JrtLcefajLpK3ieeTy8TSIflykknTnHZuHAtSQkpnmJlk6KOLvLa/lMdOlFk0ayK
bMo2sEhROx/DtEsTC4paT50OlgKUf9IDy8XFkMp8yChft0unZPyVuqEStAGshKREtIbrdZq4FgBu
gNTSVCErJOEuhFA+VmcpIRmD/TW84/cpBvUvACqSKUlptNvauFqrBAk6OyVrJqpG801/wDS8Emyg
qm77+DoauIi2GXT00570Zdzzk/5hPSHgcQu2roRwZkjhaNU77xcS6My/1XupsBaoCoR/SGgRZKDf
M7NC1p20vHQ1hGd74uBORc3Gmdz/0UjCdv6OI00A/7wBOtKXk6jsUJommKRNFgl86eTFJv9HuLGt
h8cu2vvXNPE9A0GHr6caWjF3Fv8QWR7XZmhG9+ow6vh5CLv8tA7aWu8AhGHc+tUDkxnlKt9Gp70I
6mzLD9AsYtwQUKO+LZERg7GgWZW1WNd40jxYbWvq+kzDbvIAbEZYzanTMnyrUpdVrU9H+TV4iy9L
qTCD0Xs0qRrfjex+IqPqC8FDEOIBJPsUw4J8sv0dYPOs9cEV/Ne0cQfSNElzRlLRySo58S8pydOo
7itpST99w7ZcKMykQD89r9td01RW0f1WT8zRD9InUvseSQ0v84szsP+/9tGwjkQ17eEq5uqoKgeH
/stzPXXfMyNJxoqKehUfYTkg3LEyOjvG4J4pKVg7WHtOvzM1xJq3a7riCKbRDV0gA0Zae8O/cCV7
c0i1lkg2oK596pAXsQn0Hf7nTcnPUP6uaeMRCKolSKrDUUtDrd3/8k19CCDDoHBVy+s8b7kA9Jhx
6XqhscNcnbMK5Ccd96wEUahtqzYTTAkvO4QD9+WfuI/mO8EYisfx7HynQY86K5k9ISrIO68egtuz
ki1ZkX1JJ/S4GjZK34obdHt9IyAS9C/4aHUY/vDW+KFD+y224d/cYD60bMx+9W7AxOvIxOnO/4iK
OXpYBrxe/VN2zynG0Rsd7vERbo6EyEP4C1dry6gcHlVHKd+xBHXgzXJTxu2Vl37RW0q0X89cruSi
XNiOqP1UwldvAV05591hH9KXEbDtXAM37yec3VGXGYktwoWMzPC7/JyXWpzaUWs5XI4dYb721kO8
rUtte3Bv2GNut1MLW4xT7e3ak2UxkC337jlxMmXq28evBHH7E7qblFyXAYTbZ/VdzstwMz63prIf
v/ise0xq4eUUn0xc92Y9cJhRJkhiaT1fq0RyeFSwhHClVzbLTRAga8fmwpYwKKzbZmgxx2dnW6Rz
HNI2rWFEW3rBhYkT0u9QNCofKs/BinyTtFTsw+a2L+22r+g9xvsUnqQqsATHa+TW6SvsnD8XQxrj
v+Iy2jsi6j+jdXBZyvoF2KBXtxeTKwxqR82OK8yfDbgWIZJ239g7ZvscBw6L8CCDTW0Iho9Vf9dR
cclszpG5jD72Eac+8uC+toyCoPfixVvCCXG9wkCkSxXEDtYlxItlT7kpOUe4w/+5Uqyj4LXpfVQc
QuvK5t6r2Uc8a9N6MPn+G5OH/uCfKJN5Na7A7LyP+uVFWIvHRZ45AhG2Cs8ivVjCLAtfjs3WCIIZ
0DqP8BVMnSl4e+YztrY5AY12VY9MO3gUQUf6KjYyNCi+IvJGEJiSrnJV9Y/0sWdSpO+K9nWBojjL
tGILZ8/NrtS+t/T3skMuppu5U/iuI09YB4Z/rhcK43FjycAPxC76RGo8KobSx1A+9DAQxKYhZvH4
mil9+wzAdwvc6MwoRvb2koQr+0NGe5/wllzAkykePE2CgcW1jEInjz7ImsREQbnTPYGGZJV/XsvS
TqrXwQHnxYQwJWuPVd4t0wVMkkONof/O/tOCFvZeGs94tJD3BHQ7RPKjc4JCZcGQSe856CBTcRer
BJ8g+VAe+urr0tRJUPf5fiSx9GmwUZeLBpkiSMp2gPTtDk9DM14YWld7Pem3YIMrS6K2UbrLnC8N
3+yi6mCqjwH/xXWL5Fe6eoKqkkRlOyNFG/TrmZAc5hERe5tQMIBBfbn7qpAcznM0chN1El/IScgL
N5YOi2N4/7EB2xU4SG7xv2lMjXUq3zjE7gIyL6/G25Sev70qv/3AF6B4Z7h6ue35F0z/9o/zU2iX
iydTd2S0eddRRvmv33YzEORn0wO7k/8OYG28q3GNF/TYzZ6qp/RA+sfmsTVZne1bfrRy24szoAhb
W7qFfMiQbp9Qg9wBb7So+yCjbt+rsFh6qAznQyBP08PmKx32O0l1LYSfTBrwKG9tYniic+aqILQn
Bkqb3KQZrCuIHYrOFWkYXTXpBZUp8PkG1qejqsAR96GrT7ydnqkAeN712Rh5OwYUbnvXlJ2+BnVj
jI5VOAiCXvGEAwKG3QYutxC4P6DzzZjipveRejtKYoaN5VwaMjnicWcv4p1duVfXBxXGyNaln6Rb
o7UNO5w+pDyIku+WBjddoexvC+87ECagoZXcPrssUcl3zBDdhumrUzsxyiDrlqvkAnHXQStorCAa
JBu21yzXKwXoe4n7lLeX9KCYVr4S0YldTl+sTfRQwC/fm+3ajPwc6FyUajJ1aIrNotFlsZ9HVsT+
ZzJiSFVsabXNEqSFI90L8Ob/TxEXdwLsbw9recjPCpIw1qsPTjAik4UEdejobPlEHZ6zY42RGkH8
E79oK/qdiKx6yuk9NqWVwEXlEI5zHr7/WGEFCWWXnXu+cnGeFkDIqxIyR5D0FTPzgaLItzlo/bgx
+RacUkKC9s3AYI+F2KBnxH4Grdqxh/SMqOxYSdcgN49LiwGh1D9GoLRN6go+u0Jr4Rlq3lIQ/7cH
seRWpr+ZDHPAO6kUoa0FRWePTCnwXCkmJjarsDGnzcXZ9kje87FJheODz64AD5xCWSXYJNKKFjNV
lI+rIindNy90H5Zd7LMy8/Gx7JqxpGWTpuLiEKpE4b/IOomo3DZ1LCVelkOCdB8wUagwzb0IrL9/
2XSJbkMHn/wYKWAa6X6xRm21bjYc8SUuiYyGDkOBwxyEJ0ql3L52XevQQZAAlFNnlqo2K8tEn2iT
lb3t4CSQVkw0b2e92tjHXGXSwO96PUl/PaVSCIwq9gtLGTRO4Galum2q4ERngNXh/g8x52u1vgGz
73fQfWIsEFPc3lwb42gl48Z/j3qQxcObXcsH8j+n2u6ZbD8Z510foIl8qAFHvX1MQIdHgYIJFJKD
ABPfQFLIE+gwI/bUQXy13NCL6D4YLIou7vmYpuVJtkJkYhB4CUn86T5a8+PIcuRvBPkpsGQBcr5f
saaWtlAl8HTT7e9TYtuVLNBv8f4T3PtpRbs5A3znm1qbxXEOVUtJsRE1UkgMz8rg/KBmf6HUpU/9
RyouBRdLHNd1kXNb7EI2fhq5Wofy4poC9/qk8miZXRG/J7A7cefbmyC/gP9vKm1P9UbuTxVLveo7
akREpeQPMfLk22EVLbxdKhQJK9tiMXXhrxGjNizrXmxi+BCBWlIMLalmiMF9V6g51kxPeCK2X/MV
YUybsHIPqNEoZ2J1trFp2EXkQvNPea53vpnbTmD1eVFcG3FSN605Hc6i6RDgzfieN06j5wcUaaCv
m9k3kHtgyaxPAnLccC4Ud1dedWSvaWGVWVv16XOG8w0eHZvM8S+5ifkI1Wri8okGFarkTQQjoPRt
ZYcjuKUINCCnCU/pHYc6fFXTSxnAkUfisTwa34XVSrL2Mq2wu7u8DcyKScPV6gJCgcaP6bdr17x4
BG3j1U0oJu/adI2YZ68rz05xyKHuDddk9zQfMpvaH0bmxm7MOoJ8ubzHVe7JAPzAdgvi/mtfzyBE
lv0YrsGs3XeGHsGB4PqEuuwvtdNrAeEU2nqm9a+dXQ1e1pniqOGM7ItTmTLycE7/CQH19CJmbcTP
kUIa8x7Fw8CyG4qbDzHfJE/HPrNE+UmwwKfZqepuMcSx4VLOB7c/dM5srHo0hGPgxaFbWoOgX+6C
Vi+/CvyHEq+SeffM0k9Oy/e+UQyO/xQ6Rl0B+3NLxqw6rfRU0x09X00ydsrJHvmA90326TRvoqqp
MUevaEhwhHo3HVB+76MEGU1wfRO5dmVQWVAImuk+evnrFYEqiSIxnpTMci8LR53YegC+irwALm7M
Fbn1ShnfbaChlV8oepyD3ocbO26MKHo0ag2BGNN5UAddCZ20GGaQhGGGjEw7S/vNBO4Y/oWDT8Qq
ncSLmjUMrIc5P5ittxCW9vfPNA9eiKBqCLTdnmMwjs5bU98WtPoFf2aSxTkdjiXNp+ISwudnmTZR
WoE0v33GrQJBn5sZfbsVes+rBnoHPG6GIxntdBnMcytU8zHRkIMPxuxUu3bun6CvnhoYnNwG469H
Ap/Yw7Y9/A5FIdzw+MaeluXHZWkTgjnvu6AE55C9h5y34vLyQfnRzDBJ60RECnVQsxUw3IUOLslN
vhDtcwNcd7do8DwrPI4Epg7w4Ird2rSRuEBt6Cbb39DsIF8M/n7w405AX0eMrqs9TF/7uQ8IBRUv
GgjMIyt11V86rmh/9wr7Kw1YIOupURovRJ9DlcuBPKny2RMy6h5UCiAz45X009ucPT+h1/1Hdkrq
iyY3IiFCYOEObegVOgV6/l609M6LNCF8rK+aGU2qCegVI+aiRi3+yRy9ohmSMmdjB8hcWpV4fYSK
ANmUU7eWFgY0CM0X4GZWjsJu3rnf/4nG3h1zoEdqpslQCm8Rl38KMb+PRhui3QPg1BWxO7CqEBm+
R/IcqR253bWOD131MT5UHKJU4tjB1278CI6DLnIFX8rOu5G2W4gH1thylhXxWFe8xtmbjGW5peRw
Pv2rTUQQ9DK1w4gaLFEUKr9eEpkQNjnxsL02puXj6AezEQTNhC26uuwelxRdLC8OY++gkz663km6
/YJJWbSRISRXNhTSZm46S9L/GWyh0dUD0K0XuSOTfyhiXcc1vpw+IQS8v7kfA0jMTyAcI+ZLyNXD
0LckL0NE6P2SddXGKFZucbWlEjVhPxDertbGWJR5QulOpNT33VcFLyyv6Iwz68cErR2/AUbcW9mU
Of9083Ydn7tRosPbuXHKwGrZ2DOHfy/KyfJ8BDazYn7TI9EzAzbug+HP3QnDbjhjSq8CkLhpzkGQ
OCuXwdLuo0DP/cwLTmNimssoLV5+xl9fl+QFzG7CVE9Cch4nAAI3GOmhJbygYVB6M49jHH5LHGau
EAEIzfmtD3rDt0Ze4y6O6F1anFYUnMQ5NeGycKaKGAqzxDth1WOyWd5BfA+Xpu9dhUY7U1O+pGqx
GeiCwOxzgidgBvooQRucIaqJoR6aQHqGgpQ7f6lmOZCuwNL0zudD6doui2d9Yz9YBCJqD7oYiKOF
7D4kcIsbTTrlOvdW4E4UUTkNlXyBwxhP7kt2wrv+0PLP0tO0J5dz/F+QaSkS3JX/5nQhjjVMK7Kl
B3QglM5NHn6nlrmAo6xjSKZT8gd+5CYI6slr1dT6R+JySKU/y8aTQyI6kM170yH6Vk9Nm8HXKu8o
+MxwEtaGvFUG7spU7XpnRAkhG6xnl0CxjOJULNZ9qv95VNgizwqs/5fyfU8U0CrdK/dOZMCx/xAH
0nEy1Pma4g8mczHrzS6ndXZgTgxVNQnQ1l+ycuNmVM25l2Z9ksq0PoxAJYetQOUWnzstzR7L1kr7
Q23W7EudW9/wRbG04dbWpEV8yuP9prazTWxEMa0SsxLcMc+CxEyIFH7nosaPrRNGmZ3HjEv2vT1G
dzrqLWF0R6OPjtM4quv4c6tNVFkRFNH8Ok+EHaAHZNunIQIt35wFZdmPcwh+khAflL75OR8yw8F3
Em1K6oI2izxW4q3fiIz9Fh8rpn/ncY67GWKwP248TgrcdClwaRmXdQHH6uDicnsbNoLUjXiVt9Oa
CyS88cPbSCVmc1QjN8cxkOP2BBmV5L9i0zS4bcWoLAGWAnOQBV2rO9N+TqaxV1NVBchOW+m6Km7w
VttMSUCL7KXKMGNEqoNC9BzQNTsz80oT8CBILVXWWNlcgz6LToMEO+oM1vDh9yz+eW7GQDqLfEco
0Zot9yoB6pnYScw5C8BWW4e7MMJ/6swGBKlSns1zidSRQmteGMctDhARNpny3TON9BTUDu6JjXLx
/6mnqcU5787PHTsutMbUSFwlX8f8fkKW+AoUOA94CSu6KBv8CeBBT+l5OCcmq8RPRlPUB8eHJCFf
H+bCljKHUd6fG2F12PJjIwPD3bhnhbIIUh/kW2CXQ2aBglg2Un1zqmUn/00btVV7naENVg9Tpg17
mSaxLea10c357Yymwf8lhkEJTGOkZG0yuhQCrCZNrxF226MnwLk2rRocfeyC4QmQoMaVLXnwPK5s
LLBRWKTu/nkWBKcGTTPT9d2BNxmNCjAOO5QzFkWQHErZwnkExI+f6g2E03hTz+xmqwNfuTdtSFgy
DYsn1fM3b97ygVIUGrKOrNER6zRrxyH/SrEGyBlgyjejKiHTJII+u7vg+00SMMp8sE0pIJ7WR9yU
5FsM4V0nmH53BWqR0gCAzPuq84Ezc4v2R7JaPL2eTeMjP/C2M6NYKSGVoVvhYyWe19jS2Hsq9wV/
jYZp61cufrF0ASrJwGnIWm4aXmucTDW8cSNnRQPKP24SjsyZz1Ga/hqcWH0szjbRmG+FU9LPIpie
VskuMXR0ScbIWRJspYKLx79yBgSCHCtcxATWY+NBmBOs5X26HbTkx7BpmapP9aHbu5/ffxY0QQn1
Fk+lYSsJZXbu/7evrDH0gLSXiAu1JJKGc6hMFihyVg+ZGVMhvFydCtOnYXbI7Qq/A7AAMqKXXq5z
fsOnPg9VxSa8QMpDdU/cMId3zjsjMf0iRDS9ajH2HmN4Q8MQ9oq72y469MsCZAayr//jpvYdIHdf
e2VuRiu+LguZTPxBrFV9pNoS/8avIggwKUIgNxDWofzZA0t37moKtdnJ2zI1SAJnXERFH6EwGEXb
fpGwoT4oZgEEmdmZv4/3K7AZe7JYb8PXXcRbPzjMvM5OCpNSiC1dfbzjaoMviXy5ti5wri1Br7mK
5DE+vsWR0cZitOV87TtIFgb2Ycyfbims5JCeIhMyqxXKFM2b93tPqRc6ooX/Zbq0XcjT5z9HmSQq
VOcqw3p5TBWNKZ1CC0km2f85RuNg1RW2qQxqrcz7O618nc51CKbBZMQFybaqMzirKDBsXCspqhRt
NU1lb3FeDGjyBaPCtxBZXj5y+pQFjktJOgufxymXsnmwzdlBkG6nNcfHWfFCnLJ2W9cBjGokeDhW
8wYg+rVdENKi71FhK9RuFnECpAyDIh7Oy+EVBtLAtJkS010kv2Kk3Nu7vaBcEJLA05ok3lzA3Zva
aX6xJ0ER3SKYtRPGks6aScIgfg1x6+FrPNi40EpuUdpUliPGTysG0B3TNN9czNl6wBqT9Vzm4sUH
EsEcWzwKKaCaR7BFNWJmK8y8ex/CdeoV5vw+pH+5mPqV9l2+ZkC4Ca5OZWr7pxUKFIV5Zhj9PicM
51K/ErxgGyOon4gPZzKf8BWUyot+qpmcPq4CpwpKM6sBoJRoF+yueBPJH4YEJmfel3EGx02JhSz2
Z0H5OrdnQCb/wKMU4M8KyySwbD2lIe1vOLOko5Fyc3vfMdOyvti8ofh1T063FIWXjdodX4I/Ygng
caanBUiTg6oOS8eO4yMpMROyp6L5yxwxrvxqEIdFiOIMPMbuMech8HE+YUFl2VmP01YGere96eNo
h3dVSxB33rjIaXifjP1rSdAmKR5/AN4RIA/X7xGqNLt4R/5Lp42e6f6VJu0bCgZukpNtRiZ0dFdM
P85Z4R+8VmlRw2edSve4jOspfwf2FIb1OdMhF41DyHbGs8tOrDN7dP1lVeYXOyl923eHJIC/52sg
NPZf4Cfs3ZILZkqt2cfDk69YNRmxQH94ElOCGxD9dWwkOrmuRud0vOjBaIQldqNs4Y/bQZvsyG4c
qM/b6bRtKWEMcaqkIY37sRjTdUwRmS2U97xXGGsksKMYWqfhC4u8YRq55eBQMwQFmnfPGl8QvRYG
stz2w2bt97WEr/EU9tfeJ4dOkOZ6XGbEPyyAOGd8g6OUaKQkJPsjGdaLqXUrpmshZfdiE7GzqEHl
KzEZKjAlPYUvhed3G5Q+ApSOketjPNapjhcXD3GWYtnRuKDZZdaarVHott6CO19omzz5sNhfEPth
qDW8S75WtA6VgmlKe/E1ewdAt0bgTEuE8k8JkaTg1QsWtTwOg2C7Setav3k6NVrCKTNArpkB2kro
iD42WMRp/jUeKZaD1Zv8lfNe7hXj1wP/jRyTyTjC3Z28l44YUwuGgOd1hlTey6c+AFU7miloVGyZ
TnmiCJfJUF+FFA1u+/ml4idQ3n9ycDLAjpiREuAD4PKq/cEwmbJXq+7NIl9vTm6i/9Xy8lm7V60B
kxpNClUNNdRS4rwgYTjwjbA3JMwg0FumyzhExln4AofS18DAaeYDTWeUqAAr7VP8zSZXOnxrU9aO
rMencY4XIWuc6cOSOR03FtDC7AP93FC+iW9tPlYaJ7fLOO5oscoEA3ltyU1fQuea6196eRA8bClV
+x38TZWIYswPBRGECJsc8NZijIbCOGmR0TOU/Ejmtgg/FVyBAXLdsxAa04dwT3vnApfcIr3Fg12+
io6eiOSzLHiYDzzTMsZpZsoA2jaa02IVMgzmH6YTRSAgBb4qImyTa1K9S5k5Td5NCAaozfRndwOH
Vsa7+1nAOffwzl9ncsdN8WR0lyxPNBjQF5FuoCazW83J/XkHFoo1mQ22/XYlL+xSTr+DdxmRUUvA
pqYfUrB4aEYskiAxP53Kod91WJzVK1LnA8Wv2H6yx9sjdzxYTt/BPCvsi1u0dtXzVTyLn0Ze+72b
5s6Q+fwoZCXyaD2k2qDoqgPqn6p0V5+tLKqvHRK5jc5T4OwKcZr1WuMAqY41NXj5P0owvuk7FSj/
kV5MoDetEsdI6dTcrRwtDzr7ALEOTsucWK7QUggTioXSBM6/ZzX7M8Xo4Gpv1IsAHZEh3Dm676Ty
Ij6fT3SiQN+taz3gGb9TGJuRn1pTQMNGi5X2/q+olcAZmSxaUFB11Dd6/VJNMAuL5FtPNzS0L2KO
UFBTHG1qr05PQJmre/CWih6SIKICI0YJp+Nn41H8LuDZk3aSVC2YVlt/wtiscYrhSN3ke/yau2os
dSXRmAM6Tz64ykRIRAqDHzH3/uEw8enBTqAstpQJctu6hFs6ZmsGlcYlSq/PBnt6/11fbPY70sRy
tyDryD4T6djhHQPgP9c7foCRp4Amar2oJ4xk/bQIXYKJJwqPP3Uy3zdTcz/++rC0eeNgOV8CPrNd
mX0ZIA2KTGLnQ7w85hk9ahJWfjR0mhY/KPJUjZ8iAFH/9WZcR1q+0Jq8+MbjYYyeaVJ/JsNFivq9
RM639sT1UL6YEcQN0HCmg6qpgmOFzB/XC615CAPlWj26IPCwu+LUSywvtge3DPtSEyL/4IbmJiLV
1fh4lhxH7TQKBwXxQH2T7d1K1vWyAci/wo8lhtOGC8h9MtWjtPENjgrl5d/GC7chlH7HH2gFtW6i
FGQlV3nVAKzNKJbZUK9mmlGCbOP3opUq5NKtH/u+HvEHz5V9hB/m/ehwH9IG+q8d8lgaUfVufeCd
vmdLgL6FDh0aajb0Z9xlF31C8NDKyGQBzpI4PwgBHPbgNACDK3nBwlwSnO22jGTUoncE2sksM6uW
i7KnJ6BfmRscKLmSkh+/uoNn1hXGgUULwIUkSGJybGNDPF/6YQhHaY2JBxI+yz0qq/MUpyZomkgT
vzlaFDmQ6thWAyxrMjxd8qaxCqN3pbdJTMwXCFUz8gdgWF4e4xjXSFWN3u9xLvOxAOsUM+3rP7Fo
5Sr5lLqde7E0RVj2t1sfA9snru/pp/iHo4q5/xlzSIOfs2HOex0UPqJ7GuKqj6tTztt0tT9GwudM
21QYDS6jV69R6XOJ8DGp/YVAp0JL4P6H9wdu1x+8CEztZrAJenhy5WbqO1YhmpqzMVLIFjdEE+hs
cWXgWnmVBj6DDT3kxYbKFmNKAwKRwJtxukBQbm5DAL3XDVIeRGzE55ipkq13LMqC6H8gSB7gm6x+
W2cyI4UHMJqGN0XC3HWsgqiGqkULFou1Qqamr1HagUIIUAT4HANk0jiqmiyiQD7Xa2gOKnb4ZPPI
/BAffLkiNuyOt3YGWdemLWk5r2uI1PjQuyHjo6KPKfg3eD/5+nKWRbB3H/k31f9CWZRv4uYuDSW6
M6/v6oonQpTKsdMF80sqWCCxpCzc20hFO4tAFRm5gD+vx9asi76rTbori3e6laVDQ3/SzhJouLhr
jqf7vO6DRjNQ+8/i0yHINRtdG2oh+9wEBVohT+oO5sMfG/62h0/yTlHreNDTSU1zLpmpgeCpp+MK
+b/HISr4lInV4ZXD3ttQuc3pnSvaoeqz9YzAxwf1AOgjk4gRRcmAMpx1rweLDN9qekth8bUX1U1s
Kq60uN7gwxshEs8MKKmUVSbcg49Mje8BPSJcJ0g9nUMNH98Se+IwFy/4L9uW3LM98Egpuk2CTAnZ
i04Nalf1+5Dkb1ULKUBd/KXkj+NXKyuaQu88LDsM5Ch2XmHXImrpCjQuTGR7pWB3DAoqYchN6Y7y
ZWRKhUCtt3zhYYxQaXRSUm/1u+hvdluW33kJ0mje+c98y9ZJjPDqwQyJgo4kzbcYIzK6dqqn9NjH
RruICJ5zwc0NW5nKGApal85Hn9DetJeBVGDa+0259pdH0Un6CrGEHRIa5AmuB4AXgamhD+XAvXgb
4UCixQA/waiatYfmRg/205wlfh/wQaoLQ8cM2LJMuos4rLLrym95f7EU5UKnSq3T9T8W+P26bNCB
lJZtpIyLkqn4nmCvicaoxGRV94k0wrKJfjsQ/Hbb43vvcj11ADQo7ZAM2rq1alZRP1FGmgvukmZO
++hdYKtmzgPuy681M43/NpkVh47UTrYGqx1yOYhLkoIbcrSTr7Or5/qAoyP46Nzg0EgJvIYcGZ9h
qacZXIW+O4Ff/rolsZ1aqUmlI3zHyAIvgc/kAwvsK/vmljGBWdIkyv+TEL3HCFV79gMFWrz7PnYa
fXSushGfxYx08dMUJmJRA34MRgzKODqvLbE5XrlavqIS6M0/bZdDoHTCFv8fsbhSSWXU4Tfx1GaD
P2u+ntq7geaCCPS3sAXbxXQMCziUTPw2r7ZE5Vm4MIvYIpKMyQclXosYpKt54jTguEDbojwJl3k9
bvqoGcW9eUkwdkF4i+7tKYSuQdl+1ponbcpDbSW4SWo+o8AQb1aaOojZGgaN1oF0slIf6Uph6sv8
raAfjyIp7YCItR1HXODUdTcO7qEJg7wvfTs3hOVPLmAOaL7zlkxuriCjul4IW92yOVmPvVEuA40m
3dNbMvGxZV/akhHngGsJ+Qye+0KJIp+vaafxf/mwHXI8gWP/CB5k5GKTzSm9JHwPGMayXYyUiWxr
935NkpHFFyNi+JuFLx3zg/KHkk8bkK1my5KF7/0buIAfvu3Yb7JU0PmPm95CGHiiy5soQNu2JdS+
/3B2WlyzDJYD73s3p1sQKkYMwZ6j+5D6KqqaoYR08Ga8v0x+7+3/Jw9ddVf8UODxaPp8bdSMkrbq
q/L6GjwKlI6VsjZ59aTpVCBQQ1M2lVfjk/grbpctzo1UUe2nCPKyAEm7/AXO1Y7GBci54sQ1kZuT
1EV2t5ymxakwvx/N1/6BbtVwrtfE+R/6QwXgs4mMeeReYu0cnrOoGWqHJ54MV++L0Kl4F5FHV4/2
vTl14oHiqoK45XPpP1vhSbBybH0GXHwezZITweoGrAjsVcAf9zIDp7GpJ4TR2P2+A5+cIvwZr7zo
GRCDuXWM9fvqJMvsOQ9jF/m0gexob8APOrwOos2MKoVV5Zx3FVjKRezf1RA2MAVUhr4BcCf/KRA/
gLDXrplw8iz/P4Ta3OMtZKlu7fTnC8lZGCEeyRHhN3vHhu9e2fBPbfwF9JANj8Ze9iM5JgBc8reG
qFPH3JuznrJU9Tf1e4lhIIzmvrb6tn8W/iirbhN4Q6FOlw7OeXkUwiRFF5DgTxXgFUfKEHJc8xE0
1ijmOC6EJrn9PJjHfwWPtLZJHySqOYc+zoO2VXZUniIHpvCH4Yn3K/EqDDrwq3pFNRN09SiF75mS
q0ijPOhpACP3fFG/xVl9/uQEb2Byq5sbqucgyebmnz8vbbmZwq7mjuD4HXcAoixqrzq3IQkpdHWo
B90fsR3x3JFhbcE9kHhajIPYC9q5jN+U+EyNyr+qi2p/JgTcZO7D5tWTeKmPfhNsPuYTvPKcGdjp
L5Veczijr9f0Z1DDCoIAG7YgpnzXA1jHuEHcokOTXcj3alPeTCUBDkMd8ikN7clqawqMEV6/qDkf
aYsZPo8a9SGsIri+PXsh8dXZJL8pYFR2tfYb8zc4gpSJrcA8axxWrgrlLunc8bLkt54zHjwkBexR
/iuGLsPD+ARn7XpQ+hqmmVcicic4uQykH+hLWb1xtxPVFR5fEqbPzekYpaMw4YrUde8/QAJMb/SH
pCSYTTg1nNE7mZ91McdrYpvVlmuaQQ+iPlIFyh8dOThQok2cZM5E/M4K/0oIGqEAGJaRJn+MT5er
ySUR1vgpSLLwtro98fn83GWWHbtlbrRFe7m8bEGP4eB1Oz/SXnNVpZfKM0ETtiM1D8iqYhF4mPY7
cBJotCAx4gNbqUB2cNWpHn0ie4YdQsoJg+I4A+h2RU9ZXRnknMNbK9uknIqqKv9xX1DmZnxlrDc9
NajTrJrbXahEsOHJM0u7q2B7VsFQcWcf8jwpHMJt1Jw0Fo/ryEhztzykotkFfv5fNvrQjAX4XHhJ
pGN9N1t9rttDgQNC43jOds01Y/hZGNT1HNnPW8bm6KC2/D7HGk/jOkn4fNEfxI/mnW47TJCoXaui
vZMdvejNdUbR8OyEZQKmMjreFYmqhUbOtr5cxON0q1fuefCrz5si0P6lY9dXpGw9NQZftK4Wr7cN
Wqs/Eyub04mmXtF/Vvg2F0/+7V1uk6GokG6SnA9mWR4j51qwNLD5J7W/34cFJbUCLyYYo/IZGPxY
bZRjtSIDt2wUFmQSltmM+z+aSv/itP75o0KQvdRXEpofEeHG2NuWdepz5i5TT2xzyo50mHkBtVsx
wty/EKRtvMsYTmNHcWPH92UmUYh8X8BAwixPiZS/w/Ei71c/CjGmqtvt/z6sfBID9U3ZzkIL/Sab
5mQjlmNkGikGeIDUsssqOFfrVQ563w+4zOf0GYtuRAhHi2nL6MFi6GG9hjRIdVdGw4WW0X80svt6
nGOwa8I5A89Awok3RGCFgFLd9GreIrG8qnlcHl+5VHR5ToyM4SqpxU0rhRgu0xAQja2iKDB8NiWk
+Lq42cddIUevhsMimzyOf/MqH63BXFzGt+K7HJpIO9grNgJSrz7ZSnqkSbJ75/7aoLWVajhbSrWc
yZoR8gwkLgtiVrG+NRD5ayvNd/oOY0+hREm/JgKJrUqq4M4ZJJTUKf+9ZGEnAELnepi60ECMBR81
SeTfiNgF5Uv6Xk10JvVlfXFcjy8doLgQETNp4GRiz5BOQkjKoQIP9IqYiz0qgfTCX1y66cKVWWTo
KbvphfmU1suyBONXhNJpILWEYixfrVzPKGGZxwB6pPJcJKX+gOrloJgmdT4gP6VTYBFXal1zGGN4
Zqpgc8FT0hXdK7qVtTgCZPkUxc6hE20vxflUFFKWTOFYDwgziR/3js50CcTSP/f9Waef/Ryhmgii
fUoI/Y8SdDj94qqR7puGj1of0ELt10TMOUz5fERKb6PnzcP4Jg11t0BQh2horYvtaSSYGd3Yqo8u
LTG0s+UWjL+4Ojf2/X+v8bCNlOLaS5gWmwcFlvAzMsX0KZMrwX9Q8PPETvqiiheRWcYPME13/lYh
oXHMb5dQ7ud6XXmo9bbDXIVC5zkhfoudxqKtOZQ0ejT99NahNi7sNekqBB0aIHTr7YqGSYUwMPkP
OxiXBaPEw14FQaMBYRDjILqiCLYZ3xwEGHIKafHAzkoNYk4essUKTfZdVdkEFeSX87v0njADHfQX
sbqHkwMUQjsotCR52mNnxaTOLf9Yg4JlxY7xhYvofB6l/n6Q5QtxKyYKBlRVhBleTNH8RZ+uwy2z
hXu+lHoSZf3oxbL81XOddF1Z6KftxFLwz+V6tgL2aBfzlHoPKN/3fpXfadWhqXZhiq7BjoiJ/8v7
H8VKNPXBjTej4q1DgB2TryBNGAdxxQGLPUka6RTjgR+cx8eJx4HknwWfDNLydn7WYL3AD9hzrikl
zomrgexBL4mXo3edVaBXcloO8rtaQzTSrxgnM6Knl+stg5i+Ith4HBIAC41nWfLX9L9ErX3Js04P
kHTMWVlX498TQEbQ4zOTow1bBtQjFMjs3brmwR+EG9ZPNM6xLE0L3wsaKKCTCPQMwL8AOBxDqOqw
DCv9NJovQ9G7R5gsKriMYfHSw821to9UKiPhTrHO7TQPG/PQyhjEDDBRfM6yIokkGDd8akMrwNo/
fxJUZfTA3IydC4294FJOx4vdfse9Hk9zRlC++t31dC02b1X0KuWMbFgxNHRD3BM6GMaT6eWIg1mo
HzbDkw6yiTh1Mip1LZOzbRH3n9RFZdcXSQNXsQyJGOHSfahVb275fSnID9JGqORb7guq/rSPUjEF
fkl1HRrVqzt3V2qOvaVCY/K8poOVpKxxxQ/t/E0WiyuW5q7yB4wxboowN+i9IWpR26BqcWnhF2oz
q9NMIZRfszgdJ10xgP1Ig9XhYVDEKrIyuiaZdkG5cm4BbNucr29Xz/Iu2J11T7sTIAXgN31zTEoc
sUAS7VVzmpi4bvypNTHG7GibhXCg5ieNpehHfxLZ6+Xc0sD+pCcvoioML7uM5a/G9oICsCPU43Vg
HNHfCzSNLUY87wl9p0osRuYzcdPFKpmkQ0FZfZjdvmiITKVKg0m3QUNHjdZyab0h8XnDhLxIYu0d
82ZeJx3YKAwO+SvgQ4L4pIJHJ260RqvCV5Ut5/Lsegdalx4xTKsWZKjTGKJnLohKTCE2aXN7HjCb
QdYPrEPqfV+GBQb45Zh48V+mkJJLRbiDy8OjntTudlljm4V5c2dsiLCuZmu3haKXmp7PAwjvuuEE
fs9FLrpZNRf3uFYfuNV7cJkkrV8rXyHWIMi1lIYfr1ZefWehoULhrXko6MBFbfx8hIUtiEc2lxWn
DY3w1fmN0vSnTq3DYCaW9+xny8H2z6/fpJ5j3MJMTY6diZ3aaGRTUve9M4JU5qF+/zU+Gue559nW
mev3dTRQuqOPyiWGERCdzxY1EMrK+7V+QK08OzQV6VUwxhbTqKN6y57q1MSqfpcQX9jSU/przb0S
esFcVlOuxX+ZaIHA6NziMOrfgWB3T6nu6pINtkVRjs//Jby9ECKuIztcRIqV78be7edA+p+MiT2B
qjmwr0mY4Jo40nCVgpNk3FB2whXB4y+zITCou9IUQGu/7+qUNC5VJGrod+bh8vwCzo5lvw0Z3kBt
xeXVZJ0c9jMVZEdhaOYFW47inZtKEDOSyse+3Rj0Lx23lYweJD8WCkfGb1bBcoNDmE6JxM6B6HG5
jXMLKuA5wwgH7RWACMRGNAGpnCLMMP58lB8c8tNfbfKDuiBaoxW4BOhFU7BDEewRUDssdtgKVZVE
dL/qNZQYfVb5EwXHNeKwhyGpot6DYFR2GdswponowQEyOKONpNvy2Sh3ObW5eoA3gUW9sZ7svRy0
1h5AA44Yx/xSq/rNDP5XovMwzdfzC2uuUmgWLcy7nLcmEXIuZtKRLY0bp/OEItFpCTmDAhlgUnSb
DJFRjGxQcQEe/ikdyUaQhEGlVcF5dyW9ptRzj2cAQY/80hWMkIPRGN96FDvzpxqWnhwmIFuBhGX2
3pIjT4cGSF2DXvf8e3Bb49ldjUjAms6jKjTAfFndh5POOGigvkx5hm1Nlmvy68Ig8H/Or7Dbvzpj
q995lU+tvnAflp0DIcHxKG4hMEDMit0Cjhc7nLYVHnoWxCqNl0XAHQKsCjSkFhm1XlsHkTA4S/qs
dQHvCbiRezforNweT1FbPAWeWYw73Sb4nETFf1G5dmX4vBFHEYgy97SRVVfC0CVpxzItJmvn4jvW
ohaafO8ePvyfsS9GhAz6fPohHJgTRaJqGZvqKxTa+JHvvcYT7s0+fFqBgyNyrvrG/yL9c5STRrh0
j6wvaIJ4+0tkfU6UYSArWJDCRubl/O9721BcO6dl3hwj8rzZ9hkeE4xUaYizWVKiJ4+N27Ix+Ag3
2uSAi91XhJKKwrAN3nnrQ/VyU5V7Wviyt7pzXBP1442y6W4RYo3O6wHh+0/x1UgiYC/mTIQnY3zh
WrV7sMi3DrpomaH51EbaMykGbQPnNB2KL0zL6wr7oA9m4FN963EEcdD02afuNvnYbb7MPIYVLRlb
MgK8olNQO9SFlBzHQt5elBLoSGrY/pB/frUxkj7WVICY327HXbVqE3ThadTup94Ip+v+UVzmOxTQ
/H83C8RJCkiODahgS+UzuVkD4SldODdNCPMsIJ0YFUjSWpPQl1TvTFuLtrNYrzXaOryjC5kGFokO
7TMSk0ugkVbiGpMlmxvhtjXYqvLXmH/NUCVgmIGZcTod+sCO7yyMZNrJs2OUrP3SMHP/JsFT5ekh
DTxfYHFCyd6XTzyzEt3XLV/BE+hvcN/6Dt94Xj7M0ZfTo3Voa3NrSM+9pEFzH6bMQzRMKRb8aCPU
jWrm/U/zmxNWpylDDT00+5DRnE9yZfpwigp1a+O6QI9+8cR9PqqpDeU3ZRp8IV6lKSvT6OpnBhsG
/PSCstUyjKv+DisB3FbWFQkwy2k7j9wWYzrD9KnmRF1BGJ4lwNQinoVVjAgQ4O87DiytC5k9txFj
OiwT8Tnc4DFXDiAz8tkb4Di/cUEbAxT2rZ+GR+6bK7WTO5j4p/wpqT6Y7oASFmr0bMpb/C5xuPLV
8olshL2FL1NiZRoso+IUpt365dMLGWjSNR9k9DHp46dQowRgDdWWJ7HIc8oO79fmvivXlh/Y/1ZZ
UFIcGye+2phDsz4vqRKk/ZiVQ/fLvCWAk6MjGBmpYJx3JqQZLc18ekJQUd7YS+rjI3lAMPdUa9Gz
8wJpN2Dccoli9A7AbQLruB2hqZKqJN1yyjzXdhuNjVdR9bqhg5EcVUeCqninx2kYY/3meEwkkgVr
g9VsnwqK8lD/7tUHnLmGQu023oJP09tptMaDtjsENd6W27iu9N+KMcWKVw/p/lJsPmLG8WiivN6O
KZQqc2lyeInG5hsbk4tBAVfQVrwoH+nC4wnKl70a6dPp3Zu/ZFEUhoVF7WR8RLQc6U0rgg1S3Xsu
vn+kfW2yQPOtwDQyvdHUnEpQtW3Te0liXLfhHxp9OMbpyjaDGNvL9qv3NWM7I3vUZgfGj2V29ZJP
XVQT6l7BBJsLBCsj0884tgb7MPxJTQ22yk2Uc2vbhHAb9i53wMqk4vbqzeiHv32QR18AoJwM0ZrS
XrQQ/pcx5753MH79XgmoRhWHZQ8G//P8jak6mH9wbvrx6g6YtXV3nP8nVBXL760oyiUOBOdR+gHK
7A63QPACH9R9kwDlMAmuBUhDr+wwgI1gaJDIO/P7fsCNp4CjdtCTRiqvEUoVUeCwXHYtivl7AA1y
5xPuVdhLBgIJfbjfDA6LgMsmRpbogVzaF9emJCVqSshSqp9KYulkTNdBiZnNm+nJcXnJoS9rlywA
LdjGVll+FnIeMj0NpApza6zB22sPuJEOIT/wldPrZfdnNPqXrXdis15G+JlICg9QTyMt/uqIx+IL
v2TDq4KbASZDywgO9pPcTGmcG+CPBRZfPg3KgwU1r4ph89M/zU3nuV/4qIf24Xw1s5V1fCLj8E/F
SvCOLp3tlmj0lOaE7SiAKEkE5Ln1WXzzLkz+OWWVbJ9iJZVolhpk5ea6Fu8EA3JKEa5oa0hjwzEI
7a6Mnu89dPXk3ONk1+UrnztP/vrjvKFvvViv5rEmpZoL62cl+UjIC8XVHKL54hYM+RmxIUbgH/LA
Y5H9nVeUJ6nud/mgJiLFJI5yG89P+R8vq0rojtdhxM3BE7SVyK0jX3Y2gly3bg/kOOitQDAgZMEB
xuLTnXZ/+z8gFWcXluC1lNabN3qGGoDq/c2HtMjmNRqv4/Nq7HkDtK+k/FCB6HF8KNLrJfdJfgLh
o22049YWN+r2zKC5vDyk5wJDcvGgmowyYerkbxLGhdWiDJYJBIFxDUhnPZAvd97fFtDJV5UvQsno
3YE0h4+oCMJWbybHIJwzNk0uuteGelMaX23tzCHkXHC+1bc4uH1NzB8VJNDjQuRhRyx0pxVGEonZ
opsSV4r5FmeqqrVG1UMp7encYkDfU4AO8Xk2j+SSEj4SiRErdEd7ymXgV14jHCZ5ogTx1IpIJHgT
S/DJh0qxDnI6LDuRZDLKtX5NbYBDwPOlKv2gRBBKmS97yerRypLt0MDtjQl66X9djJdJiNBbXqyd
vBejD65KPxrV8sVPIIKga0CDMydW77BsiFMwW3ARaM5/z92PhDqpwyDgfNH6qkZGiffy2xPn5lnL
LCuR0b0wOg9kBPzK5i6aP7Neb+VMg8lS5iXxCzsFmU8M2yAi9Z+LxLLciSXwZ26io85TvL74t0or
YG9QDB7ZwTJt9fc7HJlSsBgCBgIjmMzSPPzS7btRoCx1jp7Mye7z8wlNQ2PfMP3a02D6jWjdIvY7
1ZkEv4Ua68T/VB+GQCxIacLJJSM8o5zOdFsdkX4PpSuFglCEBjJyNQWGuFmOjvGuWpT5cua6LEgu
nHyW+/DrZ9r1ybglHnb3cy0S3f3FutV06dc2Ipls7pDtVIJqpAj5/ydusduWTRyzMWNNhaswIq9P
X6ysAc4uTzk30jAZi1X/IeIuqJtgsue/38CRmZWMAVKwMjKvolPjvOjceMBKkWOUK85OrxePG8iB
MYJkqgHpE5WT/kNNLcgSo1AnKV/Atlce7xT8XV7f1F2KdxFZWyMRUC94aereRXVN5ejieywG+Rel
1KTIaT0W0VcZSqsK83G6UDb7kyAbs/b1ESq3DAZ8x5WMtISyHoUzE6R/3abeOGlie8uAct6Xdvg5
foDI2cb/qES5xgncdDqm8fyLu8UdO7tofIHoQpBOik2HqXkwe510dEfv21hAGLidVbledeFiFmSa
zIlekangaz+eVoE1vufNvvPKReun5E0z/QQVojFcrr+yw3okUbxCiwaXhKYs6vVX4TDMFm9qTR7s
r9oK5UtOJVtzKA2SRQlEQ8bdW39SJRGlzDTId8ah5Lrd3UcuBD9xFE4D9IF3vO32ZJyAW2pVJsq0
zKrVxVZ1zZ650uvBRC3wZmSqCED9bRGeJ1M9DaZ04QJV0qcH3kIP8np4RKU/BfchZcYS8wxgdITL
BTMDiAnT8utG5M20XCGD+sUE7qP39hL5j2k6mZ+4CuUblWJ9pzyio6pa12MXnv1cw+od9b1GNJ7k
VEMqTYGJn2w18YpbO+4FQ2ygiJ7U3B4dm6gqNVRRirvptPlXClPChP3Dz0GJUbeF5VBGg/lkRYcX
Tn7YCqqw1bwXBOo1fQNLDngrSZ10lM1P0UH/A+K1jWjBPtHf5+PX+w4K8otP+G4KUcSCMq9StrEK
GVN2lAbnF9Rx+ulAU6uavy3L3GotqefQN5DyohzHAVGuzGKmTfVqwBg2JG+ZUak0nId6cymL7vBG
v5MYkGDdaokrDLzNqmoUNR3UyAc38OTUJmQkwsCS5N1Bq+OlUQIBa00t/3u/f+6ugu+Sv9HJf9iq
fH/1bkjmMJl9XBF1rREO03oQcBCGdTapNlU8ufVqcFY6gvP9BL+yBQNB2ws8rDRkA5N5tbk/OoEn
VpWj/JGD+sgBsiBNHs8zwgr+eo5JKO/xGOplXawo0dK2NNN9X9vZ+IEzt8fkjV2T4Ibq0fAV4hcd
hlnp82euLXrXiH+Px87XKn8nYEXXeUptubpaxCvx2sRF/DMEcVjEbBNvbAoip42hyflE9YlTcJUk
VGmyNb5WKmGRvvzHfRNERzgSUEk334+Kjxj93nokAgvcgkcjTWfe+CrOURv8+C1718LfXq2Gwf71
3eGyaD01g2Pey6SAq/vIH8/96UHTlnaed191PQ2z8ZNADIcDy14eZgvIW5enZ1Rf6XSHLIlHL4Of
mryu2J8TQI6z/AvmjldxXeYvwPyIQVhfSkxoOKo+mqfzJ12pwO3eJRflZ+tEX7Vn4vHZDgax7JPk
uyLXde+OnmXeWC7Kfiv20RXTKjJAEozxBJhtbSABFA1tBEZsEKqQCEOJc+dyCMS6+scTAgoWx3Pk
fwpgvF71H/KDlrym3g+/k/DKMqGl6A9dUAtC6tbYsrxMMIuR3bK0wFxo8Wmj7raOSO2Ig70dW/Qg
SkBqevM6ue8BY/OqlrR3PvRSNK0dPYL9dJ2QLSXHxl7niOjobxLxBmzBZLiZ0CF1jVQTsObH8Igq
DguQO0O1+vm0GC9fSDqGGDyLNIQYBAJCtcFLL9zkHwUxclFOQmF5VAokumlIZcjjz+SpYodXL9mw
mPiwcifgen6/ejCiKoIPZjiUU7h5Sla9q2TZRV/qbc2iG3D20h0arK99KiX2N7nSI3jdtwyxkMWS
kiWHtUmT84oHs9eZVl0i7n8zs1A9Eim04yPHGgpZ9ZuIGzhDJVVUnXi3ztSBqKS0Q2Av5aOCDZbY
MJX4NrXG6aLlSJUBEW8Pi7tUA08yTSr3Zha9qGVpjFFdzdEbpLOf3VWeiIOn9zQSS4XMyf2jze36
1TeUPMfmH/bOAeOCWCzSgHsIhQ1Vn/81xBPPf6UJUizaacSufUmBNcepTu/dcG++pIZ2WjbQYmCP
goxdHYDNEuJArQN9LD36u1AOgjPAmI0Er5gsIt6jf3Uu8I00S7vFlr1FBjsNpRxAED0h0ZJL+d6/
TX8ymupkwznYuqEny6nnlUi0Ts+L8Aptaa+MVxdc57webUA3OGijLKValV4c39GGRwIntW8SnWqk
Sgm12yGLBWh96+IgH/PG0y4TXmoaZR6q3PhSLGM6GFQRpJ2N01NpVhpjQts5mRiu7r5/jBJL1AD1
i+jROBFKhQ9LiSPPuDKLOQCBDcbIgprCX/NAAZSaGGIQLbgg+CVV4jHTxaEyhCmNhhI6ZMd6TtUa
pUPIJF9fR677Ngvqrh04TJAaH1vMsVqTqtfe7qeZs2v49ICZK2Uh+OGsQcOpRq7cj368eltepSwi
DuaIxypUjCmZ9jGovDrYnw7A6ja0z/HGmXvgT9QIBqv6t6na61bPsVvukblSQ32ZQAKc6GnfC/gV
Q+zZWnZxRfwMJgaPiY7/4MoJeKXvatn0ev3jOUrDfy4WmVVvlSj+eO9QYDC6ETVR40rNtgtz61i/
iPh0g4GLFV8JRZ/+CoY2EGwOwZp4/OGipe0K2gpgWoA0njjbhlUuqfOQwyHZy39T9lpZ9CksYBhv
qhKEnGJnsMh/MYHnLCqBv8tfMjAh8UeoJSw9BdH+9rAR4sm0OM7jIb5Kgx79qTiBBBsDCBFzT1hZ
/NBM0G15zlXt1g5wjC1CTUqyR6Ijgd2lFJCY07fHJJIbqBEwZ3Zw4lwO9U6J9NxsixJEN55nLhuS
1AH3GLGAlWdFk5za9mEW0xVkTLUZxaO4vXA3yW5rXdF9XuyOuJgtaH8WXFVx2tGXiKZmufu4zUkA
1e2Yh4uXFU/KUcpKnA35ovVRwVtGqbuHEHJV1rQj3j9EdABPHuWktVHrWAOrANXaF3ENYtU2fMeV
Q3FUY58HrjiRdUEMhwOvzfN0PtWH22Bx2rFwLbucP5IqWkyW3jLPbv3TUiE/ifXZDdt9mas7dGin
+D8V1HU2HFVopWvboxgd0+0WJhkbJCzY3bIaX5BCYpwSro/5rpnANh3dvKI3/1f1qLZTsVYkaZaI
LwpSjVbRPZCa9a6/z4yYH0O2E2/GZoMkZAymrXumZxjerK5VvdRduzIcxnuNfXBAGnN67Y/AASUL
nmSdOgUIZE6XLOCo4YnKhHDzUlYm2M/fevOziuXwgIil6EotpxvLLUlHo4jKIJY16NCcOlBJZFpf
E1fsvLlM8tLlYRCqzxxcs1Tzt1ftS5TfgJwYFt6YUlmG+TD6nVGQ4OBRCCxi+uqm58S7wKpKkYv/
vADLhT6tNpVfu/atsbQedfIuE+U+7pw0ssVFv3nUEW3ZY7GCJHS+WvuJGnWbnrJhYV+ECmuPbebj
8EkwiXCof/D5Yxs3nMoNNNE57jgueokQqJhowkPzDxz72G8ZJGIyfJftngC43JVw/0x2t7aXpU8W
Y7yLQ/Q6Awh/NvDL4otKYV6hme4eBHYEWTPl8sfOeDU76Gff/pEc2HgCgb80vkj6r3EFGKGGc2jR
E8KhlgkNu9UNwKSTKa4fl9mV2I87mbADgadklMRWrTwNdRtTE141H/QWaOlU+57RKy+BH3xLbLNI
n/q0Bzox1We9mdGYdjReE3LYGuuErwnCbTeWEE8X+Xob9PIOcUZS24s5ssW3VTOzLzlyP3k2oQWT
XIzvEH/+GxU9/mRQJDhs2ZgN4lHl36bVWTmBTDQqHTnjFdbaB9thSl/j4+tVH+59XQfflj3lnBe3
Bq3Am6D7THwuzEupMWNjVZKtQTZDEQNMaXx3ARPyzpJf/QbPkzLh/7rLDYBm+60lCgzJbarA1iJr
PRpJHiKjR6Npsl8kbwauG0x8M4ZwAiesxJUN2VjnzQCAwBgWl+JNzB00R+02TGwjE1kNuHFfyk+/
lh8Gu6vs4qitNfRfGG5t4emKzk8k3Lfk0aphY+/2925tdYISa3X0uVGySa0t32uZ9UeT836DwKRQ
r3AeYFXvrfgdS92dsEFLqGtQYNE/zYDjXJoDtFjpZ1CpZKR+zWg5CP2Ekacf1mLKQ+HufDFP92dV
d3AFl8ranTQxnDKcFqW5O91dN+LXLAJfO+x3rP/DH4saqT9NDF5QF9t21YgNbJs6hYd7eWNmC/8Z
mxsqkRWM+QRrAWqrmQkG0SwQP5arLT/51JITJYEwXTIVpoLP3fKr8GO+UdXWQC0JV2cqwAIxCBej
2onUSWCbUjA+ExsTnPnzvJtauhV0HAFKmuF2xTil7AYoqTbNJ1j/+BAsAiA1dPgm6VbqY/BV27xF
iOjFvrAScm3nfAUg8vuAXlPOZ94sxioq9ptfpGiVOyo13m9UzPs9vG/Gs3yQjhaNuQtDJ/m/fH5a
Jp6bsRYICMwkeosjH6vM4y7KpJCjOieD91p0nHv7U9tpgJV+N2sVW71GD3UUZKm5U8G1daT3MRS3
R97jyGqlIJEMyrPbr8nt9Zmvl6xMepPGPQExycbNVMSd6hMFn1J0p6Ccx3jp3MDC97HLGMCWidI6
5me8+H+5Lz42e2uwTpPT0+wD1FEnttyXCby8eMEZ908M2lGwBQ2mimgM3c4zAZqq/h4mg1s4kSNC
S1XT5GXx0JlZM4633xJRHBhW+9iikK7rfftuBTmcwOiYa4tTgc8l7M7mclMRnappR0jSoj2GFCTr
Ab/yjDvewrwr34XPFq34gRDuivm/GWB1kpTfcZriabZzSyVR0pf5BisAQlJyX0cfncMNaMPOqR03
2Kr6+o8OMQ8iSOzrj00s4+ASeicE/BTUclq+gWAKTqJ58h4tPJRS3fjVRHySCL5s710tkUGxilup
PfTKwwSxBqw7HlX0xpd3/EmnmdmzIxdDWEjjetb1rgwJGg4cXcPVfwF8LLdAAFEBV6OvKdz569Rr
2nDG0WMB5xHJML6CnM50fFzsWnvBdEYYKI8S0uSTWO2X5WiWd+AFKag+ky/112uNXFSJfBDgLw4Y
snA+G7i8ehD5y/HaPL/WnSLTO6/CDk2eVFRbQdAtuJ/RjGD6a2Atoe6A34Axgggt7cA4ZGk2pa3w
9aRfMPafkaHxbQ+fjnnDVwB+fVLYVSzGqCzW1xJjsy9IKnvLtV3N3esN4k37IbztV4a4R8OYsPWb
uOkT51IAtOCWNx9wuJt30tpD4NrPiUcMyj9ifRGzfFBaqhtyIBW7qxpSIF6kQsICw3Dv2hiZzG6k
tWAnAPz1aktzJ6aSsRHJgJU6FCnFv466mVLCVWK8KgmSdwaDstlH9baYm+eHwEovt2Y+aSLcWpwr
V2SB8DxLLJ/wjOggkttO2j2xLnDRPrflBwq4grO4c9JRXx5wT0htewu+LlRcGykc0tYsrtj5VrqM
2I4Sel4Y3DRuYA0g8QOf+c87rMiy6Lv4vY/6mhSr/FzaHJD9P+9iy9tYxz4bbTmp75HT29rAm+C6
0pSNnKhNcFUhLbzrT8xf1f92QolyWtS5iEAFRgn+86OaoY1YU3czuRCrPGlknLDnA4CHtBPUhESu
vqPFpk08Tk86Jr8LZ6wvDNfm0vKIz6o2LmCeINSSGydXax5oPvdpnVAG7hROeNlz8X7OvnTUKybL
+Q3Y3yA8zRnrzU2Z6Ck4PmtPPifNtsDIW+m479nzQJNtUYlzyff6aw5evfryRFxcChiE5ZVyj+zk
1APFU+Ar6gcIEJZ6BjwtLY0V49MvFCeRYNK2nVT1eJIjZY9Vrfi1gV/X8kqCjrezFO9aCLI5MM9/
Y0ece06oMAmburXjFFAy+7zw4H9o69rwca5yxqb4JpB0In/s/5420hcNk5BOIt7mUNUZIdUAZ2zB
rxVyo6HVVjAdhIExfufLQiwlzfiNK9W4aST6ILomTPotYBxk2HMAIVbEdunv4oJopgMtxThowi2H
XEtSnVggUOjy6EG7RfrS6mImg9XBJpgfNMVdWPzXPkzgwiT11H+d97QbQfwFSqM2z3Azrmf2fdIS
Nvmc1U0rhVl0N1GoYLkG2Vf3st5P7xCjmohyRBah7LxCqTshwOUfKYe+X2msUt7y87MJiEzMgAxa
8MBD5UC1W7Fu3slBhekAeWLaII2C+i9Q1Bi1/6Rw0tZ/kaEe36n+zRSnWsLKzTSaSXK369fmqoQd
5PEzuaLRvB3H3I26+E7DN818MTryaOId60EvRCGeYVVssYUc/J8eLH1GrQer3+2nmoAzZ+bQjCwj
OkRo/0Oy94glP0FY49Ym2JeGQ3xjC+OswB2J41DdzGJkNdn7dy2kMoYgrhm1OyPCyMYDkqjX5Crd
eWnxL3zwITFgE7smCEC4vSAKs3V79VLt7MPIxjaoSvZpLVkE9nKzsHA8UO7tu/+EV1kekiE/miOf
1jVdOey09JZV2za5frwXxwd97ZRIJ+QRGhTvyvS2QU/li6dFEYYEfN2eGptAqG/50DoeI73w0knI
jYohibu5jbH6gYDh07MAny7lDZLX0Wtba8JLJHAyNrJf167sX6+8Q/9YRx5kMzU6EPtm0bEgE60M
G2dQsab2jDrudB/V66C1xDtMLR3HHn0Zq1ZGcXuqxi9ARWekzAcORSutUmnbjkGyUdYXqcCkUTjM
eVMJVpmCczNLE1w/LYFPUBleK4LwyK/DBBmsjBvR6BVpK1JZoChlrJZwUuBmB8Yb5hzIFsSmqryX
r2AFDFM53ohLKljQrrzEUAFCFx9irW2hDnRLh9QjZFeHPnXZB99wJenVt50DXrdDKuo3KpGnpcD2
8EhXEn9jV7fdbAqwATmZnxUJNoYxnOGU03jyPO7w9f+odZBkRwHbLdC1n2syCn+xi4cIRs96rpcx
YIinB5oSD9emXGDp07FMMePfKZKXnHRrOyYqi18vBtOFBiyCZ3lV699pWqUBKcrB7YOKXn0KwQG6
LhMVrE7TBY895IsXOpzxr7E4UhcTmrWOBlAORl5ptjoIUpPqCNqPKG8LrGnMw6zjV4Vv4l2pKFTR
U0HThv3sOWzm7oY+ZqaWUHiNuJS18mevAEF9a1RhOYiIT/d3kwYkyiKuXYpeQbCnfHygvLWT7V94
cP78oUAeNsOcQT9weoHqG8ebBzpw+4NBtO8YwKDHmBxd7LNplgAYL2Jy86g8/hr5pQIo8e4PpXZu
rc4GwOgZYYarCjOH5CtsId188nOx8gev2QE6yC9pYeLnLU5plZLXaelKbRqd4ie3CIM40FxlGZbQ
kLtIaEdGNat/FJaTNAkWYvbNrtyNE1APsB0/w7hh0zZQI8QtTEBsEw8R8qBpga6MXyNmGNjjWIQD
OKCGTiz//umwqtI/PEW4t+JEPxPyH44tScyfoAD7YxI3ojbWVsKbUURoI34LV+nwqzc1olw2UyuC
rxNiH0/ZxDsYNZ4b8/rOZ53ytjKttN1E90bVMWvQZHry+PN4dpw/fLgoqom40jXNGpMb79jGijVU
eSnmvq6ZVwZ48U79NvrDfJnr7mp45iJhG0S+Anknk227MXAJGR3KMo+bqn466ydicfAkvkFZ+T4a
6g+P3X6BkCvOI0tCahQ0pUyEnu/xovCxf5D9D5hBTRC+oxv9edYPtCFYId/DyVbg18teH8i1RWcj
M5uewKiSjznXMo3Bzgt6evysZ4oGjPXZA8qZWzahlfmNdR0Bl6rDdQfsj0xijqota+4aH9rpmPNY
MoZiT9tX6TCw4HKszmyYg+YvVxwdK8EigSzmGKsRXOuYnRGK6QfBMUfS5gIMgaXFZzYWF82cxyeo
kh349K4d+KAyk6nZQHw8qYf50PaOdDwA/m9yurjjERgNoF0z6CXt7cCfzpkwAtbavsjw52gqeP/Q
ELxTJ3QqowKqboqtkDE6jVlgEKZMXfg8T/nRoDPaHpoRNQlyy5/FZP6vzcqE7tBEQnhSCLjaExho
rX/ulN3zcBrXdBpq2S9E4i83xJnE9fJJf+qDZQJazDm+lideL1/HsfBJ3vxVJD1/0bVmn/7eDTru
8oE+XlTaBM4JFGp6bBNTE4q5tl2bTXmlz3UJrc4hPtxUw1C+f17XyZXEIOHxz5RkrX/4oayHP+tn
7dEOYXQCwSeAXpRAa9UynFAzlkZjXeUWJLJR+QhVT3cl862KPxcMG3MMZo44c+OgIVG8B7VCZ6P0
kwEzfQDEVfnviAe+ATMzpn3sj6I4e5TvxPjsecI9Xd/VWno8J0mfzrU5VNCMtmK/hv8ldfD284ZF
zyhE+HI8nXagq+JdS4hah6NkRSCyG7H+52nCRvRfKXmwpQUkNNeHFCKIVFySizCaYLUbJstXlZ/d
OpXjctdgFXtYip44nQsA5zZQJAEZppJ7E/1pJBdOM+BRRJy09hMoWXMWhZ4M2FwajVwJgwGDn+QZ
7U/eGIC+ZVYH3awScgB1pCKNK077IV3iQZsrur3QUF3ZlmkA43CoM6OHKOXAcRr0mykMhgygNlwN
76VNv3u+K4yM1wbTxWIeFqgZdZANWrFGNyCUnxQTvJYm3L2odPU0QFNQB00jcCjsTeBWvXHyGHaa
2ZO1YF6sBRi7vfCEIYtDmmBZcNerK7y8NQvpCQNiG4IDC8nd3e/XntRzWZezZ3fJMKqFPQB8MHW/
oCHSH6zRDYV7+96sGqJzOG/K3UtMzXJDH/mAPQXrgW0tu8WQjXnyJnCdsDpUIjHXCqbamJtQUe84
LXbWSEG2wbGzfYmkMU6lK9VLcvp36oFpxWI0f5hZK2IlO3RclUxyFGCBOk9RAN+gRnvGe/VaBYlL
AfYNFeLTeY9j1CmYPBUwTXsuMayxQNiLc1I9hPOGMn/251WuE++jtPinqFB+bqKSt/IDc6T23m3F
sefeGUROaLRUoKaP8RQk9MGCMYgTPTZwgrPiuDcV6T2I1MY/9sDpTzXCXFooNt+u1cpA7jf3x5mW
E3tYeSuTWi11zjDg0qQPUnWx/B9ZhJQ7N7hz6BAi0bcSShJLt+hHZYROxVddlD6Z79MgpZU6XFmN
GexTnuHp1j9LBW+2Qgt05rkWbk9AAfs330+dqg+g/+3GbS5G5YcUG5tFRWr+TTBnG0dQNZCm2p/S
EkfKBgZJPNFjxj4KsPrreAHKCRrx2AAgNdgppG2pyUZr0x9zFS/T9ujmX9Igpcu6iGTDFBDt3Tjy
iEWLYIYdUDGlhTSm3a8m2YZ89wMj+PY1RghXMmCe4Luni4TQA+wQ8i4lA06Wm8zd4wc0acitcoPW
zqGw4FBoPWbIfYiiyTcKtEs748VLjAXjueBQRNQo23upI86DfQYfPFaucNWvzOTwLO6kULfO3+H1
aizmXezuPCoHrIsS8EqvyVezZKHSqD52UbE7BhNKKzms0BO+w3p0HbWy7fVWfKc2SYbmQ2aYFErM
94Ls9HYd4cXiTUST0DULshfY5xcCUAjdLCITwwaGMfj3kwkm+Avxx6dPYEYkDe3i9ggnI0OHy/0x
DRXYpIb+w1NhovSvZXHvzcS3VmBhws65LzoLZR5gIo4DJNGsrlV/6g66ovGEj68TI4fMdjGsUMjJ
x7CXmSotcddHd2zidOLweLb05B+XPGGiGQVq8uwM3dI/IG/s8X6zSZOIs3mxknid2fNapUDMorkY
i5u3NvhZLbpxKn4CqAQB6BreOMJqhSBFeeiJIBVsng6rRco/DMkWYCRPxE/2J0ZFBTH5IaUXTNTd
FqI6f0QyP1IGYOzBBePkbXEt+D/M9232nGIt9pQVN4L55CZzmCEnNUa2nq1uYit/V+B8/FN7x9MS
RJiAKudtbBy2ksTmBt0rl2im9WI0tpe3raW65VgFBTCb7rfvnvcWTjSNOBQ86yRPo4bQgQKZGXsV
bN/3HJmtGTUYOoa1Pi/J6HF11qhcdWRD3RDRz4HpV7ojjmZUSmOkCEq85/9W0f3BBAflJKOY3YOJ
O6g1B5fzwpSKBdU1FleQ80G+A/nS58BlJ/Fcl3SI+lof4OqnaOXa29hi5hWMnid3nQXHR4wfEzTa
ibP8lEq5DEQE+tqiQUMNLeRzJpwwN04GMyr5bGn4NeZ7jtZv+Bf+YF33zft5cbVSenafYYpFFQ9r
GUyT/CtfZBLbN47c2xH4Qa4ihObhjMxCAcxL48RtwlkTvRlAN+kg1K26CC6ClOp3p610qLTD4qbd
9ylvbB+TGU/7xC3VpwwyDRYcnq9prBgoDELxDXDkkOR4oTe1jTY2I6Jh8BQr8NZ/7q9biAykn0l4
56tNoJvBWa1xlwO4jWNY2oGKcMxE8LwyYYoHmQ6gWySD1/NmEJwSwFS09WdZH3REpuC21SFl3EQg
HZfwBuMK6+rWeUVlr6R3uaEmh2cPq6++dKFEJZYLUGJOrMSfpxx+CQAOyVESszu7H67BieZ6dXHA
SQ57+xX5T8KJ+JSKIonOCH5yMh3UNpcFbqGDxq+wDEgMkL+BJVZQZajgmDmkMBIbNfAhHcsRYG9r
0ThAy7mGGsRW2f8W/n8Molf/sVu45TMusM7Zjs1Uh1YZ1QwpY1rUL3PspyVQmjI6+SOOztb8+wrq
AS5XDrXZqUlG/Pb9qceaLfveUmcqQDpmARHlRPC3P6JiM/vQ6yXq+FCOdIPb7VYOY4cHXs4D1vUR
fgbkHttFwkkTxexfXmztDDFfPyQvEO2Md3F9PQDx9KuWh4/87XqT+nhexCMLtc4RwJPGVjjCnVvB
/m8DUICCort2dxLDjUNzk9vbLX4cwa2LwdtceNtb+AmL4Y1bF8moBttMeo1a+b3frzgmsfgl9XRo
/C5v84OfFYsgQHC8fBQRN35/mfJ3ZZJefAVK6v5nc0n41nyGtoriv8MJ8qzjzaAWmDKkZ4ZEA3OB
c8+pZ3gAD+nITIOP3TD26FCaSiOmWdjQ0MnIJABx9ov2vn9+QbkZ1h7ZkrKYlbRBWX/khjNiV+ff
EqRbUHwy7s9mCnf0xB6AvfG/ALcu2t/1uZMOT90xMojA5QwZhyPv7M7KY/fYplvIp3FC/JS0TOa6
rM7QtJKt5VhaGppc4h2uLGpLqEz5uzCom8xDaAfM7KGtMQXlnivWElvfjMSCf1B1sgQcNp3ElWou
5UC/uAGBLZAobPO0Uf+vuF6+9tDbpPyaFiq3uQhDtO4tfy8ZRUO4yOxF7UNZ11mqd75n6rM7DGRS
rVtYdA5EwEah7Xi/VsAvqVPuFVYvmNY1qFYsgUkZRAzCLcvdoDUSpkD6LRA31EU0FSAAmiPe7gon
NgDVlZjk8VdubsLRKCayG0amYKu0DxT4BDaMf/uImFSSoDooVo+mYbjP8OH/VE9srUfI7o5mvrJS
ysDEqh/eHHytKxWGHVa3PQ9Tpt86u4+35s5JfzhbN/RhYr8RbLTpJOJ/ZEVDzqpa+vQo1RquwpXG
bsKwV18AUGStYGIwDr9TP3YgRsedcQY8RrED+RoIu7mEZfc82VMGth/NwwvwwpVKzFAEWRsl9I3v
0/SZi13ck8tcGfNslEX+sIjA3kfW/5MT1qnr2ZEjjxgT2mbmlE59R/4OJ8dDrTskhpBA+3T9xGuN
6Q2OOCpNnSND11oMbb6VyfDMGYVqtdnSGBZdW9cilRzBc+R0E0bxWX1tKMsrUwGhHeiuvfoSIVtf
qGjRwuFRWDdkrlyaiayWykEofhvp/MewVkaWWCVt6pnJnqpfwKbJ5qJ51Z1M5rVvlPbp/gQyvUSx
ZewyFbWClGpQDroy0ryDC6RKff+p/pCXCzxFE1kxITTi5CFhWG8z4Ma2S7S/pa2GrI3MkZVXSX/c
+NBxBqhOnMfNYlYEJBoE1WgIiRSny/pGJtYZySrKX0/3fhf+DERddcwlZT3tOTjmGweegZFPwEhi
ARc7pMM5IjpbcspJxAdUcsrxSaJ8e8MxljeCq59edU5ZnFXu2psndDBSMRWUu9S4gCuwmZL6eSS5
Vs/+ht3dFI9p0kWyEyd4m15AERRhaIMYzhJNjmHr+OKRYRfoi+Z2gmg+m7HUXrevrniMBVKfq7j3
RwKi07nY+1hNQhgdgYjoaLyW72Lx1LXH267ru0O6hor1W6YUi1zD9QtHSv1b3u3h7H+YNRZPGUiX
IK3XImqsx2UE9Ko/0BcfgMIWWTxJQoCSPOB2f7WwVa05tjzD+f1H8+tp/7nFrDxo8+LQ42xM2Oj+
zqrOj/ctoMGzEka8Z5DSIzVU7quI1yFb1qwONZzRhCbqe2pOPv4qxtbIlLcGWJ84kr/t7YZqHP0P
UdGaXrn9FUm5FkNvtJdS0v+qV96u2yoj6YXf2tkcOjrAyXUVO4uFGl/85GjF7KRjtXzAC9P9BG4J
5nj8WxgBnZBDzYDqiBcjzNy+CzulYiTKamwFY3m20rn2lH7PyUJSNRnFnpJeuZTjET3XeVeicks8
DYtjjAqvS5k6dN5gzgMa8zAsQ36LpblpMb/YQTRT8oJT9btTlWw5YosT+aOa8fmBU7nKTeJ3C8Ak
xTfSXnxdoB5UV3p7VLAXhaDkbRlieVkNU/tPNfqbnaq5jZw8UXSBp+Qc2VPd5ZPlRbe3FajvxXk5
Bin1QtJHK7m/iu3iwxhbHqvqdZnCHhnlAXRUGNUcqizFxr/X/4sksUJF+AqAQ93PONruQRSAsEdh
R8BbDyDPQU7WLXAU/7FVGMgTHPAmFs9mDXOlmEINs5dFWq0hKSJ0+5sRfPymb1dweo7n2gmErIBs
dY8REwS0taCzNGz3unDAcUAE8hv3uT6JptY4nb+hgvpc9Ft5PkOzHnNOhSdW2ECO8PHTamjckECQ
OB0bBF88YNKEjDFhMn9EBg59avSFIbnwnDCRx1QYDOh8U7oxgzCTsawbVwgGxi3MnNkwPUrgbYQr
xxXilWBBFj+D9rW4k0xV2PgcRHblePU77PC0x5NC+Nwpbq/erjkOMlOxJmkKZG1drl5gMxk4uHS3
9JCIihTh63NO040Jo+3hKIZKhp9r3BsSyb+w7cpHQQ3ch7ssl+FNlR21YWtsQV06EnbWzcYw/ade
20MSLaXgZdFXSP4LeuP+SVs1XgwQCs4mllC6YRHN3mt7rMBcXsYTkg5ID77B+QeIOBN70QVSfyWc
UEN+6fMFsZprNsY4F3hE5UeMaxmr5rFVN4rWZOduX5l+LLTPYA4I88qMVadnMpCw25EyJmbIDdjs
WkvpNoE8OrpnujtI1fXbDkj/0nWKou9/7Y9AWV2T75059mIvXYanl+YRPtu3bQrSRXwMJ4vekeeX
KJY5R6EQ9eP46Tihx+u1jSH8/Yb10mFKX1XTqgImgUtwYKRDpgSZSI9gdrews/a3WLOt6hIkJG3+
Z6tSM7Ji+3d9GBKLVYQzyXLUKVdRkfYcI+NEC7hRNAb6yYnD0wgK+KdwyOXHJMDk1VfrYGV2apJH
foTyx/4NBdgBxK3k1hfT9bsMTUE1NOK6yZYUnT6YwOisgGYafkK+i9Dfep3vKglJAxpEK6qqZvIH
Q9A6FZtnxQi/VvUkCMwkC/NO5TDjOGx6YRT3jHQGMmm2F03lqnbgYFhrMcQf2AIzUOJ/f0chN2st
BMnusmSD8JBXp4qHubq2Kq4v58umriT9Zm7K569x0Djuxc5SeVaNoAK24HBAQLW824QWVyrQTiab
peksLMknldzTETsg0QXZALE+CHbT7x6HP8gI82NopytJbPmnlUtPuPWYLsWNjpcdmBJhjbNlJYsR
IYToTYtCebbTkaYxusX7MoJbbIAyUse33N87b1XSLL9V5HHLtYpNjC25q3yi6CgkP4jk5bVUjnBA
ftMGTrz5QdIs63w9xcgo3WpOwMdWcP7K9kZaEI5lRwu8cclH+SHrUkeZLugglEOQ+qJJ1xgV71bJ
2sssh12LYDAwnL8jvSuR6CL3T/WgVoL7iIT7jobLmcy/Q5Urq+ZDExfK+6WGsxmOsOQpdDIdIaF7
jRyqU1Aj90ojhHltYCHUsutSzSBWbYbBIyl4AjpkEtNDKoGNUe0FQ4sIRq+QXRZvQo/rM4eIswg4
SqArvy9amev6+q0I+Ho9eEh/r1DbqDYa/tO1Ds8F5uAX+jWk5bNE4CvvN7q7VsuM/IPIi83JFyMg
w3anXsvHP7MNQrv8EY2IQzWx5skUeqYBNExI9pQBI/kuKj/+xHKfHiiDq/MvZMRmglh3kfghu/XN
y5jzZX7VUPYDkryHaONC7VImU+A45p/gc9CYEyqYuuOn/JqN04lHxoX0JuyJfBQSPK7Q27TaFgWc
DmaLOUZGHGRzZLGCs3VmOO6U8DCoSu2luDoRGOlZb+B0EkvT3ZAdLkyBqHetFpvrzSqHGvzYfU53
IWh+/KTeKOmOTdtMVqJig4l2bcmTJDfHA9Shdcgd3g2wSzEvhIkqi/F/+rEp0mpYJwKgv2D3Zg4K
v7wU4iD3ff98jeZBx0CEGlGFhpYhKDeZHtgmEqbKzuI8QH95ymh7629gr2kWq4lef1tDAODVdJlk
dTo7BOuYO3FmmBaHAkdEsMWlSZ0It9m53LZK3ogRd95lCuh7PpQTJ4jh3Bb+VeGjMhw4I6WdW+MG
FOJPSUoRL6vBOFX5rwb32UtNaJwfRxu+K18X58evx8OTtPc8Ell6EOqbjn/Yewl0E0/zxLDNYP6Y
+oKayygTw7d8NTsOKIEDLIIqx51k2VopfrSdAjCiT6QsySpdM+/keYTQ8jl4ihAm4QnmCVxnnm6W
zZtvFZDYymzZpYK/5M4RrXfyk5xdP+99B4D/4trBf/C+VDq2UTf2Zg3Yeji/J4SnZ3vphvnfDB99
OknIN8g+HSk5JIbsVoo230n+04gfGNm1O/MKoP9zvdULC17AJzAZQ6/AXJ6bCzp1gUBibmhHlOYh
e60iOCE6U+xSU5JhudwjNx4NnDFd+rJ1307kq+jMYlGvvXy/WDfsLu7P83hVeC4HVwJ/tYCgsgal
aXehGwdrRgZvqDdVxgFqbTL6Gtu3tqojJ8Q/C1oUqDRWJ3Ci129jEbPXV8gGZPC2rqGPQ1mKxPZj
8iKfysgiNwnVXdwfCaneldL9ro5/IiJZ07xW+si2zYnS7CGozr5MRiELZgAzOcXASIsqcu3yB/6w
Jmn5qcXhKrGodijr97ek4u8oKYp5w2GKLI2HioPdODBm0nM9bAeKzRg6VDtGQ5IGZTftkOAjucrq
Df/sq9GQaMEVgnA7GdDZl9lSVDSF3MVaqO/FBX21gTPRYHeHS7S/EZgSJsCCekX1SfxdRsvzfoZX
SCfhEN6HDaHVtHrJXkF2YmX3C5UUJ5w8wZ4P0ihOr9l6vTV8D9chmEUG9c/qKPeSFeheS4t9d/kX
qEkBB+qJ/5RGqCjJcBGiWyoBwh9w+NSjSdrsXFwq+9is5DkY/zD/lMblk+LNiJKGAQSXOuGzALGV
CX5lD6Co60dAV2d8pnMjdQaNbUPydlBJWydJuC+/+4ElwnaVkUUK6RzBL+kzXLyU4u/DlUHG7e5+
BcPrNR2W2Zv6WuHrnv665dEgO0KQzwBO7Bv9u+JZnmWMnPc+4colD2WAlYkyO3pJbD63S/dfCzUs
V79zDdZZAhk1OKETIPmOPRrf4TIgGcwREAslTYEr+HpTMYMjPgWLVVZigKNRe4rTDchfqGCJeTIz
Vuhv1bBFreHpCWqIelYmh+rPuUsA4mgzZAD1tVpBHlWChH6dbnXfj2xJr++Z1RhJg17nfjS7Fzca
WQ9eZyLNR19J9rnETV/e/Ra3DYVFiYuKTW1xt8CDKVwptc5ULTPBhHuBbIDKEfnXSOyAYMc0WN8E
aZPnjGUQadBcIIMuPI3tjt2khVcV9atqrmZzkBazwEOB/iUi0bfejFwCC3nBCtqcH/UQ5VTmsa4a
bkuldRVAwDUAD4KRHKUMcb4Qkms7TfPuu5mirvHTO8y9KIj+BqgJk/cioIgjjq2IpXaLOPsiwP+r
yghaR3R8RuAVlmN7dAdAUsVTwTscym1BBmv/sS0IJRN8hN3nsT/p9+wOeHPcX/sPapHX3xMiPBm/
R5iWiCg08DIVD3y9dfsUv7YfZrMIqWm+x3Wz1n9ZUSsyyfSeBoC5c7Ftf+bPADdkrVtf94AfOPWC
a8DyJMgITHsh07vCRuMxGduRHJeDzo/bmFMOb1s2lxRI5a7W5RmO2x9gNgSS5OiLrTflOutWyv8F
10tSSzr+jeJHtdM795tqPMbzb8x3LZvFT+e/5vInHrRSwt3gSnlbVZ+MsmtKQhWsHPz7rb5wVq2w
PdSgM2zQ4FMxqrtk1Iy3hrV+pSWXOAchrgnDxwqrHB0QUvntIk3j1wCKg87gbvrzatjYKBYLKOJz
LsgrANR9DQK2+WmUjq0KKhXhaFj0jS9Qb3uKEL+dbS7A3tWKkifX2tz72x8ufHcPTjn0vuL0Em+7
dUCxW7S5I5eJiAeG1qQ8UuOA4+eign/bGZL+WunINUmlRIv0TKcu/JilXKjRklfZfBcQjuuNbjga
z30q/DVQCat7w3mLrXEyQtLX6RkYn4G4P4G13tGfXzmky6lSaNXSZTLhxsiI7pOQOoFnRWHFtXgu
10Vjd9hRfLmwH+uNBSOg+3oQ6PxGxkRS5mkclxBl2gWaRB4Wm+NwJEKJp1p9LouWcUp0UYHUDDOq
C5wxz9EhXs3fWBK6pU1GAsN1lXlyV4nJTSFYEeHLiRL3nMLLE7SBV5eUgP8nnGOS4qoBt4Nw0TIl
Nd4d/+Upm3anox0/8pxngGqPQbBdT2VzulnhBv541HhPol1fGbNg7W9+h+1R6BhAPRJROCj9QQUz
9oXQ0Uzxj61G4YSiWMzwNleqg6kHRbo2rDNzoFM+3HVxqnkClxZMuamZTEjT1q5WHjddQApxc0V1
6R9EqImgOHXTvAwJ0Rx3JBuGTUsMA+ckNhIelTrKXJs9081PhaNqKPQ4Fsg+dOEUTXUdWOjdcuoK
iGPnUxcctAGI7QfwPC/3rzoGNKcyKHZSS92B9TP/bJ8TJJGjNiMSxLO9fzKs45XNm+4jAnD2RuC5
tkyYBbxi2q1+JRm+aAytsJ3LvGJDRjgwbS8KP2Mne01gtgxzEQsCWYch1IjF4SG/3oarOzyRGuf1
0BVsTGR++TsrOK6DoOzX0OyOFnEINRaL/bf71SGLVA2zoLPLilu4m1qViuQwZ+vq4kFGt17ik+If
JUDrlBjT2laG6NJNvdZZgkGHPLfc69S7GBQCEY31a3Db9y1BhsLkATFScJsjJVekxh/oeIwOPIR4
uWrWMXWI5Xyf1WfVQIJE8sb8SVM7+9EA7nTsLMrcHGeQyK+0MTDiFSesBJ0IZer1eMdVnZk5FZmN
aBOf72WR2OJg5vvhqe5x0DP8MNcthkKOYPuG0LmJN7jxXR5Q3LB9ebnLQBNzC1NPoO/YiE0LHeOL
hMrcC+gxBamNCI1zgB5QDJq0xsP8tg+sCvflHAGoinUFtvQvZNgwWM1AHBdInGJZ8BKl9VmG7K+S
CpXgFmX+e/oy8iOJvHlkzzKiNAvlRZo800DVfp2tniE1uDJpiimtTj5KlayJnS3CmdFwcNyHQwWD
N4lzXi9E1gVZc17+i+OZ7hoGQiVkO8eetXv6v/ToYEJklqSh/vP+d/TG2gTx1tdPPL/t35jD6RQb
qP3gH/xLc/sFOTWZQtssN8J4WLkEnOE2e5LWAnWblXO6wMKqo5OXLdsgolt4HUc98DQQg25sikA9
Sge+jayjcxTX8pyd6ryxmuazQl0ogRrvFWl3Fc4hbYQakwBtBtyjZKZGF0rmYw2N2aelzkXFr+rT
LMsW1ouEs5f9f2lBRN+O4djB7iDnblf3O4jmg9VXtfZSPNHxPFp0nIgixvz18n0cW+CbyyJTLqiA
OuaFK4WkeuQuxgEVcMJWGPVTkNURNlhtinqLJRtcWEAt2wFRRvUgAwLytydmXTo9x5fY5bf3zJuj
F4HWomeZ3cqoVL46vLW9tdzRBXASSXhOgQ86fUVH68XNcWrWBRl9lYXX9QeleDiibDptYbR2P4Fw
Zjx692TNaicKfDGjq3B97ydkHzwqb8jtRCMk55GzUwXiJLxDMcyyHK0wSum8yswJp1b9krZEN9xT
oLyj9oltL6bNFRk88nywbUF1iKAS+t1pYNw/l3EU8ksxbS7B+LVONq5y3yOmmJCB9Ip+iuELSdru
eZSaogGtJm1JqgOexPbMlArm1QUb0d0+FC8De2l6UNrNtJpugPJb5tCNc5EBO/zichW7M0oKj/dk
f6xyHjby8J9GJvS3y9r2Agb6YbFDC7BrNStZTFr7Fghu+hzXlBbGIrLkq7y048mG6wZ8mbSbhLkW
N4522atfrWiLIp/RKSE+o2qj9GRk4UItskMGgpHLpfuSVGD1EWl4jNOcYjn5zMMC5VrJuP/KuxuK
uhAJ8syS2GwLxzjSaAVGOKOF2SXHOlU1sTAVdmV8LDZ5sySNR1R0Mt10nlx+4qR0fsvMeG6CrVd3
G65susR6fe6QuS0GZjr6ifHF5cMhJjORjDBwnEmZka/Tb6KupyW8UpFz76Jsy5s1KVW98XbAlbGK
xSHztxqOoesPj4GER3GHdSwKDpf27LQWDh/cD79vbVf602XkQq6Lrve5ZvdIJNAlPg0xgQBJnhof
BK9SIPKtWQXWn8eKf7AC+geBI4+Ie1nhTg0FuyQ0NBQpbEP3O2KVDPX8QWBAqcudV7UHQommtE4I
FcFQMOF1OZ0CUiQBxUQ4J6UkcswIkd3I3/Txzp5H7p+k3V30DfBK6fNFhVGlvveaMZFIo15XoUhY
CjLCt1b5BeeJonrVB1XLiYrhUu+9rj2KCHUvBfxUttpQ+VoucMq8WBPgXxsCmC00seNlLHSsQImq
lltTFnTHNXmAHiEZO/7Bu21dE+2bdmF8O0Awqx08EIxNdHxLlTunVP+rQvPeOZwyEfZefS4Fzm0q
n/yBrsC2s6TgekCKBRPtRts8+y+23cL7jaECuTXih0LB7lIe6UhkIU+WziG6y4CAPWoQ8eIv3A8z
RXMubOFfHVowTs8EDwjEFfmRpqCIKd1HJi5OV2ma1Tlemc0BJokv/m9DDFOEgE3JglG5b4xQ89WV
CVY855eP4iJLFfmJP3oV49AuzRlQBnQKHy567eGv65hrtBOHnchagLNJ4LAi4J8EXHejZnNyLTyx
8va6CjfJO47wcjB86Fni8PEaULaqX2t9QtdhCgMh6W9aGXCEBGNewKE5CG1tBg/vetdSyTub8zSm
f1+HVWIa8eqIeO7/ohbcIjp9KimJK5C5/qZFl917ZqI3loboQ5Aymg8TIMVKLxpEAGB9xUzOF7/d
88y5FF51NNEgGDK0geRbENJOcRXwl8WvVBR5scxq2GT8KFSrE9LTQWi5ov3C5IA9dScyI6ILSu6L
SCudSE1tCzqkkiSGL/fApSr+tILHFu4D8hXqOLJ0xG7TP7/ZaCaJsLBXvMbTefIl6LeulNJOVuax
biTOB9hDO3L+rxjOLMi01O3/id/TH7hdFv0G9xlc9fGx5mUA0EG+rbQVXxsMmYRK+fMT4lTxkpWa
KhW0EX6jkNF0aY204i0WH5kM8UsvJY7Iel8NiZLGAxQ1vT9s/Cx4Xu93sknWw8LR5BqJ/2N0FunN
q4f63hdIzJibV3H6QniA9w/MB5JypXCUBtroo+W5beODfq8wkxozK0oYa/tlu1XlMxbVcatq6nPJ
UeSCeQy5i8I94NLp6ppB22nlRrsyScCogg2/rZnXtWJ9J0RBf7+zReZ5ZyiYSStHYIE6IiywZx5Q
jY8KNF7EsS+7nqumbYmAJKJFmgnwrDRrQrSBbco7K1VO3BgHNKlENCc7jH+4yxSQBiGSsBuPcpVr
M7Wbhs6RMwhtD6L/wB6FQ9L2l7yvP1aKQgz1dA+fGVWEV3pixdMgW0BJ4i0tWqK+UwGwTwppQ1ZV
c7MO61KRhVWDvJ5zRO9P91qvDFK2QOE9oTjmaifNamQo3VJjyUUvAUeOtsmvHLlEkd2UK4VcJCkj
4G8CojUUsI7QqsUoaHLk6QRQHTZlGFXbBLhQHt6iSrwKTARuCKkSfuBbEJMNE6Yo/jO3a5OszyKO
SdPSd09e+QUZVeg5u5eLjexCEZb1o/k+KqMFVYCqCXPmKd8r9ptg/+dipnFTxU5XYJuiWI4RKk6C
Hm+dthZNpg23N4lCgzlZvLigXsFXitMlxMDx0CKkRIgLV/1sfNah0tENiTnDpqwuNnImg2MUtR9S
0TThkztme6Uar61H5t83T2A/ssXBJvQIFqgRSFVwQR+atipjaqPeExAa/hCUq9fZFdV061MW4imG
VtPeCDv2zVj145ZZj1sofGU0Qtb/lI8GHqHzMReEUrD9ypoq3xf54nUjsAOMbRCBXFy6nKUMz8zh
CaRFZOmE5fOkfMm1O8loaXKElDxMDTQoCotpwZyOKPmVKJG29fIKqzSQ3hqjh5bAif2x39snO3dk
TPvEgqtSiEAmziRfjtf+6HD4ls+E+0qEQK6Q2oTMsaI8CBaAlvGfy+urng+o6PgiZrCj7HS4A6rE
Ntg5R6fjaFAevT9kMiMc6GuaRnHIA0NqOUKu5C4WgQjmFr61kJwnErR4Cum75vUHfmudsM6u+82C
nPuOy9Y/SwD80Dj/OUZsFUrXZH4m5odszZWjBjAPkNuomWsZyMJFFFopMd4ha3jFw/vFACJDy04I
2ksbiGNqGS3Bc6tjFzGOD8EfVnxWwCQDoDjgmxx1MWTI4BQWWfUSkCX3bgfLcYbFFpcLYj4R8cEB
5xCuzuqK5KgNqgzZ/FTkJH8Xe70FOUwErJgN+T3HAHDEkB9QEUda5gopXxv8z7InxxxGBMl2xu7C
Gss8Bfz1WEJdnMUWUxXcOVUu02mfeNmY7WFCglRTi7JclJsZgvN1cBnRKEdi38ouZtYsrPdIWKFf
mS1LehLU1ttP+5ffl7wNn8Xl6a2mlUBmjuaskvIpnElssHfrhnPxxCEISRcZXnK1RUR9uAndOv5s
fyde4wrk6i7pXQXtuIJ1f1bHNPWq3AxfpNiznyI308c/G6svHcrY2r8uTLDEvmAL6nwbs8Rh1Ea6
jNyquc8ZqfSSiMb+Mz1QjJLS8OoNoeqqwfReuqep6CFksQizPHWktyu3eG7DAYI1TzQBaYHkUfEX
ur0srCPckChM2UyFsC1XaQcHjS2C0Pg4LOs7WzvZpUrMecn0dCnFE4q5lx2xPUiDR+V2v+lhGNRR
taSYwhddHO9qKJv5Qn+B8VNelMcVzm28KIQThJe6Ubot1a3d5Uk/R9XwzoXvtWE3qA5e/AsZshsI
P7I6j+kIyzc+HvZ2ngqTegqcHxyFhYAYQZk5OW97GfhWMs7YF1SFwCjcC5iWM+NOpG6ulz2lVDSN
VOEUNlBuhFx2/l0C3W09E+LyxK2bax15zTfL71vfJ2G8ucfvBjHTayktKAOrsz2qFv6dQOjtVuyL
k3uveiTnNDHtpeYSrNnvj3fdd41iMKLkNdQ7bVeCVM4l2B+SUTwiiqolep2yB/Y3oT0vbwk7C7vn
K44rrEkdwQTie/sPcVZ63DSei4lAYSIEgUiSUAZDNY4GcpfEv/Lqk3WfV/52KCm+Wk4DfVC5xyF7
4esgGlsn4U/Z+J2gQBNAqYjvI9ngYasaehjw/JqVTFsXLHLyYWBl3kke9cdBeSjscsPM6abjjtd8
K1RqAj0yj+/sOKUQ4Bleqc4lwGkUiiGZYBbCehOwR9vCJrj9ivtTPuI9XRyHp5WqcpPs7mhIgE8D
sMyBb/59ihNxReKdSpqTW2LENe4IK1W9kLGr/zB/Eu56/uPoA0CRumku59G/JV2s1xj39mcjuxFZ
Nz7XF6ZVKHSFgDV4QYOhnw263yOltHtdbFuL7N8rvPF7bKEqpH38VtbA8Cm4tVsMkCAzx/H9sAC+
ZSdXX368y6aH68O0yDNg+3lTP4liiARSQuPfhqhwcGKFi2pno4oZdeljl/3GBtXDUZ8LWn+9/SFO
2tsBPWta+gBG8YwhUsEXzkeXXjLwQ0vMyS/mNLxs2t1KDL5TNRN8Ayt7kV/kxyb/cImE4CkNB9Kg
FVSC5PxPOIEms0jhC7nZnm19xxVJqfU6RoTUfW0+WewE76Sc8cyK+qT94/xW3tlxoEgDRTPny42p
kOon2j2oha/wMdZNcqlzRO5CPwbWjINH8+VqvMuVadn8BaCGTUbA7oL2yJ5HXgJnQAULwhGlYW7w
mmJq/xh7tiQeSA8Wz9Zp07lnjRfn/y+ewzzZsaZn2+OhrKQKB2nFT9TNS/tukwrnUJGpYqUZAdP3
HOKO05wRaOI4fMMD2hOzfAAc8a5+vQHixUaU6BGjsXSIcDvlwnaYyLL52VG1OFELLbRioztj+/zZ
DiChd7shnaLfxqvgzDU5tG7f0A4v0UmZ8UK33uR82dvbTVQxmxqwBFPGiMvmAeZ31+T1a/fswY+E
2Xir6w0ltnZSHFKbeZa34cf23SHeV+gY4hz47+yLumriJEvsPpW98aaQGpTcGgIDPm0Fl3Yj9lb8
4OTBHAzGYAPRLGYemCWpLZmmqwtC08SACz2S5U0gIEH6Gb1Z4T0+8827hs8xkaghRpTfpxIZTTIO
7OKo/7gCPsXjGcnoQ1G8xbK+seZWpATXChSR2P1YrrjMdbO9p7UuqNvvxlbysFK5K5YUyztqfjn8
hHvITSofkGLVMBCt2OZ6YIm1QBXY1WCokpS9mMUi6CBgP+fm2x3hWHSU825fUKwSg7FkMflQRIw4
APz4NPqrLhFPpGY/wlE2rP/zCWS4BbRDNwAvr1NWmCkQEKW+dDr1m6vOmmopLoxgvNZjYSreBGnA
I7EOf1TsBuRAjFjxDc62Qn6lJ0wGWOl/FPtHS/ZLFgwoLuOYERXKVEKg3YlIJcL5HVGRdkPSNFV4
G3veMJJURBqJUQ/WSnp/lX9/MuUqVQWjVOBXqlkRTO85cabh3U0MAcTI8L9hlvYEaZbk1aMowDoi
62qNmjY4JHOdRTTwyCNS9vyDFjWtf+0EF3KAVkC7mdl215cqfMR2Vgf8duTnFVaJ/gz53TjtArZT
11VWoFgEnZb+gEe+6bO1jbe/bMnHJ8WBr3ItCHg4c7Rc2tJKLUGhc0JoIj8o3vma4LfQw49i+mYT
j3Owg/MFiPFdiGs5g8hq/LDM88OKZsKpHZYtigjqHfg/VyCgaHa+CL387pGSQuPhobLBXIY03dRi
9YUb0Nc9ayuMpjX4xegV9DefQCHARlLjranlfpXa9wkHKP9owGtG2ZMywkGS6AIP5X6UiU/gXUWV
cBVA2cLD3lPqyEH8B/udyw0w8hClLjXv5TlWjnJYf/nC9YTEJQwSGP5NrbKhsy0o6BqLQ2vYzD7e
wGczGmsa/7ggmRIbUimnTbxwdIs3dcwwT0oe3zW4EHueSCV8qc6vHxS/fug1PUxu9OuaplUVt7Tq
JSANiuiMF4H5TsbTQFNzbI72tIqh1r8BvObzKowdVntf27yZjFV5zJirYKQRat1NYNG3xOwOLf+H
fVZFfgUf3IINfHrBRz8nEELdELTl/5lShFbJwclHh9ZVpFrWiQL7sefiwdZQ/Zk0PWQTSxph2dlu
wNho9pf3CvKN65KxZ8QqaIx2o6bw7Fai7alYoHVFBauW3KgSBqUp/0+5tYbu3X8dmQAVpl+1Kk1n
Qlq/yvJLBt/QaG4rVoGapE7866h/aoAaBQcc9AFt8z7FLa0O22GM8WfPNomFSO3lKJmwWqO7piia
xgQXv7Rp0yXaqdgSHb9kvfexo/dF90UL/pLpxPoKf1tEjPtXMCjDfvTP0drpqy1/Lkky810GWq8F
x1MvV6IdXqnRNplypBijGVUfZiTFPEJVv5gfrhkrnUG45lpJVrDPI/AK8MJtYCoZIjTasRdJ3+Wc
6u9P23pCIITMdj3Jf5W+CeJh4Z9m47NHrY4UXdekajf3LLi4XyjYTeGXn7I5gd6lR5ZzTEY+EoCn
uYDDO7ZRhsYrul8TWgWTw860KuvWILJAe+mD97517ZO1cojy5FzOpvv4+MKWU13HGt7W6ojOI6a3
O15Es5VT388eKDqEBiKySvjjZV4e4glzy0cFu2VDfIX3WVhKjwtT99QtijerxQV2Cv8IBY/TRXjL
YqLR6RBDI3kHdWW7+wew/XhOmnCR1Se+hVcjGO7gDvbXuffgLvLghewac+I4Y64j2iit3bC25H2Z
rT6F5R2aJc4Nn4anNdw6DGntQH14CKXTQCsRbbP+LHftV/cwJ1J5Fgi0qWqvaay5aPk15yoR4PmY
7Jw8gossy+N195lFsL4uNQM4ltHLaMXde2CPUn37355wTGOQK4dbVsUc+38TESTD3Q6DbTy1wjdq
XelCBDUOZNUxAwVLUbT2a/PpfPQt0a2+Ut0q0FdoLk0TqcVgb/CsDqUTg2tgDtlTTis6Cvny3waI
e6zM8/vcL2n9gHbqQrSfV2lbQJBT0U8oRhdo/dGDRVNfrIc54mTBNDH5Whk8GAt2Vgw9kmbDzvMs
GeMpGJimM5z+DHa36hvSepWNg/UjsS/gxRIP0n5F4tuXDDGZhhq6+KtAjN1MGoULu8Lmq8j966si
SRGVrkA+63PNbjAbq4kXg058YqTFM2w4E1h+o1f5Y0F/MyluDclzGLyaj3mU7/xiVIBkC4+rXo+k
ZucYAIVju6f02w4KtjdV2EfrxZpIq5tXbODx3e5CprF+FKyu1YrxmlKl8fUAq0VQ7UTgclrGplt5
SZctVOFlRm6+N10ljh8RdTt5mF+LeccZZbPAUFQrvxSTT7bUU4edoWNeKy23nOri+dutptrNGd1q
2iBUucarvY2+5Jy3coSJUhZMjw7ZVUfYht2JwId3/MwlaBcEAEd26orQmoTt6gN8xcc1ZcpjG1mw
U00b2KZdIG4WByflFvC5O8vHaePE2ZJO6c0ndmbal4iTvah6/BOKO8GxqW/Wl6282v/ZTmyde8vL
Lygrl2ftI34d4VMwRsqmpOu31OTaH3ZtK4uISb2is2i5WhxZGew/G95TuqzsVcIe7nn2S9h8/RBu
QXmhILEQ5wSifFgVOI0SEB4wbEIfyY8fqOC/Io3SUT9/ojbmigKTtHUo/oHnwERJ6nO16hApbYem
zWLdN9glP8XZCW51FLH/KNEme2lN63Gd+S5QSfcSJbu8rBGzl6imQbKbjZ0tbUFfXNxELgaUv/8i
tC/O2nYzl8muiIQeHpYhfNdyzuLyF4S8Dsm9g2Opo1n/Xn1dV+fTTVFsNn9Zh4Fh9rmesdD77jfd
SSys943zJj0QVItzr8NebSXWbKZcjXHoGRbHj0XAj70ybWu7eb9fedIgXOtSIU0XEi1WSxketvw5
T5tpwqoHwePvbbkFl0V3jkDALWf81Vf9DRZ0BApzLbuHO4oHl6rjVB+mi0OwEhjhUHR28LzLQ/YL
X8JAgqr7C5WMAz36Q371kLmSfB4K5UA2pMImuOVTyTx51wXoMNmLfbDzuCg09NgiBnd06J2tmQAW
Mgcgl05NYRYOIe4KjjpygL1ygpVIWKtrP0g6BvPtH7746k1sdnyfozEBVXhQd7Ecv15KqMxvS7Aq
b+P+4UsAhhz93jwsI7S/C3hpuvtaAWFMP1u6D2pTJNzidf/dpvXE4PwF0daz9FPjxRlxg42t4ZGq
qx6K6lEAO3kIMdJwlFK/q7g7KJKrmW6wTstZF6YZ4je+J23N0lLMfoLa8bTlqIfn3tZBXCZj+16b
8yFLJBfTR2/d/RbmzJK/OzuCDDQyXwjWX9JnXzfZ0ZYidfZpngJjWwscrCGOSM8TzSUhOv21NFJv
Cxy3Ua+RR7z7nX3YaMiwBbOw6kq6IRbuJDxrG0wHKUU/m9r1+wa+4O3fX/7Fcb87bYsyjrypgEpS
w4ikWIqs1Wvp/eHR3FFQ+uJKS3AaM1gXZCBVLSQWJKyRgLLLMij8e6TE73nInIzJ3SK058iy4W3z
fY5O81nE7WkpqtKGczlcNcJTZJliH2PWotexZm5B83KerIv8hkrZ6OWHXiXjJaT29Y886+iyRqR5
ASfKwRNFGnxy9EWpWcCKI7I40zmgv1GviwA6IGHorB/f1xktYnYbhuZMQFQ2N0pEruc61AvB0Zm0
B53Y71se9W2cjSLi7SJ291DtnyxBUXT3ovkDhxZ/eYlF7okKp/S5kI2q44Z/opEX9EfxZ43GE90j
HL09sA0qdxzKzHOShqUfKc2eczo0sUlbpJR/rOqpR4QO4iOQxwHbi1GQDDApcLfWP5JFkR1nz+07
zxKsKEJronbmwKOv3dhkbEod47GQjM3F4f7oEoDza32NEVqyYUOkg2eOo4sJQb6V9CzpLCrDbayL
4Izwqe3t8cwbn550GVGr5hDA1eUIIhJNTtZOLuBUy664mYWEwDjBykw77qtsi86FqPdPe0K9mPzf
4KmpIcocn612lxAWJPD7iYQAdsqPoRBi/lQORGHDFCIkvNsRTfGNv2ktDCsEvC64C+d/TI7QyNgb
hlHsLPcP6XcwvT79Y20K7SuxMr6NTrhF17QybXU8cduQt7nI5jJp2tU8rsVSH7pmt4Ni+BAKNkeo
NbfDTu9ZIgt2bTZl6smYDEPRoo03HUi1j6mgJTpQQfpG+RItEpsAdiz5RrN4fTU2pGhGcip0gVNV
o/SeXu4afKva4vGYGYXknLW45arwiBmkkjd8h6V6ORcACfXvLanfz9RlUE+mbPytSvkBYeUJ/osd
Sr3vtfSCDU872wmjKooh6ozdZlQpAN7v9IWsTIPcqnKyKAoBQwV1WLHNr1U5IiW29RNmTcNrI/vJ
rCHNpwqPXh0INfLH85dXwEFhpjywIa8GJNMqKBl89Dhaw1CmbPgl09imBCJbiYT58fu5zRrjkJ+P
4V6fFQtmiTL/mjovZjPsgYZrKbIrihKKYM1Bzvi+CCoCPUvf6PFwnbVzLrBrwABg/sdy7d6BGJEl
Zxrmisvk+H5SDGjUfkK3gW6HNXeo+qu24Sw9N5xao/N1hgPZZUorAQZz2Ueml/jaZU+bEir6Bfhk
Ys3oGN5eiLySdsxNWacDQE9Cddc4Fte6hGqgxoua4b1mBuylKxTSMORS8RGLwfhBN7OuXn5sHXZa
9egQLhccx7iaDJU1lqpzV/yIZo10/EKMM6xjBDgnCRfERHMAaMn030+PaT1CmgPOurhXlmpbJPIV
tMtkJhXY7Osi/V9zFOO59QCoDIE+y0QZbZI8nYtYcYf3/qIDvW7kQUoC7ifZaRg1DndyFDKuhQQy
vSQzWyDQdxDtHtBw2YJC68+EmtMn0osmSV10rV2umFMTKjLCQOzs6N9FvAR7+itpQ2lyb2XJ5n2N
bM47UXT78QLlVWcF9DSHyKWly2SrguzVCWhG6d7tzpvqXlZSjeO7A2ut1nY+kEHFvB/7SBpFGFPN
ihAQZ5NaynjZojt6SuFCl2pBM2T3egKyzr2Ecb3m3KfSVhNuliBeC6djLmRUQN4dT6KLTmQsMEtn
1cpveyB6Irv1uNX9Er4rvUCWuP0B8Cc7TAnd0261DBD1rr6SICuqjSHg0hvGgUOGqGgYdPpyZGMH
9/bRiiI4ES1JNEZ0Fhl0fLxW6Sg5p70vCPuijOBExb6kIehTFuLFHZ/qOu+hW8ROCXBC9OeDsIfH
tDiOXPnQ7EAS335kNtP+GAjL9noT4h1K9tnJYOYwcUeVvhYiYHKCGEGWFU0wM2hDNerY1DJMIRNt
nbl4x4WbRvf+vrjysuLhXzXjPZygFd+wJoJyBriaJOxDLOgERiUoi97Zu0lHwjq/W3m2nnJPMh8c
dcvck3iR9iJRQiNC/rUsdR10MV5/DWNYqstX/bYFMpD6dXNNAgVhtuYyepJKvY+J9Vmz2WwCujNw
wA6UPdBvcDfgg7v1krEZZOo06XwL5EKFw9LrTg+JyoTLD/7SwtSyYzlY0xuT9PuwxX7BP10TGze8
WYNtPk8EdF4oo9JRKGO9Wii7Ebx7P3gsncC2jc2gdVEzHplXwVHd+x13euYS5lJ9rsJeIcrn9SCB
ea5CFWdyM14fLzolgF+/1a4SgWNjhLxUzSjaoiUsWn3BKrV2NGfxuBl4JJmFgIVdj0DuDHrvs1Z4
G6pGvEAshqaUKi2AnWO3QOkvRNoRjKOq1f3yc85LCLAUUs4kn/pwlXORW9KYR/ISQFYY/Eg9ZQpC
ejX5gPUkdINgbclbpcPRNPoZNI39cdNvWS+ldjCUXatop6y4fTitCCx47cVG8TmDN4WL5ih2hD6+
RRRjBNd19onYyEkVoL5A0IfiXhwUZ9ekA9U911c3RVKfeJoWDtPJM0hGU+7iQcZNYHTgZqNAthhD
1ZzFlnGL57gU0BgxHlwQ3sL6qBCkhZJHlmPzQjVL0wY1TsKVjuhqNSAj5saMtMxkAryWjTwX8clT
1rkd4sc0oy98EBTEVp285lkzcvb+foCol1RLQNdVW9XyPBXmPyg9RHIsRRpVjmqiUPvCp8k7ULvs
ZZaH/8qOQ9aTeNoXgePFFbB1xvhj3lbHl9ujsxmFl/x/glKwDqc602PYd68ubno/FoyV2Bpc9IMG
LETrAiBvJ2PnMW3hlE4iP7TSQK0W/L5Z+9KRnN9xiHFV/7cTx9ZvNgo+UqluHaXaWsUJJbWxWrQe
LOhYzhbUlGu8He6M21xZIlvnt1npTnEddjFE1592a/7c0N0WGdGwgNr4r+KXANQ8sm8wdvVpjCKw
l6wAkI0pwXrbhqHf2egnWEKXXUE2ONBcHFJltBDD1Q+jyjMdb0cCsQhCpje9LO0GXQokuWcPqt6G
XQ+J6ZwB4I0GDVbOKBgEuzkbrM4mhZFSDnAqS3WznmWr76iHhpx3mFGofvFWyC+w+1PweSlTA74b
8J1Is5LC6hCU+sLxFKHpbh5SINVW108aJ3HtNqOHqsQQbS4t4gpYQFc2qtLimU3/DztlDH2oXfaV
UYtibm3eEaPeG1IgDCPrlvcgBf6vLZEP+8e8yAJ+u61l1RIel4yep5m6DMuKgOm/D8V90Tlttb2Z
t0wzJnLzQKHhs6xr4Mlc8kKmpTXV4lY1qXzg1OSmAtPdZb1zLh6pm0Oj14mkcB+s+4aZnLhMgJYL
PV+oppoAptUW53f8oogeLlDxZx4tnnybo3S+78O9H3VdHrBUPoN0ImZi14oy89z91uibhNEKRNJD
HwN0DvtYiyfEFwfp4cyLLkIMrN/30MDg71tTjvAUY6bCiKVtxeADC5R0uKM5GDpE+V7yxjg0qblz
SErRkCAQ5JyB66Q/nZYyL6iy43dNeCEPNMkyj/B/flWL/LgqkBVDs+IO74zMSyPyksRLFsNP2beE
iA+xiLzDV5LgTR2HBRktkeEkb/aapL8oVs48MKojTb7FZGr2t/Il0hMly/93GrCPeeHj/w1JS0/o
zmrQLQAyfi94slMjNuBoCpLNFEqrITb5JbV34wK6zoaZN87UuOW10rDSmo2Qnf+1DZxGcOKgSAjW
IEXfyvC6AqnZXUgaVA6opXTb0TdF7gkxRRMiGocQba3wTZl2/gdhUYwcSpFfNqZg9qwQ2/9qIApJ
5amXO9fzXw01s5T1OcQP495eSclq4izjMrFZsgvA+49hndbEFdNwd1GYz8OytHv4/IcGfUE1yPG9
qAwp830OhEvI8Q1Qf/p3tVuXxsxtFagWYYdCoea2ZKseAzqytTMhixPS746prX+PFzhpJGndk+SK
yRbPcW3TPNUT8ubIkgOMkUdFKoETqwOE1Vq1bUcEuGu587Jfiu0wPy2YUl4aObJ9ncEpf/054xCu
7sObgygqwMjMby+XnIK3pb3iyTmWZ5UXrUk64GiF4B0vJwaXsuNqnhb7x6ux0WaMzFJymZfI+CLk
tHlAKccXQ7oiYz2NrKNAlDcjjQnQSReR06QlGN0vMbxLHR10GfL9jR0lmpFVD27xifm70fmZABHE
RSMR9lhpCoZz7hKEpBb2SZBu92OH35syZnzcRDMHG/YMl6nhaKgQ7vi/ds7zwEwCbfhovfkeE323
zgXvhACwtw2R92iPyRgERFnPEsKCYVlXBaEOFqHc9v4DhnZ2eP3PYmPlUPgQw1IpnyFOErKrZ9uQ
dDvOZkFQ1zyFaLp0zSSkegKOn3wv6U1NHkY4kiy3sjf9lg8FUXCxRE35RtwkHYTLug/faHZhfbxb
QJdyyNkJnPYWGLd53CNPrxQGX603Q92bdYVH9eCSPWfw0gBQnWdFBPSdDbGqK+QXYgrIIjAKvOS6
+ZDWcGgE3lVMsqqjzcMwNUtSoEhwfFmEwUIhj9wWhnYQkHhFxZw7t6nlDFu37sqSzX+qBeu+9F+K
hhYBsRWCX0AvmBdyrUadt63VvYpBNBu2vbhQlvLM257jceuQBqaeesm1xlRPyhzauSiy+X40wOLt
dI3bu2D0a+TI0QB/+8y7x6x34XvkQeiy6plKSCb/Cyemz4t2/vlkcFyYD8fRjr/vjS/Au7rZhgE9
9bP2UONsmV0mbNWdOW9DStJ3WYOQhlIF95fdB8IX+v2ySZz86gpvJ/R5XhCEfNUOfn0ZbKmpaEAR
S+OIDnI0UAeqNbKWvAdUOVnR4cHfd15z6d+xy/rtHJa8xshLYDgBFZS8j8Z595wbnWu/Gro0Yfm2
I/W1HEZMkf/Bi/DHp+CYM0j+V7rXys+I2gUMTZu9NC1y+xwqHz5MtDe5Lal4ZMM1a3fZifE3S7Aj
lhfoKrRZhFYtwQmqbcLYWBCOH7Opb68R/BXtwCYSUiDBPfBJog/7ztEEOpKXlrmKaJPrJdmLrMiS
96la6kLocbZENtAp+JYo0SS3It35zWwPe+L7+owgOOULRnrd+gc+tbHECcxpqrKip6+GxqMfGvDc
WYfbLNJpHy82cUk7DmREhRUjvgDhR+ExpLFGMu/P1GBfj3XN7uBVMFp+axMtZkUZJXtQvJaczO8k
N3OW9jdEmtX8mL9MB34Ivv4eUR5I1+GsJuGk5UYMuaKjLhx81OhmUoEzua14cSxjZKm5+KeBZ2Y8
003YnHlS3iOBsOg/shegusit1Sf/tAid+NePg665zQ3FbWvosJ1SvAqgDG1QxhTaWL10cCietqx1
EDT+TnMI3iByR0jioXFCI3aSsRa0nlG+z50KPodbXijtVcpnwSRgjUEXsIc8sgC7XePK+rMyI17k
vWR83F8zFsA6LObWrKLet5s1BjfSvWVnRXqy5F8YAKl1F4q7AG6x57Js+rtQOLg+QSFWwqjchZyI
z5RF5lbJEOzTf43/gYxZnBUY8k3RttUdCZ6d361Mo28ieu51WXwLDNPFUkNbYZnDKnNXLPefBtuN
OOidGbAY8MIJCZS/VkL+qWyS6roAvMqnfwVlgRL9jcG9nU9c9/fT1QkM6s++LIGiOeM/DgxZ1S6L
Gb5cmPHy636yGB4KnM7udqA9DcuqDcoe21+RaM56i63hprf6MxYUt3qKV8Jilq2l6nBJVup8nUsG
77sUTdK/Bflc1wkB5j/1nE8WxLSQGcmxA9FTTh25hK2aQSYY5hSTNXzdn/cTWB59ziFg0nxlQH31
HJ3ImYH5Uh6OEmVrqAEtrVLNLej6IviM6fujymGM7VJQoNDWQxdBoH8or86rm/tIIvaMBkjXLEjT
6GUlNBTiHIZldu0FmY8Mq0bXscljUmY0sTYqctn+CE8bomIy/lyAIqaQnJhbkrG0wwkVd+3RFbm8
D6qoxb/ECR0YBe3r+FLupZid+wGAovNYHwIQfUUvYLn6ungcUQrr9a/rLMTzotmybF7ECjuvpkDP
F2w7cOidCZ2mquvuXd3Kl7z9ULlPxxaRyiPEavljE5Ji6uuCvPDs0uRsdmFrYQzNtUhqryj8lMpy
CGIHgMEfY79d1ior3z4BwEdrb+vgdaGJV6foP4FDdFUPcSaoL7O+aNRA0cJy6npSYljhgLl076pj
fl2sfKdTolP5x83uoLCksNu5/hrsSt+T4qs+a+q/9qp0N3+CFHb59QhoNtjL2qk/snRHJrAiwNku
S+03RM0kh1OW2dEaM16yELQkzebggIFAfujIxkgwPTVvNFvFuvv0pw8tsstglk22macXrHVHnUda
+h4Z1YG36n+oBwJlv77PZEfwMTllpry7Mt5sgbwwcbHsOx0+3hc2dJw59hGfFUNdxjEypu+XKbmS
mlSPtEdUWU2jyLIu+YAbAA64gL+G3LeVgkCra624i6fRvW0RDE7fJWTChbxajvbPBBDY1acqH0qs
0K3xyMcLRguIYeCc6ThwXorXQ7dZNDGhRjsGGe6QFe2Xep1IYttRw+yD/l8+iW8QBbwaWluAetqq
kDIiDrV6/QiWWSEMD0NLTQnsrn4LfyDc+uMGnyDrZzpNvSWqgfkwsjxj94QbiDO2/9d7GICq8982
7BBsxfS91nFhGtw88BNAA4DXEvcVIfwxHsc+B43QjR5kZRkS+WlniSny6EpZoe4OTHVe6Lt31B2S
Wapbzyk6m//zF3sX1uOWIeURFD5ih0CN3NIKHtc6Q2nfpMAd+n4hwKtlcD4sLoQIZkkf6DP9C7kL
5Rz1L5ADBG+tiBITe21kNP/FXIXHkja4a8wOgdz1Kc+8dC8dnjdnd92a/bZvxSlKX+00Uo8lJA2l
AMslZ9ssdvesOTfiiCd3j8uoNkGKobNOWiWyKQ6iiXdoU/mFWGHFmwbsGUCTeSwxDWk8tv41qpnu
s4VZ0D7P03vvKBdoGfudYHgIy8J0aULUXhvjM4FbTj0n4ptkl/wdQ5b6Bau+onzwu3GvtGFiTFbA
V8J2o8sqLBELIsjjEaKaYl/E3gvVD4y+Dj1xOSjkGJ17DnVG7PiLbYXwJHAc/RVzYFGl1ZJgBMSM
Ixwmd/kcvvfaynvIkSozsuvQ4aOwC459czCptX97fsj4FW79l2rWgZCUN7EyvcSLXeAw3JrvJF9v
KidVs+a9aEPpXd0q8Tv7WWA+G6QwzVKlWxTftrLpsTOadoMNyATG5il+kt/nuePTfbrIM6qKp8Yt
Tf6ShXg60N3bICFoooLX4RvRJTNhBngx5uNlhsmD1D1lSjcaj/5EmSJy3FiNVlc+hupVq8vVqnrE
rnEyBlb1StXwQJsB2p844XXa26EAXYzjU/nYA4rOZIuvGgRnxpLoGPyRJIDwjEqcJtVrK/Sx8Coj
e7nfLMRPGr2DFqog+wMSa6bPPnOoCfzSK2mMaiEnMqC93AMs2X4kIIj/6HDNfIHGZTOkt+iHi/o1
7zbrnk9zWiw39Hphug0r14e/n/kxYTS1xVTu2wwpn3j3/RI4dFHnymNXXgesYCYAOPUhyqTrRnQu
5WsaJkpzIKP09yg611lheoAMu+xSYvd9muhZZunQvbUkq/myEwW3OV+E/sCta2pRJLoPs9vQJgkD
Ey5AVYMBzkpLsrTfk4DJNF03mYmO1fzwZjvRqJ6W/brAj3PMASeqPf9DjtEhThg77eO5uMycTnuo
6EPLkgqhj8utmbK3JiXMnUCHn97ggMeaMkE9I2wZZCdenXje2Bu55miyro6W5bXhcCptGS/dS6XY
DofHOpq2x8Uz9GRFZMHGAr9mSghYkwW1hWMo9VjnLK5/p3hC6Rcl3SDXoRT3fg4VUuqPMEqVUoo9
wP155TjcmczBCjtACtOvY+eeyeZMzKK/cdEVMsDzIRojbQzSq+MOrUYM88tJIYJlvxJOYMJk0wCq
3yV8yuv+m0vRks6VB+k7FRV4c2HXw7rab5Sf6v8YWMo3T/ZUeZWNOxkIf2VMPusQS7b1F3J59M3K
ML2IF/VxrXhhwWMi9Yp754oLSilkTOvCgS0cHbh1HUeGVQcdZmGzu57WSMFLFHXZ/wxvpFXi61j6
gspYtltW4xQELNFoXMIgMOGYA7hY7MdlGYfKJgiKdJOnuFbS5E/zGe2HwyBbTtaf3BbgKS/IOLUe
VWwGxbUYzsoGx3icCkUpQzBRh1Nrq3AUlEYQgGksHp0Nm8pEWjmeu8FGKWdFi8IsBObTlX6fLzD4
MIWkzo/G1DqiJAY1YTVuGbbOvX7ojiMUGWKEs3sPWydZz/Lq/WN9gy7Xu5cftw2SpO8y9BbNHPmN
+9gntv7p+wFUXe5gp/8WWej6z6etWUqxmh16FdFS9dcqDa+qVjCU4HmqQLSMUn9BfVxz064Mds4w
tZWrmVVmuCguD1lUfiIPWX/eZWFDDOGtPVJAy1veiC0Ve5C0VmyM+rz9mgm8w3WU3PyaoEZbu07k
Ge7Ed+uXLygOhwsrZCFGZEGJAA+Y4XEd0MLIXIWw1WlCLGtapLMGbT4UjpfceBqQEwm4G8e6VOrk
lW6CVMI5DLyGAOhnywxt1cO5f+UMkczP72w/1thDdDHNN3f69oLqWufIpOHf0gEEy6KXquf+Npte
dEodb0x7JMoslH6wWgO6uXm1+HdbTA7LFu5hx7cejSZYl6OvGi5OxW6fnADTRnAwE3yrgg9Z/pom
8+5AaUUBoA226DtvAdvrod9sZcPJ3AUFeJRoh6tfAsjv5knmHdzgVYYEBUhqfgVfeaQP1u0ktwmS
tNi7aHjEPNmF+84sOVJsYKoakFhA9zQzkP6DPFqv38gf1hfxQKJTOQG1iYocu4SXmuA8uDA3kH+1
aNxaZf4MIBfVaiwbAgTHWlNlfwHKNxq/XNHb5/LE/riVg6LFW6xOWxEKBIkolvUYwQXrzOFThuwP
+1TetNQ6Y1ij6m56TtBjOo8PpusDZivaHnjCwRWSh4VFpqB7t7Gi3fGb8XuOxVTv7rQMMfQBfVZf
YHdfjlmXIqjtkr7PBITvaGmrtXCyP+mBD9+tdPK4UmG3fpqGNw0hwnpVtl18h9aIhAY7ojNxf7NE
SNXlKgFzREqp5sbvUkdIn0Yu5wysaAav9id8SNHSpt9dp8JvxYP408zT7QbJ0BFlP+9F+DoQmUPp
m055X8vcqJZGHlr3W2MHYne9LtGTFBf36IpZ4jPKmZVvGA9hF25bQCwuQV3uy9ZU8o2H8jdxPKuF
6C6Im7sAXjy6QhEjcMhp7ChE/tqnhl3xHjkul1A9KQBEK9Dg/s2EIcQSJKPfiH8Y+uwezHQ8aqyf
qjdFPImkSDH7TQFmGHmnoJYRpZF2SUYxFvZVMJd0DwhWsDZpe50Q0lrHabLuLwtScgffIOvqPQR4
+vyRdjMd6pqzSS5pHbZAbkO4zbtKbRbdaANDgNZj4qKBScwHBslJsvN+lwzCSd6kQ8gUvNws1U8U
DcfZHJdLy5vYgbi25xEh91bFuNzau59gBJXOZqURuF6wUZmnou6RVYkbV5Sc7pVRG/lfQl2wbwfr
JTEJOaBPTe00EC7ZDimuUwYHVITq2wOhx+GTyc0+UT5ZqHBEHsVRSfJYnYXTxcOPTThJ6Czh8gec
fDVGlF9nRC1F2I7bAH+wnEZWoAYBykLyzFvh7DJjPnFr6D26FhL9c4db2J2V0NhP0BDKYJYus61H
3cneYvPQ+Dvyxr6hKXU3w58iYTVh18zNBRF63FpOZm3hyBJOwjCSNNGW7Zk2fADsMyJIFh4X7Ij2
IflvX/vdvMLE9U6jeER1/KfRBzOchEOE/VaUNy9fyJlEk1GtMMiO98Od4johSyhDsJN4OTT9PPBv
AF+HTRG2B7O72oMJygYQ7IQ15/HfB/N0XAozI/z+HP1oewENH3AFAPvCe/QVgEG/qhfEPtM6W/3H
ephlWYtzgjmPS4WGyAinTgSQKrATG2MmJVF0uqyQOF5Gp0ZYpXRPFvHe36r0yQ5+0OMrOlqhjWu9
l2h47k9+rhMismKDMrshEjAFxRkwI4t5jiGyVLHeSQG/d7o0vkG6i3bFDU27+RR2WH51AEgns4xo
bTbUUivdqJB6+wGdU5ryAWAzlaQd3IzIhWQ3WIFMPeSGDhz7WAAB5nwpCQVvqO2sGtSKugleLVBx
lknGIPflsXffP249SRdPOBJVB8Xw1hWBY2ePJLwO0PBn+l2lRmkK52cHojeSycSLdLzli2Xc6SEi
NvvTDmHuSvGswytQCIXuhteaqJlrAAYc91/DthCwr8GVLEbsx20E0vkzVX4KgXSqQs2Q7G1+Brv7
o7I2qQnHbSx8fzu09BPB7eXmfOHqYwt3yjoIFOqj0bRKqEt5EqalH+7pE66mSwfXROz0vrsG3A5C
IQ2TvVcbQ4FimWN4eHitnY9jdBTEuFlBAA/sdxT17GvJzKjx10QOABEPLVUQdXzFyBsR9BNmBoJU
aQGMR4TgfteSMHRGNG2/XHlS0cgxDxpXkaCrgFQtUAQtFwL7q3SI9ssG5ssjJb8W9vzpBktbd0PM
Mny2N3CMekyRhH6t3mKHrP3eOlUqvNjnIVuH1Zj7nnRNJ7VVFtEPeP+LHXZ9EWPLroafFKKxFCa4
m+CKBg68Z+OiUSakeXKIRo0/sV+qzCZoWayGXFn5tFgruqUUk+ph7Gljr80/hP6GAM+xLRAk3jy5
ctLS0FhhIgXX90m71bLnyvCGEZCS8NUJ0+HXTzo0SnAY5O1/lUpXhH+2m7ZLu3lsNeyAKqSaKuxc
xL71Q+pB42VQULTrRjEPh0EB8X/mD6uRRsvYIEk3x4hFTBjnO2BmTfLK8MUWhWdEfl362rLyIaWJ
CA9DG4QHdP9sj/Nior32pEtxYpXzOhYm3eDwkkeY6yLpKjEs0VPWQiJwJTo6xuQfLv/9J1Eh3nnk
vlGE137yE/Kz1Eo1T7LzKlbtyVAdbMDcW2DJYGu19R8VQQPdeIfArBHCxm2WGxXua7F+pYiZxTcz
4K4oADefEg8Sxs9UD8BENLOE+L6t3di6HXq/TMP3pfW6QNwTiHqEWMcXd8UnP+WO3i8L4uSHYU98
ZS7JDl74k9MLMeufMEzgAMP15hWRWB7uSsvpzTfXERgBp+BsH2WCoETXvdq5QPHC/JWC5n2mTUv0
QnjKxicMr4LwdAsUqp1idU0qzuNTQ0ye/D+9de0fxy4D6S09m/xE8UNaBXAhYCK9RPgQS8f9MX5v
WVTSG1OLfpU2QwZOgHCRPg+kC55+rjMJcp2ZourR94J4cJL4HKkQmIsrIObEaUWCUNSSz5m+Aeca
jpWaSJsE2SXIDmmu4G0LdjsgPgigQOdXdY6PIdsHFCSN67rEFma9QrH0SzpszeUc8Eg15vQDJRuc
z1IdLTTdz7BCGWEHLBT8dORXSOLUGt9cb/Qw0umAsVW0T09OYmS6bR/doU/mi07IGRzcGdernoJa
fnNyIbP/QOeZrgsj0ztwr0wfQZP7YzoM4zicd3FLrpJcHoVEEnV7X3Su8qx+ixmP5fFYNYDRbYRq
QxNSSqFly7OtKEKbOsFQnAeRTCqK78qNReGO2lUir+3DD7IPkHrNxp7VXRuXkVOw4DVqfutVT2HZ
BwJfknBYNUSroaUULmYkpO/t01Hpmuz0F6VRWwxvLdXhohfW2KgXcatqgsHIn/AK8n14jotqtdaX
3JAqrbIYh7mmhFE0IZh9tT4IpksimwZ5oZn69evc1FG92Nyxbj2GRfavGLwscpYydjFvqH7jSLkp
qxL+zxiVE5/KulhhC6RkuXnMlzq6HJAmMaUtwdw4676zug0ETebt7abnUfgSZUddajS6o2nkCzAL
BEjHi/niKoYnSfit/Om1MDeSMiJL8nk8F9LCocnWgdnzzJpUmR1HYlsLHKavbC3lWnY83P5SoTNs
QsKq8kCSCvQ550HibQ9aBSB4/o4Cd2KFrg1tf3m+Lm97Phh16zP/t0RKlctP6wQA8W2Ba98rlcE0
bjPcpiTprmw3P8rpI55hy8/hrbgoR/5d8a9TZLvDn3XcNcsezH2schZjMRYpx+MKu+pZUyrQEy4X
fbGKx6Y8nC7yMOeI+xCO2Au4RIcs3ohf5s2J/Q/I+XYEpm/l3T1ZW3rXgq06T1yXAA0o7Vl9P8RE
hyEpWLfMMIjlPr3041foQsrVWE8TFjXFk32yWFkg2kV3KnHEPDkYFZJWuyNB4/d6qgZkYeQL5L5R
b+goMahWRYaZAmme0agsreMwbaeoKZev/wzX3bSVknv7Iy33OC5cmxYTq1HiI/GnXivQ51vzfy33
EMyu4np6QmF30rE2lY+1TEFAjmlRFRMGV/0gEfBxpY7W4GZIDKRwmlUwvVcfYMnEpnOi8YeGkb12
76Wt5oHWFG6Rz3fU1mdJTAfa7fNVCRMMhytttzATfBSIDkFy2dxDwE4J7Skmuy2YcKAjgxIPqoUV
zT2uox0wfC5OnSLx25Mg6Q5v+QnxyI48eFw50TrW8uaoZAi8gL0HphFhedv2Ww7JzkuaYw0DX0Gk
EA03Ia+IFSOerleaU03+AQOj0uAUYUZWfhO+YwVr6LShlaU6k+TZ7CW8SMANczo04+UyORMiPe0a
5fPi9p085l65hKmhOePpWZxudTLzDTsnWt9bT7/iHuoxf3w4DAUQyY3utp39d3FUzGfUTTSYrsmh
Fj01YemWFfhfHK8JsvbF2QBQ9IW4QzFdpZmvLutDRC+L6j3EWz3OjMgePcaRRn3lqWNDQKuAt5RK
MQynq7DlVMl+4KRkG49Pj3mvMaHf7AUFX9G2gwbn4NXQ3Woji/FePK4SBKBa3+Ek8dECeeif9Dci
T8fhBElQJ+4BiEsZqVrDL0/hGNrF8dMFa94ViE9ODPchxC41xScqMc9hEYJsesPgjNvn6Y+rMdmv
/W33tlqGAqmfS2TtE0r6VaCZOBZqgaccTYz3VBYCesPuwEzGQp5pdO2RFS0xBUoz656DQCkoe/pG
zTo0+cLAJ4KpyE9Q2k6ZvUheWyfgkJStRa3OW0X7RG8Tjq9wKRSlERsD30i8IdZ6t5QuQ0NoZkXa
bkxoHmvM5ThQbDuxSW+K9fNKJQKYKGvmLLHYTBQWJcCPEU1Tz/lVQBvoK1sAAqCr3lHfMnvrINGv
bxQz3nmkWi/M0Z4Ko8nAbiQ5lH79Qpd5+7kF+3MdDMX41IOmWUozC112TlmXdGn1toriFgltLSNe
uV08wzdyQQhgPxqZFujAsn88onW+kFNDCxdaFtTxtTObUu/nv0alvtBPbhchXKcqYTRUgf8JFsy8
Aah9HpcsdIruwoKZmoVGCsIlBDyE77Z32r0W0iCsfu220sDqntWm6sBb9R8l+kjalEYpj9iCc/4L
clKrEqUkJ/wAgD9JoNhIiPqI2S2cdevjn/kFk90OSFWSrS/R3GK7uahreVtDgtFgKpOcqBIGx07h
oq7E5DQwo9bEHpdz701GkT4u/er+h9w2VabldUZ9owlSiaP0yXd0SQorvCzob7Vmh/OcnFEL3hoW
NoY2CDjO2MJ+fkq/EbagfQuA8OwKN+890oaK3GvQbcAOX37SKcp20WZoZ98SC8c4S1vEUtOpx9/8
2xLzRR7Gn4VjfqHMrubScOd7HMf97b0vSvx3OqVVXSfQhzAaP9VEzgON5xlKK7HnLcaJ4TUpAaRH
Yrso70jApQ6dRuhsW20SSbSfDI0Wvdf7TGCMAqg+q4FNtR4K08yS+x4nBuZV5QONNYGqfeCUSeLR
5HhftqUcU7OSiyUZ6YzY383ME0Sq/WvzipJq+2571u3X/vf/RolD8wQ7T7v4wV5Eq2nEeLtYjEQu
II7HDb22qYEIOjUuhxtSlJ/X6Umyu0mHvx/ae3vZni/SRlP1ZZZZZmM9fewUxA1NaHI8UGM1iSwY
Iimg+WDz0/ahl7uBOozIpRWOv4OixuHzH7+Jv7hSDLULZr15+0wEdSfxckTtVxoZ+Xbq5YIPiRec
3GlOxNyY1YvqOSUuqEvYxNFLqtWFwrHX+9sO1R0KDofIXfgfdMVsj2rQD0XcjB3IwUpkzMu9qNpO
xLgTlJBFbVuCn0/6ofcv0d/6rr5eHD6qsef/68+zOpCrGMvBeGr5jJjQGPi0Ij6Gmcgpg3IIPldj
yYwoLKD24jNtFb8vMu6qXGrJccCWtCyCoZHv+4xKvd5d4pRo4ankHrIGlGE7UtIc4AmaXkwWOTWL
axTtix2oMktk1tU41C4CCYJdOKqqU9YjVaGZUXSlG5f07VxDQLwaKp0dpe3eAGIJuHXpNuCbi6dU
/EpukOrJIGi28HIWHpL+7R13TmtzAuAR8SOQfJ+JAixuUFC0b6DO51YMyWpOI+tt9S/W/aKCR8Tq
11bvJAQtnSIPaKHBjZ/8n+Qrx6WJpLhhcT52s7wul70JFxqq0FD9Z5pHuHO2E+wB0UnmMzkjE/Nh
XPvVdVGpWxY9+doK6Ly/hTMIKB17BAyCKi3qesqU/dttTxgNRMjOYyYf6dgLfm8uaJeUAmHVSJge
niogS5G6gxJoHZ+o4l3/oVcr745ACmwJwRk8jmOD4jvFu8C0L3UgeknVEcWKU5GslzmD/+cjNE4j
6cpinRKDjozg8thmUbSn+hUXvmRJTk/CrikcesOtYsHJNPhpYeVDEcNOBPowj2DieTD4V7rrCHEp
F8OFv3JgfYgNASAMBSTCPpEP8bLchp3hYZyI6myf5IElBX1vwq7vQbbKEgc8uM+ukR2zPHC/MbKO
2WB2XMZ1KKaH3/Ybrs0YOLKNHFex3PtI1e67JjSzPP/3BUF/sY1wNK4m67VyQAxIqftkv1g+o7HW
6eS8Pc0K9KwyXQL8tj/8JduVq0VRKDeIDSGQskwNYNkEV5pJ1d1DVLUJzZNHfsi83QCG18iUw52l
qTfgjhTcovFXZAnIJtc1+gVxPvfQGJdN1DEBLnDh4CA2ZXHGbiEyTv/WBk1cn7f29oT3Fp2d16Yx
MEWYSG0RM5aI1v9Ys596jaX1H531+QktS2wDIMXpEz0L32Annvjptoou8EYPaxNVG7083tGqtbpo
WkfzF1FeA/U4e2138StbQVwLgRYpmqeouVIO4GFzHxuH+vY9lWN99G/xGCclp8d6Uv07ObvjWmYr
OCf57QmR1D1rxzuN5X3Ihc4tCpcbF6UK1xTW+ysZSSOdHBQppUizvGgFchPpznousAJKiIQlgzCs
TLzd2FXsPYSOEPLxCD0JsQ7sVQwGv+i9IJSz/1+vcdJk3v74E07P03vzLCbjcMu1GonWxEjDpdNg
wxXobYM4t5zUmy1j4wyHOrTC/P838mHTMQ4f+kmf4bS3hWN/bdZdNt7P/2gCEJedJ8iqxy93ZXKI
wqxV+nC42RZ0kcJGo+GVpWwP1FFTOaom+haxqNcWNNACOUxIsNHfTIqqI4Pt0EN2P5MQtfHSuGfr
KXrDnVa06rf2q2EgZ6RX9Z2l4Y3MKL8vcU8e0bAfM76xXNzLOH5MLKvZtqTUoWk4kvlRycPYHU8O
B+865cylqatrKfcDmODLObr/P6NGuEB2mauDMlziWquID9gmeMExeopNlpQNPqGtXsbZQwlocII1
Pb2lUIUOpDa141YuLJ9RUZPynBx0q4SsGN+dOeJ6evSzmzAi4T81K5TizvKa0d5IzMg3kZMsek6t
4uHonENJTMvyC7yQoi7yh8pgJ+uu2iyZDL5+kUGYAE4RO8CG7Goy/5fhL6wPNBEP14g9ASbrbDYm
spVwBqh9/WTfXqgM89TkQshda6b0yheHl9OMiJT8Rxmo3l0O8+mwwI/2FkdHG77ucKkLO0+sWqjd
rTFdIaOBTubwwGcUxuxcaGHMjyYtzEXZj5qQPWGECyP6zBpY6jjnM2dwiQKamLVjUCZqnIIcPv0w
EVlf1h7SFnc+Co4ptI1i1I/9rBFpcCoQVPF0/VhIePZ9d1AtCZ8iTH6Tt3wJnRaBL0XiHRcp0GUk
Xqugv8DN8iuMkUz/zeSKKEZtNm1fc8o48qva8YAPQ53NBeWWj4fBWlMuLSF05jNKT/jkks4JWWC+
27rQBsCa3JHtrjmN6t6u3jvQcLtQbFcrHj5XsjB5WM2MkJZHs5pwjFt/znSU9wN8oBSlO6cxAgTi
jpBB1/uUqbC1ACYSS4WXdAUzTxmMdtgEGKtKYv8kvd9lrgv8whVPvE72C3KJ9rNBmBrLGLK4MwaM
LtVJdULHo0zG+8m84GB+q/sEGAluG3Jy3YCUz8hspJWwN1Pja2TxM2OXjVGIfItRv2gKHRTSOn4Y
k2pYzvwerEi+OA/Xa/ZJJ1idzi9M+asH7XFr1lyfYyC8Yc0jle5GHlzIJmjroU+fqwPpBKfvpXvN
JGOSKKFU5RCibk7XB675DEVEjgCmBVCV4x/VGVmUvhjkXE/tExgU4HOEE9qaLhEMO/vbYwiPkhiT
lTXW8hhS1C4XPO0d1XaWPb7SnWdpr7zOlq1w9rSlEh9DQ3d3T/BAemp31dqgctPlbJVoZvd0K3b2
5HgW9EZDmcyG5Gv6rgsE14sSz7IrZaOIeeHaw6cPDnZF4yZyXo8W70W6fvlKarrGfxaWtyAKOwcQ
pKsO49ikd+oAYZE0UotlF4yb0vvV23aii8UGHShTlQUTZHMEsSe55En22s4F18JlfWr1eS5+jdX4
+hvmIwzly+2DfbI52OgpaODrzug386Ll86JLSaBailsr4RBjaBrXFDNhWDeUBtb7/qNrRiBtgPWo
OSYcY0uAjcr8J4Wy6BvQsP2NlNUVSMgIAPksB7Vgm3FXlT/ZOYKVbFaUAV5C7VEmsX6TyruxPaEp
xbcljwaI0O5zEtrafYMdqSwBAqif2gvW4L4V3dalNYHpF/ATLjkFRfWQmb0eNairORXC8feYNN2O
h3SX/PZC8iqv+vpFtYH2PGvq8UTdDVZJlJE4UKk5ymG2dofI/gWD2AteO5fSAw/gCwhi++WbG+oQ
7v6aW/gwyOlsNEDyCTNj04m0sYd7vYYBfv3frQaAIvc3dVMOIFH4AYykYNZNC/7/4aoT2mFViwKK
LhfFHpNnlJIQ5al3mx/UmFkth0FTAUWt3k8pygZGyOx7WtR/0PpwzQJN6dlvwzeWPsCL+2lF9Emm
VVubRQgs/xt2hP2UkJrGr0E7lZj0y+eucWGArHbwhHtYUzxfUsGHJy+mb6TlV6kcrFBjqxkrb+EP
skNcWttV95mIRwGe/8ReuV5c1bFzAlircp4W6z1W+EgfGJ95peFG9rDKW0597mDP9q6YvZhtw2N7
s2K0mw+UHYxpbn5epQ+R9gnoBLAQMIerGWQgFnvIXkizYIrykKAQBNrubJu7euPEBwjI0xQkXfCO
k0g0D9Enu/X2rnWsjxNUovndPR39u+42HIX/f31k0PJpPXBwE9toOnHg2RormuDtmRsjest+ltDs
hDhS1CnujKZgnXzk4Wm7LguZOVBm5bPCYAZeckLQ3o18iEjocdkkKFC/HhJSJYsb9FWIzsXzNSv0
9bSCXcYSNzsWbSxUMRhJkWMmTrBj0qDjZT9AnnCLbENhq/Wge6hxeS6sUVHDnBsOrv70luDQOCFI
TeGmPH3LXk1JVZvhLqjYunxHXmF7CapNPb1inq1ehYYWQtYgFy/qRxLTKCX+QJXZpnWYFFQ3mhXu
j02RJaEopEuKzpcJMY8luPc4Oenm02A7ojC9BTddgHyYNITfshdHKLbsnvYxXmlKiLh8yL5GmyL1
F/4kR5JlOcY8lExI2KxEzikrU8t1bCunP2GLXechdBDrFMqAbeuM6u2xBhaYewUVN4GWo6TxGHJB
eN903F/ufGDHTxwBIZ813r180uShsdEDZEEpAs2FFnc4YipHqrAgpsp720lXaQJAhzi+vfyc6IAI
702XQSKWnSMlfFtoGp2maPKOadVRYA0L/vR8tzztxCITpTMFVG8eTfSAAWQCKkapyuyjVPa7bNYl
7E1Krcw9DOzqYMaBaOFnbCWprNBExKXxDF4D7erakqNvZa2L4wFjt0hXGupsEx5y8zaGofruCfdW
UyJ777HTEURYCVngIvrwjJ3ApEtNICUQxfMFPUyLHXgyVFG7pUF1/kZBs9TpFCAUZ3Cfirp0IZ6d
x8MNJ2EpH0o/Hi85OjRB6ttfd6Oix+t7z0ALZOePNldE/GIXNNpJIsjYjy6BXi37LfWaDLWLLsxa
VPjUr+Mc7iPSXJ9UGExZZdPEsKTYrv25GJbHkzeKGBUNe7DrtnoRAdhQNN5HuAQ4QyOkRiRT97or
h8GIpVRupaF4UfvNKKVMVTnk4nGPndeTjOzFWpkNS9b6ovqpCHvaIvsRUsmOx41q+p2NSKYzTxYo
UzCCA2A5MZji9BpGoLZ0dBA3GaOqnqZ5s9ktU8agxA/i7eNVpfztnSiHXlrmXuMDVJjBhO6KxLxq
npEpBQ/qq+OiAcn8JrdcQTmaUEQt9PHybYavdqzOUDZX+RqZT985tuRfvwDXpb60EwALhHBOkjMi
yXDrDDomBXvE4Tf3a/VrcIG18PPBUCk7899L0dDicabGw+zNIKNtlKzcjUnk3RVvckUeJOcXGylz
VUSOsuaVXH4QqVWrVehtY62uYspG20avDCXOBAEIFIvKznyJ2HsuCYQUzDrktj/MkeKwr/7oOYix
8bMgFO9OCJ+Il5XzBrcgPWubPVR9RoAVcsBl/OE5uymNHqwt8GDI0RIBPbwPVo328svpwOrcb5GQ
WXpiiVeHI/u/+hjNQJqbtZykIqAV7hm+2CM8JQv7zw57TnhszRk0totBzma7zzV02ZFahc/+COew
MA+0hX5Y/2HFOsQvjpRNZr/ZrMFigdqQKFbyjSw9MkFHaZD1VIznnLQmgAf6FpkIM8SzsSh+ZhGQ
GFo23L16Xv+gdlYgOQw8M7VdP76A8FWrLnTtjn2DSkEYOMfF/DW2u6j9quICt/UI08cxa9cX0J86
vwSc1LBlr5Dazst0pT+1c4DxoGdItw2IWapqNhQ80pyZBuUZIFdb0gGj/nVk3AtzrW+cSAm8fGsv
5R9IlrWcUHrbm8UN+7baCOKYoxTlzWzwavKmU3TfWc1RdSzONkXEdakZnAw2dj9/ZoF59K+H/HWu
SGbveSlKDXho8cWWe+GzCFgdj9Ct75I0ttVRTLCF/k1rOiNGKicD7D73WIncunKgI3YBeCzvUMJ7
iyTrtZLUuDVzEGqYb329TJA5L0uQPAWP8+HfPwBK9CzLLrG2JF15amQ0dxwdUwXFOBd6DP6ukycG
ziTTVQEox7rxBF1M1ldeWKRuhqNn6G7jykvpkQxOXz68r2kNNBEgjKZrdBI1suCxkcfTgS97FfgW
1HRYMeuJRLzLhVH2QJiiU3UwDPz6+Za/Gm01tpl+G8mdTUuWp59on4FXi1BiVjxHxWii4nX6++8t
7n/o+Fc2MS2sXOaTWziVmgJLBYumkvED0EUozqIWRtkTBd1qMjdSPLOVwZWB3Yyupz3jL9mhgbN0
wY1TCvn1yYL3lSJ/ZfaVn/sRbhqy6DXNYtGhfinmRjwebNwaeuYZSg1bl+vfijzAgXf/VVoDiQlc
A6HkjVoTJxfXDV7DZ6XUAEZAykjSLRE2kkc3p7shnQ/u2a4hwS2gXyYJnELJMfOD702h3hHRrzW3
kjJHiYwRf/Z941XW8qOYqDwi631N8s7i9aNJzCrpVudzlM/1ifjinP0odkfQPJ2Z31g5MJIfLBdi
Um1IA9luMDv5gvrDhqPhl/oISqCJEygL8L1g+AOFlByQiuq5NkvrK4NzK9LYvfQwFegC8vEJEVCS
7RVM2b41/N2IeUuuolggL65rq88r2vCbr7kW1oxNBCDDFUY2znZE6PuhbQFxE6ZoLNwX/pANMYZC
iY1qTntRbKY4Lna9RHBS2I4QsL0Zg4QaA44ih7fTgtruePg091OSZuNbV8WHYRwTm4MTcx/gFSAq
I8/0EZpE/mHr2UhfKtll5W0wefQM9Bm7l+VGgCECSeEGqOzth1ocgnc4y73jHdfaKFMez9aP1dUc
ZvRI2T3+yitRQBZParWo7P8ye5ph5L11naGjltN+gYUwW5PeP4Cx3czZkamtD+Hvjy/u+ZJtet8V
ln0WurHMSvZlXUkJmBc0Irtw+1CWuc02iR8A2UQ+GTuzHjo1BtwzwT/lVr4p36qsPsN+8Sdm+zRu
6DHC1K8f9W5uW04z2N10VhwX0lQrITdhIm4UvIOSXYIwyblMwQ8W16C35/uqdBlnf3PueakGzswD
qtnCLm9ithHpXWmzPbiaHLSJiv5C3AwWJ5I0WQYmb0J1uk9i2nKtKMQMgA2zErW7TdGs70sZZoRd
xkHdLkythpYbZU/m8g02WPAkIrq6wXl+wFEraJLw5OPGblWQ6BETANWvJPyzGzKwm/H8A7p1rnyc
sQgXgsY5FApteo3qZfsOKDyAKI/gEtAjFFPCyYyK52Zwsjc/cZSoCOj0g/bbahtAB3/qDucvWH1A
/9V2Gm3b/P2i56f4+/vD/RLBArhQdtbY8Sew+njJNGVB+PQGJhKiCwgW5zelcERSf8UN1KMWCjqp
3r4KAqDZLrpJHb6EL9RfW5WeGmPy8HKEt+GM8RkBHqLMePHlg+3GJzMy6xQVFhPW0K7fX2V5/9tN
Vf1rz+bCOVVWumaHQw0Vi21W2LQ6W2jl+5kBckkJSJRQZfMO/TbkNm5ikkg0eODV2XkNJxvDXDZc
NAtkYee/RjeozYL94Sxs4FBgrfO+aChm5yToakKHdzrtZRJdhA/WsokOymowFyhpvN9OT2y8RZYo
UTmaQ0lRn3fh+ohi1iiPrjosO7XRiTaq+4GXaPOQXlfZ5JNNjTW81aKRbYEvlXWibuTgzYbNxeVf
JVKDY5JRCh+MS8KrUJlvxFFAmczjNWKfNiKbTLPwlPRjiTNSw1WJWPVFunETA+R4a2Lt5cFFFCsW
utbe/bSIvr0AKRQPyEoc7LcXRoqW8+IWKH3iqyF478u8Zu8iLvvNxqglWnirYzBZjJLLAsiwpJXr
XKwca8rOrKoAcWtTBMd+nrszD5L+L7/84gzbLSEJhgrPov09n3EJiYhTu3usRvHH/7DhBmiSqqAz
q+um2YMf6txkZF/4sBIsqKIq2EpEI6qA7VbSGkqmB7c9+GIguaqh6BfeqI/J3TqasU1r/D7hYJth
nhBKzC3uZ+m0GF398eRGSBlHY42y6kNnBzWlTmcD7dpEuZjdNSV6OlcJdIBOul8XytW1N5MNetue
NHxbiHwl5I+OirO/kUfjl0Y0jbC7SoxFcVV7CH7xRSbXLI/0h6ag+01TvEQotLLrT6rwwbmvPlhZ
WP7hmlbtuf84lX4uKCEoxl40G3VMFassXOpT5Zhr54hUgJvrY86t9+dRTxKqhSiOVnxNIoFq5i06
OKZe8WZesfiWlGSXxYhuS/jqbfXtfYqXIcTFO+sPbJBFmFXv/T34iCk2Yugj2fij8o3Ob7MsQray
VSQRDDVhIocCMYz91IGPmXb5VEmLQutu5AMd4iHw2ZkHMzv0mKm8dOtU26rAQkvmNQAvApcltTpJ
vQyF90Za1ucR7lkr3o1WuSLJ9X28qbheTLlmnLYHnpalHAqyGrCoptg9YcAIf1xq9Lv5gLAtGQ1e
4rcGvhSCm7HaLGBOicq+jnvwBPqV3rFbmyOyu/xZIjWwiC7mvjgDVMCHyByT1IzA6BsOT6tQbrJn
PWIz+jVTSskmEJDRieAd9Blwzj0OR3nIQ4qJXzHfuQhsPA5G4nRpQsVN3LKeuh5hHB21h9/HellX
kGq/f7eB0wzAnNZVtXOQztL4qG26hMG3l/N4LYC5WMfs240ybBDoV8gWGvL2EzBsSLHfTim8UbYf
oKousSjaTNq2U5/VilASMPak+rr95J792QQ56/98DSHoYJ7Q31AEUYj6lFv0vhXRcCwFGVat3g3A
4yZGhqXHJFhN9NYGqqSRvRwi9fTZz+UBQvmM5iMeA9MC07RHmC5lG1kfeDZ1PxxXBjRnbvGbdTQw
IJ1i0n5Zs0azOhWMven9ekeYSqgycX5HCu7EYoKcKmQy90aVIom2/juiJZzZphCxdmH2xf00y2Dz
UwLqL6bTjmKXBsoLQZRBCixs0sUCVrycnCQ6xcqmzzsyfq40w18cQHZ4d5jYvVYniDLmZDrtjqHR
99tzyV7BbCBVRPtdDBDZ0EyPdefULXkZM9Kxm8lGAZsuzFWRxoOcfiq1c9IILuZWe5DtAkyW0c+X
Hpe7yje39EpAJCFr3gGN5L7gOLs4Wuy14O/rmKDnong/SUirBqNoDrSEgkETxVgc1FbL7SGzQY2G
2h6/37KaWzFiIDwv8UXCWr7EGs+h1jh7451AJwY2gmK1hQUJ8p70YHr7ErxTQ7LUlo4tryjKCUE2
sz0CL1YfnVtPA9voyeOK7lcxjLm43AWXQz+JLwCO90VXlXvu15cVz4zBHTKd2N312sviCJK2Akjj
fR/SEYSpHmzXR2KjzEIJ/U5BZGgYztw15aT5o6OeDett6gwqal57RiaJbrI5vYhw7S0Njvz6eoWE
HXjdwtxDe+7HF+J4QGtHLqx2RDxkiAVjrg9WoYK/I2ZbCxnlHCGBACH4161t5mDuOVX/9wTiSGni
Y9FYbPdTbXHNOoQbA0zWY+3FML68pYnK2QzGMvkGWagr2kmrQaMa3cq2ta2TpgKPdHlXU14qV0cN
tEfujf94zNx6qdT6e1nIwCefJaWiAwZu0y3Z47OhTMqnjf5OOTn642sEseyJljuY6rp2DUzHJOOV
I6K993JnMg1b1yrVVS4yMHh2w9K2Dph4HhOURkEUOxeiqg2F1QW7XP4lrKDwfOxO1TLUuHpTR0AZ
mqXgZ2jOD1TwanAOOT+n22wXdh50A+jMraD9PuVGGskCTdpRlTufAjJJdqpRTXFHmhkXWgBrcnEn
NrlqV1fExtIQw14THdWf8ij5dGvGuBaX1sMiV4MfOWmeAQz0cC1vH7fivt1jXGGK1AGQtK/XReNC
1jM+5xCNDMMiofQkiIOn+vxBEw5gnFlxIimWEm2RZcZsJP7mnsbjKvb3hcv/Bc6xbjhm3s1kNjXT
gm8P2tcuAQVlx8zktQ6/eXu2WGFim0pLrDMDgO+ljLoVvMzCLAEB3KN/VaM0KINmAZ4DSkbotOx6
bHzj+wNDz+njZ+DdLRsVIZacYfLUw7SBYJbfWPr7+B7btu3XRQWcF0yWipKx+E36gv3EX9pc8XT1
O4t5roO7knnB9iXeTUXquHwOUdWOpYGRCVgJJ0G1ojBjtCYu0m+TF+5uPyrRFTJfr0NQAcsmoFX0
vBOqTUCYNdpqXswTutzIBtC8YoeWDDHCIsHM/5ADctgurGV9wUtbXFkBv6ewpu4GGJHwbHsMEMaj
XS9AMz5IoCPQw/w3mjRh1Q+q/UF4Ep7FkDsxH+Fg9/vJLXj71im1l5l1XEqmRoLraenCZjqEdtlJ
+lxbHD5kslWKLh/d80gJiilnDDTB+mpCntcMiJBpxX+PRSkxnw8i0w9Gmktg0JFYZpaeSAEsi494
azj5JA58t4BgpWddcU7/srL1G5EeoACJII2GplXXlLOLoi0/Yw+S2zEFVmXiJ2kWhw5SUWL9fnbw
pGmtK7Zg+jUncIA+2z66iG7qafAD19Rm3FtS52in2gM5aSVBzRIKkhrq8Tf3AqmV7wwbm2UBMR32
0WGYb7YBlKQC/TS2CUY6pYXgPyIFAF8/44k/llh7glfGFlSWYyOPeYnEhMYY8yxsIfCMBAeig9Lk
cTF4Z69GFeivDz7Xl9csVvFKohsVsB76DnY8SuaTzegj4AJphW7Sqg0bxL75p+ZysIponwwTvvXm
TNz/ugslzbYr3E45I8R4OqRIAP5EclOk4BPcnm0hsILOcsV0yK+sRnSmFXQ8hX6owzXRIWwQJdmt
neuU1jvKYAomeqG2wkm1r7GlTxaWXb3jY9xu55LZCwoHwi8oclmAPL4QvBHQyWtPy2sTSbty4LiC
AhAxlfaTmNzVEh5BzhXMLBl26mHIqbGifDS2lqvneaVsp/TwEFKcdmn+5aGfzkeF9Sij1UUEpEi/
TiXHzSB+gHAhnI7Qv8XI1dpDCaIuyVcXyriRKqthpsE8Teu1pTq2N59negMqaKmfVGn8GQjmV1Sg
m7cRie9KUOMb52zXK+RhFeB6oGPcYO00Ei+jtS32vQVRZIuED1HOVrVo4UX4cw1LLhOF10X3xksg
ySi5/qb0BWoaUM+qUnMaSr9UkYWeWVjZi4vc/4HzD+jfvieALgZHvc5/ppm3Btl1wi7J8nTf7gZL
j5pGLnyf8rldS9fSAqPO2nF5mF6y2Ay6i+REloU3NqjhizZC6qSYT//AymF1tYkhi0wMvYZEUEYh
obC0IzqN2nCsR26LzXAaW4pyvh3tSNieilRzASsfDtz11arsggJTm0WaruCxlA88U+ErSx6OJndN
y2qy3NZ+aHf3xSDfJtEy5Vg9/2mRwg1x7ScID2hYMo1DFP+Hl/l97UzHs2wxPD5NbH/xs2ivo4ij
l2QJ4aIzROaXmpNvzBGM7plO4pEHEzgB4wePCmuo2w1rR7tjYzxgAbrXEH9HdmyPsk+yKf1yX3Ap
ajjH6azczHI0wth27qLAF0AHs2H8mPjZca7hjcsXYjrV0PWk+APhGzaRv5UjH9x863GTJNitJPsz
vexs2kLCbYZ3JAgjwmulvAcGeKnh6THdddJF1+HMLjGRZu8ViN17RbTCRF5Dke9tR2gd/UddiRf8
uwbdY2yvogTfy5OJf8cjZ6YSl36ctkB4kdG95oqIw9edSoD2yuT/UZiAQ8q3l8YAp6CPiCVfCejq
8v1Dv5QUUVQGdiB4dECteRlyHcW8qgTrJKZV3yuXNEkB06DzpqDWgThXT5Idf8qkMXjdOcGufyCd
w/uuVFV5mjCdSBWGK7ia2Tp6yOsRiVuWPt0VV/r1rkvdNnpdqPGO3n9yRjV4LNhhYT+0JCAYuMdi
rCfJKpnv6h3KNHSxPKbbk4X2ZT40nMj6uDLcsy3+bEPvjC+gKZkKexAcYYla2vdTrZrApRuUUCsK
vXy679GlUVlAa7mRNleUztJn5SpyFbzGf4Yha4cSfaNnHR1jkHfgyKPBZeB+upfBCVZf6VDXNPHr
6VsQA204/dBp1b/cnmfkNHF3Cs+faDRnL/lOLjIFzyxKJw1SlkFmdq0STiPzQahi+jtdmwxbE81p
tS0Wf5XmPA60s+h3+gnz7l1g9RlRPVTNQOPHMy7ZZxBalUNx+soY7GqbILMROnHU0ePuvdEZusSf
Zo4GQsub8JZrlMyna1upE7KiV7EC3bGjTlIrbkpC0H4FFMPblbp6pHh2uOy2tV20XbzqX7OEb5Jc
UGxPmpyxvhA/5Yhx8+EzBMMYRvE6q95x+mkKzcaTdkXSzbtSMLANPVzCHchueGlfFhZMg+81uDto
P/8W++c6DMstLLQfYHv5Au692s2KsTRP7h6GKMxWU7mJv2s0KvastXIO1Bl08Cn73EuJkRKtmcCO
pezI3CBgNSJk7kWWusNbR+sUjg2VrqJM7j+eAVTE2c6YEW877UMah5+hUe9CWm18QTo2+p4V7cAV
mfC5eExAKIC0FIzMF2FbzmlPFcBguXu7mQv6v7qzvaCbUfjIZF7k3YonZBWPlgtj3fyv7usg2fwg
zdZNMq15NB7C6LyRZEjRweqYgrV+mKEIQU/uSh1vIGNCV7F0lXnmsml/3sNHzXAFVKh/0i8S437P
grNBLXJaCncgF2Pe3gCNxPUa956G68p7cK6Hoo56asKUTDYtS9Jodve07bGlE0tyzjP7d1BtI8uk
IXH+/kMNHU55u6FlIvfDr131GaASbWO47Y+/2G0V2oZsbr6vqiLF0LDpSw0vbH0TxU0lXLOQMKtl
0E2LQMvNVP/KFXWx3/FgBGU1mmWGwtlalfqKJU9q8llSM9bJGeesDSnvSrUa0rEmlJsxqxT6G+RW
AUY04VTExb8kvpMpui1NqRn1jGIYnPIfbtXI2koekNs8M4wjrUB0+F17nkwVkDYWU20zowrRWReA
Slj1YOqSo//n9pUw6jkaa6FQ1l+pshxJFSglhgUavfaRFG23FRC/MvN2zJrG83SqRyh8pQLiyeaC
nnkHGTOQYF6nZ6Lrw8pG1bJTJqSQr8yQAK/YAyaxmq66ekP4reLTnFwQFnTYu3KGi0YnKGMRDAGj
W52hr8SFkqNz80ga9j4bPwHix2gTHgDVnDBcqP5OloQQCBXQebgmc80X0+3a4tzLRbod5RKnziG5
ie0HQGEqmP4eRDhldPQhnuvogUUF8RQt0fuNnyuvxYKtLx0mTaYvBlN41fgfKBc3MssM5PNiL/At
UXDRygyGaqXMk1wKn9AnTStkd5b0VeYPf+vcL6lsmN5uyjmTNfSlGticcs10wKOQCOE8BkQiRW1q
/SyO9cizze7LLJ9mr9M21N86qZNAMZ3Ii7ykVU5cZTfhkTZlBfshI3Mmg40sU2kB1tFAJIOdibsz
RVtaI4baHOazzJygKlKViPfrLuvQp2VIJ1iKJelO6GU7qk0uLTE13x0rCFflNlZ6WlaaUa0kJtPj
6UBhnbekNARkbhoRbhEe55z5KG6H2NGXP1j7wVPkJ0ESVp2BjLllkoFAPcf6nQm0DCpgyPE9VYQJ
tERaSn1r4gNUmcDLxUkwvPMNOGHjhf23Nb3OO45T2TjrMLdzLdNkJdykCX2XBftVQEwv+5QXrhPv
xJ9voMP3uLXQhX5DZq1etqTWzYHOYDazKrtP5RACPIIYvA3gQkqH1FPAbZXAKJCEzij4lJkJCiyO
cUrmUwtiUUbTBwGKA0W2CsFebwyEJ8O5tG339SFKHw9Gf6Q94UaYRoRZlKjAhCSPcTH0B9QffBaV
zzHdbIPUhZYVM9JpfTvukHiELX1WOGOFqpsJNmczuPWLIPM9zjnBvT8KBFe+CzbIe6ATRO9+Vjw7
R0a0XXKepdfWPJW6FUo/kfUVPuUT3Xq3+VIGpLe4+9qoLqc7hLYr0zS7GHducq4TVchC6EYrHuC+
9dhtGHCvMeO8WOfsHRdUMHCpPZ3lvbyibtHZ+cjkpOuarmaTazTvqEDaJankqL3dEQ7HdGLbEal+
9TdlPvcvnnWhwa3N7xP1rCnjDsORlTD2/V8dKUG7kc3rpHGw9tPFUtFqyCrFGaeAeg4b+1ecDaz8
ATBHV5mV1QAaLs017DCym03aqqaNLbaOPcpGRptn+FdbH4laI6je93FFQUffl9o5XIoUzBdDx+2g
qciLIQhj4Lnx2vbTIX5OQH6TVWHoDiAPURGQREaOZbRXNzHAWJMVlWKPPT1sFcqCVaX0azu5x55c
SPWBLiKeK4nOcqBK2eYS3akNf2zOw6ZHObu435v2ewKtzAR+54bzV4Y++IVPhFvWzJ0JOU3nSTiS
XpKRTpnkH7gy5bUWSEHMBgW6F//jhmQUhh5t4mL0WM8bLvFo05L42pOtMdqoRiKXi5Ahe4MM7A3M
qf1FiiuaMbttvDIdm0gPeoX8iLWM8fvmji4GFdDY/7M1MEtgrQwZZL6XOMmvy54XeqAoOzmHGtnN
Lwe48aVIDpGBNGfdeDKJ+oTuZud2m0Y5DkH09Rnzy1v6ECxomq9txbzhiwCP8lQa9EC3YVVe2fPE
Epgj1YY+6Etg9ByJlvxQ5K20UIIPuClcJq8YDlwtwFsbS06uRgj9cBHbyyI4NW+c6tvxeJ+tKtA9
Udnjt05Pk+8s9dfHENmlkPjCSlOQPz85kFxauQUuY5lOG1IW8GTChjOJykVTN7l0WPQCHqJU1voS
5LHgdYlR7eqCoFOmTjqsziM5LujFWuauJkJH2az5fQ9M1MssFSW94OKlkyEI4Hv7mEDKEkn/Yn9z
bm4Ke3RSC/x2oi3iAmpICiUKHugdY815zApEu6Az5WlMjdCaxgFZMFhMZPw/Dz8i1u1bKpVL5xAM
1ZIW1p8rSeFSnD0OFpL2y+l1qoq78FhpZ+CZcAAIi5zioaUDfB9aBWRqYaljD3HLcZbZoe1AkzS+
gG0JWL5Or37jRE2y+R18E0yAo/r2m5HF5oaaFFdjzXrYcYX097eufsdlPkkWKoLW2JDCD+aS7Zpf
wOf91axnAXVr60qjNYXRaXt3hRdXbKLwRFhHLITiQqeoWja9rdkXMEoO1DuMOwjz83nrcmzaIyqE
dmPKFJGKWrvIDn94GaeQRDXd6r7yeRh6dEE8h/lLEtuGqYVceIlfEl0YD+qbYEaRTnMOS8TDvhEr
dfK1r0WKDhTmXVX5gRFzJCgXsOGl0FshSNxcNeRHklmgHl3M1Tuv9RoNu6u2UYEgTAP95MSn4Tru
+bUhTk+olFT5pz5vioV6iEsllCXtyStjLz2ilEFCiVnTAamskolEQcu5pHH8kR3kAMSMXySkXV1+
1BQsnsyruINeg987FGiE8oSBI/EEH0nzFNXs/R0+jTid/4tv8paR6N/936qsrssKqwGO5g37qLgg
2kPgOa+M17DgVJNtlMV6screHT1rbEpeMDx9vx/ktr190FKBm3vVamZ+fTyR6zk3zAmEDavEifdo
9qNpIDrmXMSFxkkbOAgjCZF87AQoCZhYb4UfCTQ/EhPxz39ihauwkTWQdLAX3fxclTiLU9bqxU9G
ACx+FdKMrCdVOvs/8dLBjtIFduorCPc6RTnz4MIPhAGirHcNNXyEpnqCxhs/dRaufhqndic0UXUW
59XKkkBNhTbXK0CcC8/1OkLLyHYGuNkabdsJDPxh6C95DX6Ni4UX1gHsD+2IV98s3u/jjPTY0KQP
OFsMC3jbvb4Xv69FNYjVzCSRkzCo5XOdVTxS1S4rKZKzzcVmAyQ1GP/hx5s+tHajbic48SAqyeEg
1y1mTalC4T0FarTOHs2A1r61BUTsTOpHXHA0ENleJ6EGO41qOgEldBb5OC1JpL+zYuNhbQ1Xy9fR
FDi5nRjIUZ1fnIjGJU8STt8Teg3VJMnfbuxz6UQujaBpdOEml5Iy3LLPY1keDpJEXVi4V5y6997Z
we6BRgGETf581UFAyCAPsLQzZCLS8xl9OmO2k8+JBWUE0iFiOjT+K3xxFTeokhfb18lmxrPB7ibj
ERYNQcQoKvMoLT19sHJwVb1a96gUVac/15EezG1XjWLxk6J4P/rRFbZeAVdw30EgKeW3oBnG8pW+
KvuzsghQL7jUIfWZuV+QGE8tcVD9DYOnLJdK5929DglPgujz78lQR5Z1z6rw61pxfRd0SK4Q4I3l
2QHzk2ZUT5/gyUqsnk5I6sj8AjBaxbZBHh0DsRxtkGhzlIKH4Nl/0VtaDzzKzrnRyFEhmY6ZwzXa
wpv8s94r8vRXT8k9xzrUHD6wQrRi+C4KQmRuSLk9aH+xI/OKSpFOkINh+Yr7M5jhTwHjdEMOcuSA
g6aKXtOu0SV/fbWLzTEpjttbd4d3RXCZnGZqtjMuKVQGbHsUIqhqu1F+BhufJZH6vm2cb+U0neRw
EpY46MzN+FjRhp8MEPHCYdP30Ht8/JA9Gqom0q3Vbh5vok4eqH99Xhz1ZWU2oebH096ZSefVv5k/
DJCCXWg13LdjOz/uKCFd6S/czB3lb3d/JZt2fUUtXPEEikOboubiioDuWXYhGSN1ccHhootua3ay
Hmj+jRv6XTpx5ezfirXJpyqGzsWnUYXnzkxgVMnyUceB2BhARJK+H3CxCug7tQ5BaNZRkscvQksD
kbUP6127Pl1sW60cvGlIK7R/mclL+qnquY5ieAJ7iUpmqV4MiEPpQw9MvRrzLJWjm+wQywz5EgMU
T7TDF5QrjwXFWDPbnC/oiQAbkN6ISvgbxdhK8RLNQKfg1T2QzaK7YQOvdi37f7xHFT7dWK1xJzHk
5poDe2PLsBk4a+akLLaPQNWW7a+tuOy9vcVoOqWJxVqJbpQiS5oY+3sPnMAsNp7ww4ucQomGzXlt
ipnIaS6bRj58VyRs7vt0nLm5OW38srHULuEmqEO9TAxxo+wPoOy+cBdqQ/GcgjY7OUNkaXi6+Vwj
9vw6fKybk2IS1xlgIef+S631R8QqGr6yFpZwe8RKMmA7E6OQMPwlZjPxl9QXNIWHuhjpo71hsHAv
wWQzgo+WxvhjRgnrG57wlvj8NH6pzQoCWhPGK6nry/nY1m/pj/7O3YlLhTC0+WMmss038Ef7h9cA
5HI0T0WuhzKNvUiQDgrnDwStLjnsHktGUalmTu4APxxJZjjBiZ91/o3i8c8JsZaakUBQADM4UQuS
l5kzKQ5Dh7q+/SvGLVZX2M3z/qUUL5Giw57FLMEWiHe9jF4SV9N+cUnFuI7hamPCHZKT5mPw56We
RPl2II6RPJ9o08yA2D6zEmw5idrK//uBN7eWKIHEKCv5UkWKzAe/4mEcJkp4ISDmSY8M611Po1l7
MeilwhSscg6VATh47o1Pa/zjj15t0gmiE37HeeDm3iHIjVRCIT8qPHpW6GcUeK4ihbxZJlIVFjgk
ZhDSBG8pHCRRPsCgYpurFEcNtN9Xr+yFlRn+WooSBFWAn0p7IuZZVc8PmpHgk7+pz1cwo7Gf0H8/
Hk9kjBOjfwv9zwV/LQ/AC7K1FNy8/vHfzOPLSR6QsNPzCHqIhlRa1Apa8ylEkG4ICk+EjHZm4brV
ROjH7Nvq996I8T6WcjhOffxv12vheUVfCrceu8hXB4FgkznDK/18Jo5cT7f+OZQLCbE+p9xK/4TM
q9eOgG9n4zXjRJUg9GU4TF9ISpRf+IeQrtHxwFQaYttrv7rXlFIs7201rhVnXxn/RyzLnT3B4ohB
TOUF9UPz+Auwju44TsZjcXAyeGA/Sn58WHWTeS9zOZSe/fktMnYmzuVZPF2XE76TNNodQf4C7H8F
eUMNx6u5Zl3k2KdjJlLRsjyf5u/+ap2H8oT0EPzSxOCHw3c9fvaIHHA1ty3PzrvNRuRq7JCwnn3Z
PAOmTcnSyysILNmCroeTFnDwcIZ2JWLUQLdqg47N2odo2V7mipoCZoy5DwqV4F/h0/J491X/8drg
BLXMdyRzymrhgZZEX0c5wc4bwG7VtuK0xq32xpLtMI/B+U86qClcMLGOOSNeuctgjxMzYTeKNmZp
JmvLrfq5F+vlRWHFGgnMntL3BSZok7WN7Bdm9PYCySPLOS8MJtcGMN2eJ4K0TU/Eqe0416i7+Hti
i4Np0tRABoj+KBb+e5Zl1hIn+Ut/58iLWFwI5R3mYMtNowimHquLVnWyiHHjbfYOedwPldCwlLYb
yA4X9yH4v1MOn92/jhZ6sciE6CC00jO98tX+ZPthj495GXArOypWgrLceeKlJsLSouuhwa+g/cKV
kHhYcA9IXyUgxpbnnlvG7kZR3QYo7C1ayyTIXl1MSm91u7MdHBwHDYxaz2EGfhqxLA+orcyoeY2K
QUn7AUOdGTtEcXxDgOlxD/lFm0YxqPuFxWI9jC5FwvEa6U48fumQs/36kokJsj0eXTzFdPGK7OKl
3uaL2n1FgWTk/y1TqU17nsvGeKpaNHntnc9e8F5MHL4+igm30UJHVyfrobkYPRbnYyAVXbnTaIct
ZNI6kZHpyL34M5KcXHabNGGSDoLVciXozbiYyW6kJXhPCFbS3IRSOk+UXAf5BOLkq0cnpNF2z467
b7zBraSnkMkmvzY/GGSrWSc+7LcHpl2ziGNWpmnJsfu5oLNDmU+z648RkD6H3AEkrxv36qS4ajfJ
KSOBfTfSg2pqzJa5FSgae1h220VZjiNhYBTN5ngUABYRCiLitlPP7iAsFUTqzpY+7G+3iWBHkFKq
VYBz0yeNDEel0WPFcv+INRhPSV2VeYXElA/VONj6VOvLmLEomyf56fEdWtiiG5tyQaOeFhHZdIiL
L8Aja15lmUxJQrXV+oGIqD4b/mD7Er/YJZtjy5vd88EyEMdoYSV68hkb10kjBFpF8R9nK0oXhmxU
plrIgwE9YrRrFBL8EuvoGhXHLcse/JycBePd4/qoK6+ber66sYiTvHgENiiZPL15xeLO+lMtvQFO
xsaty5FYLdM1VVBOLk09+JfyVoCWZ2XTkGNh6uCiUZU+RudDJ7WS1WqzCSjTbGrw/nkCYIwpQTtA
6ykmKcZmjX6GUBtvyDGTy7HWPdcWa/2OgECy7lpwkmG56G/IU9zU0Jk3Q4hG6TW0qXeak3/Lb4Nr
4TOQ69grCsYpquRTl2P4Dv6U0c5IHBrBdJRBPkL6Z/8CLCV5aKrfiLBEIKCnrmFe04hZqt7HFSqq
EXszW8Y3OfHsGnfb7rUhNA4Prl4uUbkQMYGe3lTE9HdIZEd2qAdnsR2AvP2JxLXxNQjDuyWs84k9
UPc/TqWZciSDPYBEe7G/hL1Fk7YpNitmjcHV9V+IQjPgPdTsLRx5o+zmwSiHbB/71z6vpht18zfq
QQlz2B2sXOIeXRLz9QjLYj/pGbJPoOdppHZ1IT5lts0+j2a/RXM/Fp5ulcrF2n4lXxYhgDBnbhqB
GopYnJnF0OhY31xU+wr2lT5lZdUaJPp4m/GfqOiLvjBJkRPSv5W/bqtOPXT8uZ4s63AxDhRc0sA1
Qc7x0V6kaYJH/M1N1r/tBHVKvW5mZY5aF+TVzggTCwPwfWU+NNLhm6PBcD+fQ7TUsKtBzqhhGi4k
k6VFncB2LgBvsjuCCbp4EY3LPam8+jeC7+S6uS7FeOkUnJD5zY05oq01h67sPPuNSmlPRuKootO1
jpn5GJ3y8ZyoNrHdQlo+aQA+7SRFcJQL0/x9Y05uue/pyCgyKwxqQIF1+XIDZTGkIMkjGaJX/vRb
ikn5yYmxtxh/45iIfKYq2kEnptpWozM3a2fw25jwp4aRRpEqJLVOPlFjggTsqlZ4G3gzy4hFDno+
Bn9q8lD2OaffftQNOdiv2TuhlBBpYJ7nllpNYdd4zZYiB0lKNIMRhdz5haR7PytyWCjwcPTJZwRj
VQ7p/JWYL0bT4TZ10bL6dgIy3ymWvzTGax3UsP/LavZruUBvH3ETcXvhBqTb+65N4MTIcq8PeiZy
BSlnG1f6nkWGs/k6eoyd+i0WELPxQOP7FguopXLtbNEFycdw5ig2Q4jx1yjaoBLLhQ+ajsNg27rg
6sa1Dfvyaws8WhDgOVlVsbkIKKo4ij02Up6dp3a2Nf9LCigEEfXYy2ptkUR0IgmAfwJlK4S4N2R1
LT3jzj1nOzrP18IFEpRXJUZEmrIyXr8lao8PBlp3E1K+ewiomIvVTTYop3/Mh+ihJ5XkWy6BHfFC
DvSJ4cdBv+Su9mvoEXz9uiuqoJjc/pDmSZpRieCgPD82O5Bh4Slxno1i+olple5pUOgCpN6KUW1g
+/s7YoxORw3ZXcVb/Th9Ilw+AYNaoBN0vhQsIsY0AC+9S7RGG8o2LBYPg/1IXwv7vFOPfRd+6pbp
yOP3MWQxZF4cE/H1v/NXswhb0kCevlYeqVbBZq/9Xa794OXAyzn3f+1PGqjczuolCr5xNcHRDbb6
E/bURKv0zRZnqm4/ElBviG/87kYD4NkzJb/PinPmwcmoiiMyvLYZ1kbD6w48QQEgWmsAvFqYn7uz
L/p/fION48nAHBlVw2vsSm8w8pZZCkuKtdvKuIak3ig+BZq1my+jbPur0RMywvW06uQhQm7ziN2h
UQSj9LIUVupVg9AHYAB2GClMmYyAppzu16T79wLVsZ29VzDhVZeAm0UpQmvpWxkPP6H09eFdtyy+
vrcQo7acE1eqyHrFj0f/lqE8k1CXt6bXUiPFP9nzr0lKyNQwtmgDaHF7dka5htlBSq7PMMbdYS2c
rPdtPtMoLIxf8bGoCUx9NwdEdsALIZr2NGPeFnwv5rP2Wj2eWrF0JKLSZnx+RSfMvZDcKK5ZXg1g
NzkhJmxHs5PQaC7hzYCRnw2HnK6uRCaOh1dqtfNsGY8R+XBQQomtBJA8YBvXkCE102DPjhslxiXG
DU7XYzhUIfpdQv/KWjqP00EA7VKweBHbn7Hrq7uOxYv2BDepnJxc5+XkDzvHCebqWnB/LrrvJ9XB
tI4xv/bmI3Epfu55B8Vsn0JrtcQ/PSF3ZoWqp7TbEv/2wV2P7g2T8SDRK8o+qbLJytRmSEiU6qy9
9gg4aE1cWYgnzInbHds7b12mkmjpfOEjwYypnEe5j54KL6lqm8l2B4wS5OVHBMA0KRTHORz5dACD
TqKXhxDac69QI/k9ELBw9C/97c+U8gYbVvXdfhY7z8HweFRbLLouo4TYd5xNUnqkaF0Au0WJocEN
uwzuIO8PP5LM4yS7PoXY3vOZBvkEUBUhHCwgG6s4TfN94u4Il6aEpTVig7ijPdSnOjWLUYOKL1sP
oaiJlcPO7RtROsyzS4Gf4wBfvPYEn35BgSO6qVYSbMfk7PN7gI4mqcLCem0tKLMBOSapsIm+grb5
2R+QgZmLwm3ZJfaJV1hww1S7hDlk1KLqkdNsgz7Sy/Ai4BNwJ1XTqJvlxRqr1aCnJ++WIrB+S7aq
yGkC4Ts2kOD/CWu9dLHntBH8n9mHuvxHKZNJbsxjr5J7/s6cX5bKBDd57Qnqr8di5C8FotTijSN2
5e0yK4nawHBF1qP2r7VPlKYU0lh1rlNZ7GnURhO06bpAkXsc0vCqXZUhmRqfEDbcd7Hsk5ZaeSKq
EHPqIh5z+I3HxwqOFbtGUN3KRz4W50TB/PUy+hcx/Koa4EJQt0aPpLupD+9DtMlT9pLH3UjtAaNw
Hv7h2m/0amBCYBBAKt0MPPeY/S9tQvsijDOJPadGq9wOx/ZAecRoI0W5LiVcX9lgcQpZRSdMYUHj
zFlyfV0GIH91E5Rax/7g95+xpWrHMDjhTs0pHXu6S/SsFnBUM2gUZQht+1Ea6NcCoNI62/Y8KzEm
brpuSmLuMh/qluYFik40TspowFpwqyM5j7I8dftqhVP6gxVKdGn9D6eQa4e6+Dh3I3BTfnUm72es
+LLaXp6dSMPZfaclsDme/3mCeE+mGmoBoliH6hSJEE/EyPULkiI0gGfnl1ky5M9q5P05WkWaeokw
yvpVDaYEatj26IBdYSxkqymwu4wKaO5u/UPSZb1i3d+065GpPACZUPPqUo4nZ3nfEiNgk8WsAB5Y
PR0EGHOpaf9A18t/K7r+RAZyVlhSrUnohzP5dufaPfL6ABreGNepSM3MYzkOt+ap1kY/0E8VbaRT
e8HkxjSGV0W/8AMAFi1EP/xXyLvQhDmzEwOcp7vMDYoBU0vq0u26s4z8/TVg7aNhMS6Bw3fvrJK2
cjZGQ34kuq+sfcsojkDvVI+m1eC15seObdc8Oc2FIktPdvtH6U/iCTUm2L4/xbnT0Zgk1UDj84o9
UVVTPJvSdu2NYmh/GSkxfjVq7FSkDisoo/ZnKkBnczRbS+z1317O0sEqE04afB1GA/PtqHkKcJaR
KY4BCbFg1bpfnEeiGBVMr9rUTWFGLkwazJWtl6WkVAg1uhiL99nM0hRc2e4w6+2ETz/r5gsX5iqM
0Zxrdo0fRaECow9Bn4NXPQHt0bdCERCrQH6u6UdZoBfK7LN5Ntq1DrSGkm5LsZM7v+kyC+TMpHef
Z32pisiERAZtsQIM/QefiQkNHXq4Bgp0jCKOsyrnpbmpFlDxEf/oDWa4X8vxB5Ybi5cFH2L0qg4j
+ZGYjZeRkMZwuLNjN6Up0RzI7d47fMyRyh2n7SRQ4a1oH4Mhup21dF4kZBN1u6XBchKrGRgGml7E
opItNaNHIP7jfTmN8bQ3Z9cbT2kpPlYihN6uK900tQFPhmkHVSr1p7yiTjgxIxKtmMfWndz8Jl7O
G5W4ea1IZW8SBczLwm/CKJAq4SQdq/PWqQImY4RO3Feg13PHm8kUy1Dcp/i3uWsFjmruc2j0kDg8
cRvqWj6GN3RwzwBM5hQ0upq5OnDG4NvD07CnUD7NpyZqicfdFar7Pu5vONFt/YD3Vr4p6WaoK7Y1
aTYTRRE+pcTBwDfIrBOFODbChRxKmVJpN6qPXg4bqttjkI2m3t9dPY1F8BUXE6qxpHG8EZf/aBod
g8AtLMAhEmui2Ys3RGzjd1KfTe5EJSu+jC7c6pt7sfqbze2nJhgLJ9j2Z8RYa+r8dJywujyVaKTx
/bRGN54DioO57NaO6T/SR/klbqKhEViLMvnG1jMMWb256w1EyX2A4KzSR+mOYZXZOh3FDqlQgzmf
3ElBhEEqIIwqv2Uy/eXEEfidmnCk6ygNv2HbLxZlFuJm8IQU3TCh9FFi22AKS8UKOSKH8QdX8Iuh
6sS2JpFgKHbztOU2cV20qsN6eRYZ1gWuVjQWp4r8lMU9oNovzBhQPP/zUzgiuaMrsnU0SrTxPfvU
x9iZ8iYfUb4zV23cXrUlD0CGTUp31AV8CxiHVSMpbru3P8w2wYj1AxDzWER/pffQjS1l4o7RKna5
adBBYHeSG5VdymMAZJS01DISXK9qQa2/qIrpvjihFmJ+6PU/TfzwnGZvPb1v0GwGi9jlN4FwdtnQ
ug5mCdkJcIv3gUg2HnOcLwcOXpToJH3fbcYuEhfABMAVlACU7EVQ4yEaqrTDjgPOIXGIwclbaJIb
UMmw3I4sTVJiPvpvwuM6os4vMDvC7T8S8F2TXlqfYZ3+yVdVziUQ88TPhCmyhL0ZBk5MFg2GyZId
rsKJyO3RxFuFbi+7G91NF4ivpQPCLXZK6mXf73CO2T6xgHJifyLnq9zSDxDM7tiKmS6o8y47qUZZ
oMr2WtO53U0dDJCjIy+tzxJOyq/gxB16JMJ7Tg2p/+q0kwmUxJvmYQrFXZ7PDAXTsfka21wV0PGe
wmcRxALlu/Q1vicxmhfOa7sVHmZak/8lryxGcaJmVxf8lQW5cam8gHmcMg+mKpxKuGu7owSf5BKi
OO5awj5Y9ENgHInbrho+ufI6SeLYhVGUIicpKLZMcaPetTG8qyudskXSHzRM1NFMBDifoYp6KNc8
hGrgc7wMSszdCQHEZbBCC3d6vFWuOMtBlWy6+5Xh++s/XfU456BETgDP37F/CLVrH8OtJ/Sa4xtk
vcYrljIWy+6ixgbx5zeX2+clwXwZNnLmIkBZJP7ZkWk4qEby22oa5EYu4Pgy9HW/+N3f4rCF9H5X
pTetIx0X9lxHcFfaaPhiW9Ei1S9DVDnHVUy2TIzTCxAV60ebjbcfRdrk8FV/+uplKqS1jOfA5m1R
UaUZcR39eePItfsh6YvsE725JCUHbPJikQjV2rE7Cn6cWNlG4maQCGbIx9fVH6othPkRLPsTua4U
juukAK8Jnb5F90z6DPBWqiitpQ9ooZJkW5eOAX39hFYHVAYmZxUBrjSXifjpqDFYHLoA+949fyOW
+9KqW9UeXlaKQl2eXJLN4yuVXb8fl5FFrvM3fUKURNxzwr6S+bF9/o42MUqajQTmVPFv6Hnlk0RO
C4srR1qSERAucKSiyAvsJcQzyb8J8xSseHM52H4dKdVf0Ovpc7Ri+LXy3aHnQuBmHBFwC0BhDzwR
QBuDRoBwLEP1sOJH9TTNgM37CflSwQhuRro2oOsIHYegvC0eAWP7m8exYE+iz/yllEy6gUroA1Me
siRCR3rDvPE5CPkksraZ2OvwxRJyqoOqFg9VvbsrAZIOiqL8Ribje3qnmE8aBKEyXXT3MTnhwRb3
uMVuZPztPR75Pd/X6PiOHWUC0yInZ8Ixq1Cez9NUB0/NA++e1ppEoPQBAhE15dPVaUTVlRaRWnkP
SWjUbod0l98qZ9Q7uCVZZTUychR7gdKNbFUmMWqJINEMM83ZWkTRCbw1qvJQzy1e9TpdWGML6D9S
/CNsLYcYhkwbHg65pMmzqrHRoWIpie4DN3TALiLgtKCS278mYQ+IYucsHcecqMQ/pb56AXPmMXSx
soFLZ9VH4ttFw/6ssoASmiHAwDcXgRtWhyx8SGtG10btlW6j1+D1Hk6etpEINbZ1kQecBv66TqRo
DUhHaSBgvhtNXUJ4Ts7kFnSdysb8MO8ewzZalQZ4AZFrlQouwkMavjkHYo6D8j43cbzmMu+2VfEQ
PDGb0RFJdtW4TSz9aHrAbQW4zmhdcRu8H8PcUDKXLZU3togtBvOwz0GDs4bD8RV7Wm1quxCTcViE
eCajvkoduBmnbnK7HIfWRtaBErqdKfAfokGb5b0Mx7EMEPTdOXfcqWpHKrrJ1aFwbHSh8Y35HfZn
Q7phbkAJ9E8dQdR5dBrW/bebO+TINOW/LqqkdWgqJhD7aKkOeVuw9H09H8rJlQlVvKj6jIvs+0RL
eMdS9kjDD8uRA/TurgoQdNbKs22E5NHKRvmIWOFGgj0xv6YZ8HI9stf1x4R85MqyVx7HuP7xylRC
lPI3mG5XH7o5BTN8cr9OuhKAiSA7DhxkiXsqac396gXGD5sM+5HDZNIT3he5qmjdnFNN/Ru4vgwL
IAwJ01DFQGnyElvM4xxMv6eST4OmNYZ57odIlBMUbBzc14/Z7hbQEk16OUQgxCfo6B2cY7MO5Rar
tYLmQpxmzw+6+u10p9DAC0o8nwxotvScpSTHBcuwROri37fP1ZXFux/lib8WvKklr2XcpIX7FJaf
C26HpxFXuBej0nGh+TjFiPpQBjmyCUYQODMa58Dk1nM9v7Zkxv5L63owYREfGTo60Z4g0N4Ay6/s
y+YO0NSVhZSnrQwrm8DbWmK3mPGAn8NrKbHRMF7+oeIDJux/6aG3fI8eZDhZqNCo7bA1XI7Hm1PF
zfkUPHS2Tpj9qlbNXhAb/Bct1eSEjVzXRcSZ1A0feSqbfemPiCeRgHc0+j/+T9Fjju+rBBjvJsPy
tvFg1LPrAD1ulSW49CTJEWgtk13KYH4a4RNO8/4HPmnc186iVLRNjhJDvNsPIyq6zf9s2NFvWA/N
oCmmNO0UK0vEAATagEhdjTQ19qJQbd2bFaDneXFhrz16QylGLK/lXqqIXEr3tX9WGg+ipJPpYs4s
3zPm0n1AHUrOM4snNB1xIGgl42tAumNq+Gzzem3xZb7d4MwEPWlPwDMeQSgOy9f+riksx0EHNqOO
YP4z4sAFFOUlVZHr4TIxbQ3Yb4Gm0kJdWAIkoLn0s4EEFfxOJPcrZXHmZfG/czwIxMJZ4pzLooCC
za5JsOMu7eCx83bVtHxdrxKhLnzo0dtnYjQpw7RSthjkbYPeGAPX9ZentLoPqIq8TxgP0Zc870r/
vkgyamJRHK/k03SSgUBWrYwiNYJQKelITKe8in07PTs5JOXAKtQIx2fadut8ewn8eOBOe34uqJYi
7JKXAVgARWjeSnmGie3Q2DpCzHxHPsc61e/2YXZYe57GJkRiWxrUb1sw8MyXQJO7Nkw1lQn5u1Jt
OqSFE2yJqii1/pitiH45DFsB5dMDFQBcleHOhET0adMitl42KULEbfi0g13qRkPGnuir6J3gXlRk
/T+UJFAbQQBYXF55c46QReOd+37J7Oiqrqraqko6wQMiF/Vy6e2Ri77SPLsEPTdcprEVhljqM4/k
A0A1QlROkLhJJe+Ftf3mnwrSmTNI5l0Y8jxmXgW2L1DM9+9TTuHqvxwhHqvhJdiauvSRzdS0N9wT
5TxRe68i6xSMCSmlEp0IRtdK9Fcn7z9fYF0s3L1UlmBobo33qyEt/aQq2hI67CeVRi50IDSk/NGN
Lb0kRB0pYH0UBprXePVaKOduKX6Qsq+neN2UR1K5dNpKJhNxPTagGoV74MvwylQekphD4BBDFyCG
YvS6NnK7dSfZ5dxKwSi3y6q1R4zmFlfVm1ayV/T7/ifvtVxjHimWMAV6a8KO0pHn28TSID3mXuem
mr6m6JChBN6LY3AL5fYAchitB4NCE2Lgu08FCt8wYiV8vZIXvI2v0s/i6vSygh5nbkYzCD9PeKgI
UpyllQB/M8uadL008EqRdNZ6q9kSa5EbzvGwiNmVxKmL3uCSkMOfjDquk5haeyLPAphzEfrwFjd/
9qdPvCZDRSlO0pHs62JjxaEP6zaRceJOIKntvWhHlb0ZxA1Xbf+FQ4MIorq3xu7+Nk8FBjj+boh9
qIjM6F9kUIBvLGUzrQLmfOpU7OtxIYVrvJuP6/mw1ryQZTYezxFiB+carBoLCG2cBRZcpSCBwP1t
fOdKkJaVKwyj4JMjWCANjd6ffH/3hFP1CwhdoSkCTbLugk1Jd7tqfljoRkH3cKTdYQvkg0yzdN4a
mQ+3800cpteIAUGgJVizka6FESJ3BiyNvDwoskuXvUXw5Xpu90ov3SMGV7BVtb510TqBJxup1P58
eCvprLL2Y5+2xrWqt+Y9kQiyf8lo9rrsvOlgv+B+ilS7skC+04yLL7Eq8lpgDlyu6N2wHiIXYaGY
6gGzEChzvXNdLWBobWhNb9rH4ecU6QbPN1DROPpvLyxLtrFPFKhv+Fj8+dgA7XE+PL4vk0snzA29
SdbrTTlE593+ImvZMPHgJmPcVqRveDzAc8b0u6ss+N9SvambZADWg+J5dcEZvB/jJAYZWjZrtk9z
lQYq7UU7AyjEhwAk8JPgK2FNHJSd40s2bBSTGFuvFKr7QZ4uB3bJKx/eSCtW2mgy/dPKtwncNdzl
DGA+bllm52MwlYAVt3SiWJ7bmSPfpNsdwsaz0XCV7nRtvF5zj5cmgYdUBLaq4b0+bw9+ZhLb+nKx
FMmEmaqygQtyaNBNMkYf5ErOfA7o+UnQixHHIm/L5c5f4W1P4tTePuhyV1wfXuO/xYbXvUVFz/P9
HnMwDbNSgfU333h8rNmVemsL5rSzEdQfxmMGoErD6xvYKZsJwPUhcPr+1OtUdKYw3jljc59xmUL2
hG3R8Nw6mjNTu80QpjcwZzpHAf61O7O3+33sngwsGwAnTi/UwxGpj1aUpwulyA9wnHIOZQ5CahEP
A9FZOCtVQHvOvIb3ITdmiVWi/rdTTV+ja76JBVSjAagWeO4aS4NqunA1K922O7W3LaMFty6TSLvA
52e3wV6hOAcR1pJjxM4KGrHLqruSuj8NOIoN19OJ2COX5lS/PGmhvPdPaxG+47hEb7rJ8Mf5NhSS
HMezAop372Cbsr4GO8owGgXWuD5uQiYtOoyYSzSdiQ7tHJdWcpfz7oon4IMRNOpow7x78jvXL7ou
+mxi9AC2wu5/d5+8PXetpObQ74h4z9d2HyNFqYOnC71mniGmxt9s5YMAptL3wZ09NhBdrZNtp4pY
i+wsx9MopJhhOQV8cO90HsJ1pZkZZnws/9v58u5lnmAMpRPYdEQXIFeJvTvZ0LzCOSlAcyXWS79T
/8lNWpAKTNQnnHF5ZUa5OmpFvQmQbwA7mE95xpeljj40OAR9x1Wd9RVlfxIEVLyQh+/nNyfN+seb
upQyICb9l7Z3cFoH7m3JNZb46rfn5s/e/grZ/1sOXz5wEKP8+hrsx82ptKQ8IB0CeSGOmmHF10DR
Ufi6F0Zu8iiRdVztNo1tFeqPl8VNRuJMqB5DPsn+gsagjuan/VZaGyVhjtov9QLRD2GgWS4ikwTS
ndo81834d26cQddufEyZ9DPzQK3+KNTQM3xFqE+TDn9b3acYbzfji9t5caM13CT+2dLiRuLS4JfT
Gv+tsCKmzIokNS+5myUsg7BJxH4N9vIQKQos/0/Wpc6SUQTweRuQfNvpkKwm/o12d4m4sG31b7gC
JSBOzOFwHJtHtcNOnxPx4QfIrx3uHP5hqKLYWnazcF1kQWWygbu+bMxTJZ62ODANvWWdzA4OAmkv
opn6EZYgj/kBXGUz6ZHQQ5HUjsavGui3jp98UyNzevIutNkb5PX8Zt8cffxvg3EYPx+WpIN2Tfn6
Cx31rf2pfAJT65gQ3ccEXZg8G1WC6VpvkAkjhtAj3arx3lQHfqtn5ecejjfFiJ8CADxIQeKwisUk
s6zvF+OpTLbBN7dldlv2777C/lNEdRBGYr58HHaMjyo6cZhT/U24VNjA06+HLPcUL9lC6L4n7exW
cPWnFfSHPC+1q2rUj4GMEMqyQafHvSFAKNRrt5lj2WhWWfXI/cpJmFj7UONdS4I2xyTrhmUMY7Z9
BdNxtpv+NnK5tNz6IwFFhRhGXhrYEINZ4LBH+/c1g6WDHXYVuXIuirwJRWMzR18YFuavunrvhXHw
Bp+o0K9omzLYaFALqeYUBc5ySkUCJB8tIGXEEH7KeeFbQr94zsjKSPhimnaUhv7tnvRfhMh/pDRz
bwXkI+mSuSNa/B72F8eCZJjmJhHNkin2fmNIgdy7qvH8n87dIE80coj+Oh1hIu1Jw1Vu6IIkhaAZ
DPUrCyEzn3PeawFjB/WVDbuPlA0Wu8zIQPNn3VfePYvaz9/udpflpZfDL6r6BBQ+m+maYPPYGHwm
lxrDMeCRu6wl1WdPF6H6HD7FgAnPr1zghnPhH0gPpYaXZk9CK3rGE04v3leCZiVx+LpWVHjlnK9r
j0NEC4NzsX7Wr5vr24k0Q7L+wBKGriVpun/eQB5hjjsNxnzAKkF/H3vPz/xtNGWJ9FVa/DkzE7X5
EhaLqv+w4JtbjiOo1fwiiYxawJSqMLXewpg0xdF1kRv//ESD+X+AiYbmFjpGTtzhj6YNbNKfGa+B
c05BImLGXZFQChhE2fNESb3iyEx7MWrQDATrOHBGGeD/LHRRBy5h6fe8UbUJu4qwkdzzdgan0O3M
kmZQC77JODZPjdPZA+jodJZdjeDdzssYqhN9I3ub4cRsnH3VtB2+KdHIwaOjPiQnsOIdGj4EBwS3
fh28VvtD6AUSy9lm/Wl6PN+QCakQanFGL5LwQpiZwmXz9lKn33fWi1XqnG1HYHBDktgY3WGQiCLE
TYYex0dI1OYZbY8jTAxq618iI1vnvY+kAqokTOM4GI0+pseobkqzuKc/3gXSyOQo4NryB7QPk0g5
HkimcqEJc8A9wNjjsqiet/W59JHBEjas5gFQ4E4nXorqfpR/ITcpaJwG6a0Q3Hi+0xr03TXdn6Lr
bj9mIGZu965m9b5GgtR39GUNREiQZLQIRLXRca+Y2km++OwXmbnTnzwqTEndegSG5kxpD1wnyRge
ZqBRMA6QO6EUdrbkEpUsp38hNw9clL0PWpf0jjcIVyPDvlJWF3WFa0qbYC20dX5AnKGr/Y+VQiyY
rZDFt5DjqRPSNfTvCE49urRrGARgcV87wwcVBKbJUk3CY4U8qT7yjAUMpu8el5II3hwbBkxltmgr
oLqoB9gHxKgTxn75ZXmxAv4bUE/7OZucmkmTMjyXwv+NAekl1rMLL1n4zym7UZTPECP77bkNZorT
csRtLt9vD+FVpkt2JTXdktiOd2eLE8l98fjdCvR4cHjJVJKnJWrTsSKKaWWM5RvZpVTN8yK41g9g
sukmhPdGJUxBKfOmnR6n2e+kOYBtuCGyfBDNyyMZicozyHLl1Y1BedUX2MbbkjZhxhBR8fExO8li
KrjwyBVdgRl2NII071GuKb1uSlLyPolUWFv3DXmRsMD0yyNb5I1cy0DaYiwA6KRooRcQ3Fwd63jV
JK8GCGa0d09R+7Ansaqsgd9GMdGcUw6LTmWurWZ3ocUcQ+TsPYiRYHPHR0SEXyZxfcuSuT21npia
TFJpaOV+odJP4q5hgTxOBqtc7W8Ia3UlN7WnPDPd42B0LIfjdN5zl+0uN8RVLJwHPULMruaoz5mZ
kUoQhlkJ4kncM7eWLRtRktKw6H3y8yBlnnxFK/beAyBKlUucv79xcuThaoZDmYlYlqAO+bXfrvnv
vlbNkcxUDn/gsaLornmc6k0J34v1q9t7WYPGnLkkC3/25r5njn+9dTsCzQFh09bnVDO0+Fsq4OzG
8bG56WpfOhl+tAopcRw1W0N9sYFo9rHIOPU7HzV67g4jVRYgkS2D5p27x9eJFpggzABBzrrKc7ZO
n85dTCI/RGBKT2MYcxr5xcO0LVT6jsVYfy1FnfpDNNZbHSBwu7iQe5WPOSYB1xaryS6uNjuCCCpn
Epc3eWDx19upyqcPuQN3miRC+i0Jo06fA7lo6/1YDH4hYpLqhMuWVNwWsuT+Ox9V9hPYfwDq7dti
ZrQ7vulkDCXNlv2Zg5upA3MZsCtt3CV6qajp5iO3ZpNnXLwBYP6IGsGF/ubqPQHwC11jSD0rttU4
ddOIwUG+149oWZr9xbn0sD/Mp/nEMrv+ErBF2cGCuH5PcU+a58JA7HN9HdisUnYEki6r+0UjMYzq
eyJn9vNc7ds9iWMIW5iNClywRTJrRvwFsa5U/hoTvuN/FwiKk6oE/0+iOTL8TE7Q8nng7gYMOb8r
MvAvNMyVZhaQoYFPaMivgstLSHwcEQJlVPW9C/VTwfm6+wwlgJpPUSa72VCjtGHlvDKrHuGQBNfL
s1PR312kVsMwUMmcxxPzRbG+UN9SjyxpG+Bv0trAyQM/UrNuoh0O5R04l4WeZqw7sbSPZRvRoawx
5dYtBA0jG/g1/IAy6mBPWl4pF6T3X4m/UI4Xtpcy0o7BvIhFVBEbcxUIxrlqK+7oiNqA7HXx17NB
k09rAsx/QKat9n0Sif7D8FufqqYJu+HADKhz4/c966Cb+DRwaiYvAFQ+9rrqN0yaBvyN1zpnRjab
SVlVy8fJJBanEe74qWXPpWfDGx15zY0vnQRWULLvPj0y3vwVuRQb/7r5T8aADDJ01NMhIxSIXYiC
l/PcLDNnejBF/Ct4cJIHkitWvzVh5F1YPIgChstEo2PrwBaW1Fn9+6iYITs5nZaHYEWkBKz5sNfD
VRYYJt0WkDFf/b+gewIJ/2e2w1E2V0wqWt6BzHw1CnTM+BhWd3qeH+iigjw4AmQy/4MeTFg5Gp7a
lVKA60wjFa5+BjCB7eldM9cFCqnz02bAYR8fEc9itOKsZjrBqEFhhw9+enDRzJXtc1N0Yl6SUyl2
s4t9hg9O+jbSwJqaLbSCgUky5o/xkmPEssCA6BeiLcg/PfDMsRMn4A8ozmHfRM1NHJ5iOv7BgMsE
Lr+dC+Z9dzs/Osty/npnp+UFM9sg9qRFQeGjwfSpuycvMAnYQruZ707ECg6bRPX56jFdLwo7PymE
1C/hgixLqnY9MZoNQVjzq8lp5zRJYm6Yd8fPo+LXZ6j3zA8m2KX/BRiZMkjWEata15u3B6jh49dq
s4IUlPuSnhRTD2G11TMj6UYvrfA61cTPJikiqCEsD9DALKZND9ImbbygDComEats6J1CFVduaE4/
Cgm3ZxgVoYEC3DHbwk6WpzQKRhIA/km5yzQRDnvpDsxkUvecb90dODH1PSQVIPgPByJ+JvPFw1ZN
1ii8Hk0lrZygSemFIiIFL3Fw4bPRjffuCvqzwTBc9ckb8BAjvDqKt0j4cosmI/XO5+9Tlc3QXQrz
CyFbz038bw7wZmgyl+BQMnOK5KKy3Ug4co4PbbRDCilmRMezlUdf5XmV9AgXCL6A5NMP1QXHjwbK
YKIVvqwnDfSufE5txwoCAcR4Auzi2HbOQlZXB8N/Qyl2hizWJp1svFuE1AJouxpNvj6en8CwV2d9
fm+26Rb3qNfPEbbxgPdRKd2jfNxnUAXsdcx/LspMbCTVpQwDsnwYdnarFanwfgLh6eK6fXIabBIQ
mDgy0uSS8nI+DmOrC+g09KdCl2MjwkVlqkx3P2ti04O1XTp7Xy2PHVxVL1VXimWaCbjN+xo/o0gj
4K0ArOINBsED515A/6H3c3a+2xqNZuiNgsUGRFm7g+UIfyJ0kQSZ9lwbnMI3ks9BdB2SNVHlkBIl
bG56OGlOnQg3J5o/tkms9SJZl/NdS2w0bFLs3/OkNHP449XnziHY3sGiqNFqDrMmLw0XscU/fWnY
SOFjiJtgQ+pstzWKjlKQzQm6DIEwaypx1Ltu8gk2IczmlCxN57ik/HY9JZ0vnsyNDccJz68mxKN5
de5YGqCeC1rT8a3j8ofwqdzkYxUyCxPBGSC5ZDGlM10l1wSz3OPLEFUln354AxbLXTXb8mon13Dv
UmXfZPogiaR9I0Ub8uEtXqBFQemHIlQ9zb+7ZbLGoxrotzuOFYJvlKcxYDNFC2rItSBrQ8uGihuQ
2xGdV4BrHFwcjVCwhmgzrDVeKWcelWMV+hRmBRa9QDkfldbH7GDtfj6tAOC7E+E1dCqpFgMvUJHH
NuFC3SlFW/lUuyuemtjw89yguO4dWvV0D3pPxa7wokkkMd22Dvj8n7qY/KQ9/sS58LwemkLyCWf1
iXs4r8JfriS/B43WVvs26E4KRZWrxQ2MRlqmBJBZVXqgiOYt52R/7qpgWY8PkHx4rYVwyQc98Vy/
ctzGktroHiQiPKKvHaeZg8v6yMcGmuyEIb5M2w5wO6PfTyZL2h8qWmmJQogn34UIcOOAsRUECJKu
lDc++WxrQOO+R/BhmG+Wyowi0/8CUUhlBWYlnniNEglclBpPzQuODltoQeSwwPWYBtQhzES1YcEn
PTyuXitEpYdPRSZd4pehmSArSg0trrrnLgn1igRyQtoTtbV2OM4MVKsqgV0TUosxB9BU/Pbd1ufA
p2Ir84fwx0430dJgQwZPfWfpLud5HzTxWDE1jaNG4+eB2QRobsZRonMw7dRwgB+C784AYDpV2W/7
39H8+jCtk3FAP0zp5KL1zEU1nJcAts5LHGAVZRHCBTRiEkf/avvgOoN5Q3FLieF04x0Y0bdT+4rq
ukd3sf7NGxqRVaRQN5rwIkeH8extpOFKTZ/Zj95E4kM3gnO+c8RZC5MSPFe8z8QENqilHZE0hBZo
SIgOSzqCieRbWOfU0SqfCHrM0lkc6o3qqqc3dlc+JaVcWSeec/QjGCUE5czVC7qlRbsovpNoQCeH
wovhTXVM2T0cuEIEk+z61kFc1DLRlHk++V2S8XvkYP0Thl0WBcnXDluBJxJ1mQlh5Q5z1WAGjdpN
t1TFXo+lVLaIEI+AQa1c+KWDMlFKHUrEFvv3k8SYAMeL3YaoORcux0v1ZDz4+nJNWcDcnL+S6qvM
8lULv+/gKgtRBakULeb5l460VqgcIK15fUIMqfQR1+HLhqEYdnXnp43FEuJuZR9gRJCBgUEm+pKF
o7HtkdYNiJPONecagOvHMFvF7FIYdWShZGiR9nKBGFgbeHB1J5mVAZopJhMQwdQeudEBIlitAZ4n
h0HiSFG4HMy/YBAErfzWQiXgHrGMs7W55UFeWfhrHzDweyQUHCMH78mvq+IBzKTOchFKgTAEBSBW
i8RmNItb7wl8z/fl69dIxkfLAXO8I0HouZMrY4sWSigLHAwSy8vmivfmOiJzsXYCHa7VWhgAYj3W
xi10q4HyMiKDg141pYDg/64Jvik3hduwXmh/I8fPEUZlviIudTvuiqe8XELhhhhXe86UKdv0Lpip
5GODWMhmMWRCcd6uWsJC/7rJ+1HncTZgu4aViCeP3y6qFG3LcVQWSD++371bDnsu7odTMhxLj58H
4ImVttplpouRTe++nIu7KMALqt9oGQzSPxmViwvQlxCazydA/nPCxdQKuvca4c9gnPS5Eu38d3tk
qZQLQmka9uHo/wjozG387dScsPQrShWADVMePFU22oXewnKNQSMjRxWYnI6rnigTqDuBzGG8buUs
4HcvUOw19uxGbolUxqjYffe+5ugjHt4kpXDFD892HGNGpY7uK/9HRRHtiZ3EVRhw9nGfaenP2uk4
nEJodT8X0JSd8cy5E9TQz1U+9o9WN5o77elOhpL4h3PIWGC3+R4el+Fyy30M/xvh2Yy/1YNIuFw8
a0Iejk6IhsR3+NMi3RYN5/KOkyPn8KA3CPLYwY7NhI7o6dn5eqUKvT0UUjxRzjwu+qq9HrlfFx9u
/dbLFf+GR5mBnIKI2FBOxDVJWwA/cmh/lIQId0iMJOBAEoFlUqPnGzE2c8OjjkkmrT/njMu69q5r
BMrhs9/6FgeD9999Rd1SDqqoByFPc7LFxKE8rqEKGetPG/CBt+8t5P8jMcl+W8Z2008dLHeNgtaw
OGcksBeLMLFu5wZNBukrv6JCkaLREnYYudOZq3pU/ag+w1ROB4kQQX5s3oDSLAwTLAYEaBIJD4W1
mtim8SI2trPX0GrPa5ByvgwPIwsCHZsB+A3une7M4SMUoPjuFsfQ4DJ/wFF9+p1Wl1Ng6EPOQwaK
lhqSseuQByviRrAL2qg/JOkBR9+B+XQnYw6WqassEPsQr4lG8VMDvnTU6YsgDqLDy8JmT03xaqRO
9nGm+9CZhdnP6KDLZTNMubXFUtkNC0UpHuyskuhP0mK2YLbLWb3ykWAYE0AfiN6hdvfPLqoAXSTA
P7Y3qUNCAUMCq+TxvYVPQnU++EfwSwgfDcCg7U0W2bLqAvYR2KxZdWTrQJ21AIDjj3wEvST3RlLm
vexMNdLTxOq16tnY3vNJJ33TcSIs1WmIsqQrEaOzNkTM036ukyGdd9pTmr9wEAo52Wf8t7gVOsZk
VOHJJ2zaD4sOj2xvtW9SH/p/mNZbJljyoilyZ85/jGsdr2w34gkeGlGQOEQTKLKn4awFCKQ5asEW
3hy44r8S4l5o0VHQvLtpK5QzP0DCZzBdiYL3rGMfW2B/qq+eQBerqTuzj6rByl+EQaoQ8e4SFXkX
tr9rpRYtxJNJiNzuwTJm0G4h6ZSaZXNBOQ6s59j+RHSlis5qang2Wjv6k8o1UakaK+sAvs18fB0L
BSCAE/kY/Wuk6CFuzN0T+qk6RbEyPxkcT+LUXeI27iy8UF/MdJDmP3cqnYn8OEclWlJwGzFwB/Ek
jr0X/lxXWtJVGTWivCCMQT6GjlsrUTL2pt/w05lcv7EEagR1h3eLw5DhC3XR18QadVuRKiGZJscp
d9ePhkOu92OCqjI9B9aVz/g2qoaN3XkM8GIDstHP5ePJyIafZnJwxD9XKtjZc5+85cdE7XM9n2yD
y5nP+LNOjtUjryK2dUkfeFkMMl5iBKaflJM6fsUDccZAIOXRHCSrC+b6bHbXZvlehLPNOygXZG6E
obd1nf9Q42vNtil0v0FZL191j7x+2tOWS3sYk8cxT3lpS/gaJ2ERWQCZnqsBZ6vch4W9b1hT1fCd
Z2DaaVDWwDkIiZD1/YyjrHW2SOY6PrhwVIfZPKSmT3Vd8FHbMyzl9bn3rLrg/PcM0gPlxkDGSv9P
6c17u/cFEJI45WX0bl4hjcr3YXw1dIVvYlle6FjVstRKS0X1LUyDed7/CU7+qCWn/YaC8N9vFziZ
ZJBv4NhVbGGenJdg9Cw9UFKzlGDbNASGtwCwMlNWMPkzmuw2W79qN4t54N2YBz/59zSE6hhZdsGj
Kmw6RrtNENnCb2wQrdQ9Ye7NqtbHi/O+l2lLuVJzB9ENENEljfWu8XvV+bc5taaEha9Du+BW7FaM
o9PLlftLUZCE2OTEqpWHskJb9DvE2i51YAop7W+lGbcetshscFdZU0HhYMMbiCNJgGxIdZ0Cx0iR
IVzk5GmeZFg5/maL4sL7unI32MYpbqeUoI3bHnklu9JBH8dorfY1v4yLBSutrpo21ksgYsVR9R3C
3pRLPmI/uUAVy6PHquz0gQOu4pDoqltQ3nlwDNoHF2Y0MqRAHvQw+cImIBEPrEei21pYKiQnrsU3
25l+Cc3xMgODH5VGeeppDDlGKwQ04IrKXhEzfPH52pOqWn03OsVBn7rAL4wCNZ0CNvghLAoiqh74
FVn1YjLR19IvmVvsLSRKApJbRyRhzzwlzspbK5Md/HKLuAmmuILPUcBcLvWzykTJGzaV6qkd3531
nkJ/vTlQdpqHQ5t4M+HjGJY49yjhrFN/ZuGkawUn67BVc1o3pGDpIIr2GfTuoBfKjY8ptJNMQfUG
mJig6KTpkTi7xU5O2RmDVm6V7Ld/VGWgEzqDA6yy81nLlB2oWOLeN2Yr1dWBXZ/ewH4+qNDpKSzP
RjDvUa3gZ95A3OcEe/z96OJ3mUrLHQAoI6O2DQdnTQOivqGAaYb7iQRl4Frn6x8esW9DBgdg/xuE
GTk5e6cEM+HHtgObm/CORND0jzFbku2zxoQN1b/omAUxCFF27E8+bKhV153UhcXJJNfNYCKr5zSi
MTcATewFqyLi9L3VrtJ+XtSozCJrFJK/VAFiGtY2gDo2LQOYxdKQekOxhG4VnmKS5tJMy4Y4g/Rs
6zbbfPm2+9hMsATvoTGt2iLmJ505yr2zhaSacUfV01NEwivCNjaSKIh4l0YkSswcRXZEXW1dz1Pw
HnddUTauYzCyec0Yi+WuNEcfgUkYiNjm5OCuFcf4OPGZ7AIUwx7LTzDmTP/vgzlDBtpxLgmzWHgC
cPnlfPa4LwSLAcBMRbW/YcI2yUyXNBYsj1ItTaZKWsRyQR9vOcQTegCLXewVmvcSs/INEq8Hn9qw
HWoUTQ5/2oMqykqBOwzhHTodOsQa05F9QznLqWjpaDZg24PjbAaj0jgaozvteTe4Jc4M30BSkOEf
pMKYwyEAp7LzOxlFLgT80OpBBhRG+weod8oDxnJMk8uiQKH/ht4AwSwZ8czO1tvoMfK91LLjh+qI
nnJ8ng2fXTNjrVhin4Gdn33E6Xsro0diuel89rfaJTxoFBCda2YD2uO9Wb3BnHD/YE2AJGML9z13
3NiLoSQsjGsnrpt1TXJpXRzrrYQBJe3hD9ACdgrdiCg8Rk8fmyBAAZUlzwzeOVOZp/YdX3w5HDPc
ZfhEN4xO1AozTDvAeisO5H49YgIYS9ntb1Doscdn8oOHrhAn7xSuMxR8Tr/cqvst4OLY6zhPMNvG
4qbdz0nfGgPxfTM0L64QwbzqluNpwv4xNJgJK5CzRdZTOmc7f3l3k5+QxvKmhH5t2ZVgExRwEWiD
8W5BtOp5WqnIFw5olxs6NI45cH3LEA6VJTvFs0fSo9SKYVmoE4Qn9RB9+YhmeV6V1neW+VlbXA3L
nqHuU/nVL0SqGsGUejsbgF5dbY/VSQuDTpkXKuc6Orp+bpXdgLCox0Ebc/AKFQXmlSVgOJ9xWGmA
2842yqmsLoNsuXXW1wWjLUhFuKKLQ0D4UQ/r4udop3CZ5/rm/bCRMDaiSJmSUSe9B3UtrBIcKbtf
HpMMuI6L1CN9Y7pcsvxchQqDopI1yRqz8Jq7fcqfujZ0tqke19Mm4XyGFH8H4zpRtNDkrnyEwFMe
BbczcygC1S/jTSIhwyUrxLaRsEJXVWOAdJJFztQXw0yVBhcfvYeSiZupamRCohJyGLYlyEuA1mRl
f6uD/gULWKJ7DMwYFQ0+ViiS+XLvNZCB6K1YfaDC31JSKZoASU4aZIP5W6e6AcTAoeBsB189f0Kp
Tazq3QTAiv+v94eDM4gnjAhEOyR7mTPc2GRkNWU8OR1DqQz1LZO2o8iVNtjIUAe78YSAzw9GEo/q
PvkvrE0Yb0bCFEzTU8wgjXj4Lq3mA4yBmAl6qOu4d28iZaThrNcbVr0nbxvnVW3WldyLO8yt+isj
npzfzqkYCREtcnNasj0zZfRgKZJlq0kSMNQtgscyKKUuWe8Aa6nCtk+iUj5T0t2Mo/SZ/8Gw36C/
SPBD58QRdmD5m2Dhbw5qiIVD3Riqd2MxDf1wWwuvWsEG2H9iBDLHyU3Fv0+BlsxaQEw1+pO+W3ll
yPwh9jq/zVbqPCzVafvZAOGmPmwD/t5awupg/wPKLwQuc/SqKlzcpAgFavzVrmPS7JMBJhWL9/TU
P81BUojWOZnOKR8PG8LBgVZ7mVQEvKAPiIBfH1NogLOq70TuuPyzwiqv1eYxlx5Jw9Bl39HtLxTX
8tlS2TcJpxPcSuO7dd+U+Np2tZkj3hupJZ47YJt5JOeQRVH9tHnadwCYXHn97+ZPF0VLh30tq9jR
Eamlus6tBrfXmu1Yt4qsU/7O3+ICyP2xI53eQxUyFELTUjYk0ZATuEF9xRjkr74u6FSIOh34xjFJ
kptMQ0q9HuyclZ5/sJmdiTgz4AG1GEa8hKpGEv/C56EpPrAl4bxtJg1FFKL5dJ36jWpZJ1N/S1b3
y+lXHxG0feWZzOKijVIiHahN0NnkubhZlXW+Pmcj7GdhYkU74HRX+M2HvnwSce3CglpRN2rTlhP8
jZtj8MXrQjxCfstPSSXV80hbIZtFxO4mwH1HMXSjTMOGmgjpAPj6H2/z0ukPUh9KVy42OCremFov
9ClcysqixKOSpqz5UjCMGVGS070Pe2f6YAlEJIetEvgGHrmrXRgjPVkGq4FE73oYb12NSW712iqr
Otdm/0i0RUEXIpfnjfgVFXQC4BjoNJuMMxQa8tzbDq43oUURxhHPXRd6VbBKQRqrws1IxJqCvRgB
TOLOQ0wwODxTrDvjZy9xhcDN7d/ipErTRNlRaprgu5u1fzFYRTtxFNkKvq6EiHDPbZ8uSmLbaUnY
RgTohg2pOwyvSIgWxbfdB3T1tmndNJBzUaqcHl4EKPFs5yq2n+oE/gd60GSQW3DhVeBzfZmaDsMf
3EawH0XGpwBFBuHTjQxKGNl/a3iMmBTqHPtLAd9klIf1ZrolOuJR87A/WWbsl6TWxl7/gJ/AjW35
+d1LNQikiUj0cyxma2OZKwUwbgsKbRmn0BpqG6O3HP+qtussDtMa7FyJLIdTqeWJeOnV66tagP0c
QFOq2Px8S+JewC87AhyugoHcM6UCtmY1zbQ6ScA2csElSdwT1ZiVoDcbvGmSzx06BesqlXHILYY/
cc+PDp7RH5W9EfcgG0PNuV2vFDUNmNyqtWeuLjJH6+R1Wzz25tbrBJ395P1nZ3FXcAY4RsYdFsKN
jtoGOYqeS4rbqGPAGGCcYFYSg7XpMqZ1fAD2j0rMtfSFFkQQdDUodbldRpyAA1IX8N+ZyURLO/P8
dPh/srXVRLQScuuDRWrc0ISJGLCru8Uz0bV1UOHBvQBzNGIIUoezGgQypAnoGg6uMTUAdN7bs28C
9ARsBu9nb6reTs/Q1+dIjdk9Ham4F+vEYqnXWlRvBo5eyxJJcl0j5MY4hh+n9uI277/qb1mWA7c5
XKIHe9zWfxypgdk/uuRyVYh9y0bLWKqIXPKQ9YsYOllI4y8wk10ArtRqM6i4AXR+Pl0CQN8+uGh9
7pKg5z/A6o5X8t8pq5sGxA1xb0uoYP5EaUQIUyz0HV6gAghCxDGyCbPbsCZ/0VjaKL7pw+nqktHT
RsS7ah4MlMSrysYBcfrJ9wEN8aKSa7lBPQkTPVZ+PtPhTpXlB1heZQC0FoEBKkUILBcrgI2YrMK2
3IzhNRhvplAQfD6J3ZP+4+JQUfrB36m35dDdv1HCz3T/3JlqC2/lfxieqAAvCtSdO2EPTML6b2Sx
LyoPp0zniruGWb+TSTncqJu5YusD9oin4kUm4aV4zgx91VG6gZNjF/XMgNdgL3vYPe/E78J8jtLK
FnfrM+foafKBXa67sa8kTzD0r/AzGQVf91sBpZpyz+9A3LSZL+jjhQYrz5n3+AKt5NMLhcYhXYpJ
QmUWNALS7A+jTyEAI4WmL0yA79B7rlevKO2yhd3+BzqU+QgVHF1CoE/e8RcW9ovKm3aO9JQc+hyU
l77A3yv7dv5z7FzIMSrACicJrK+xVKuKSW9RjwDkOU5cDBY+YGRpZ5N3fXcYxKfgg00LD31te5tX
liMoucy5fLIoZZP9+NgGGsOvqnAGqZqSR0u3CbPag9/5UePK9L3LNgtyOAs29b9vxm9ImhbQJHER
i9L+kfKI/fX83nwP71/c2OK4OUOFizAa569wA9i2PA+Z5d+exPzwAaML4UlYVv1gKVTZJ04BPcID
PbOUcefk8xIMfXVH0gQeKHcLv8c4hBsfP79Ug3nEvtXe6yhgzjA8e4zAVXDiZukRfoa18X9OCK//
7Z6MopML0BqvsZ4Vv022QgTgFNbkKl6JKrVG+/wxF5lPtKtEin9AGOvbw3EspGQjgBgQEOT4vW2a
YNjsbqUxS4mSrsalBy1BFWXuIN0Gxm+xAKejPzw7d+n0jIwT+cKhUzkCFBLI/WmgTIdSXyf0IoyH
AXNMbndCGZVu8JE4SXnguZEtcq9Rgt4nB3CKTrSzXyEBLQQEFyIkt468T9G+CRESlAXnjcdV6j5/
1lxTYgD9cEJ/7b8l9O/7NXsYmvhFshPBVUjIxoy+cLBz7x/L8fxMvVhzNqyDYMDV4Wqty7PUIwzG
smbxs9zEjAqEtdFMgOZDko9p4Fj7PGnT14cRM0D0fBB3PBJviib2644maeyxLnjGexz/kwx/juZr
0/mRx7vP11gVcYY5wN589tbgQWsNg7bEh6cE/+gZgPziC8/ChelS/N9duEsTccEYqvGdyGoqKQ33
gjMh1rquR/Iu3ZFiKPFDDdFuUTrjEBAckEXyEiChbsn/VncwJ36RkYuCdNVgEQRU7qx7YADSoY1+
sXMuBarOpemjol6kfyHg7BwPzajCQaeDwsq/P1ZcFY2XzjIpzdgJXXXj4yzg2BLudJVeuFow55uz
yTZIp6MTHcIws+JHCZdMnejpHWUH4ADi4qwm7DxVqJ0LHIB4cnw4VWScgHCJG8OufyNaRO17X050
+e0Q8Siu+17cdBAgj+62tLavizEJIdwMuBIDjH3V+ELzTCiI16iz1lYBIvKrYFWbjSrMHOB3ZDOo
TwzrNyBjwiZjMMdrHdsaMkX7pH7yAGUg8UVmbnNSHXByM/OrEx7EOneZdOpMtjeVR++tmzVQFWAt
O2axz+vM++nsancpw2olW4dSDLEPJEnembnuU2km2lf38Gd4l1R2gTPvqJY42PriN0nxLeqOEPmX
o2oHjsRKaVssXrTiOjWMdUAqjZh06I0OU+rGbgFRKJahOsTZRXvw1ayaf7z/Hyq4yYlBMHSIP7fx
2VP+8yOxrSSJnFL3OXu+gZuvnwByUhFOpiSU/wu6A0b/PvGiGUJrklKRkvSExgvceWHqhWM17IS1
RdLZsTx9FZlt1v0akHOVNflKGo1wdc46N37HZdFVIPsMhkIyzb0+bTp5f03LTZWpHzSz5eYaJEI5
EssjtKcornTZez7CCSvG72gyKpNEu8R/Kl+D50zBKtvmjJgyZZNkxEG/Bcz08uB9zDJeh8XhXmIN
5EzfSPAVUwuj958BDRf+Lg3kXNqkGBIujBCoXfINoEj9dY4v1HLtL6nSqezr8HHf6mz5FKBcISvS
O7S/1qdkBbpQM3L3C0ykuh0nty/2v/wNBQBlTF6rUezG2KlT9VWhIlXwKVTcVkBw4cn+p83n5JDl
akV4Mq5R43Gm7hGszb9/s/Head3j+womKHyBIDeEq89DEhDnBfgNkRTVCoiIQaOUwe+A7jmRBIzV
KP9YmNUA8ifRqYZ61ow8Tryg0dSVJc3mjovTNzFCR5xV71EhLbsl9Q5KlbrrfA9xaUACXIfXF9t3
mWm0/aBMgVqvc393lnX6m2S4mzSbaJN/aCDWDnODHZQy2dHTj+aiBQAruzg2ktgMXINOlRPU4i6x
Osp+83a4G7wNuyGMYFc5nF/BaTM9y7hGZ5WgsnkOyv/ZVTVRGUwFyYU86eYUNRZP1ynDWnkDaBLZ
C93VO0j6k0IwqTnPMC3g5XSsHRiqQekQzOb9pMOWfhAFU4yKBGXkjMOF9QCa2Zc+2OUU8xkjGOGj
KUVbMWfLocuzc9njEdDaj9hMuroTtLSrxtmL6UPW7UUFj9tQ2cxi69RHsi48dZb643jlp8WHdztT
XsyP3XSqjxK1HEQUavGtEat9fPcQxj8FPDnj2fqXVkgP6lY/WsmuS/mhI6rMFNBbGV56mlNXbXau
iLf6OAxRjKpnyAdK6qV+je32/Inmbd2aVG6S0TQSWTlGC5X7p2Ndqtaij0fSYeLo8UxT9YOEn7v0
XBLVQd0jsnR78Lvdelf5KDkr/cCkiJtUWJ7HPOEIL6x3DFNasvPGOwCmr+oQCutovdQVuX+pu4YU
bv3d3O6t+zIxDvlRUJzUkvZLPCH3kGajKioDu386ckIG0/q3vPoGGPD0+A07YJugHj21+anc2cka
CvsQZvbqaDkRMz9moNw7OPRn89ebjKKIIxrPKK1Jd25k2X5giuxNjOHDgGtzZbNIYD9DhkTlIOtw
2196C23j1M32ssu8hylEQ/NxJMOBGnJTxRFADmnl3xsafCljjmg6T/7kX2QHChl0P6iNUAjSF/Iu
btiTCbNm1tFFwspu1LjyAu2lgXdbWB6wwwXbMaZHZMYcYb2k5Lioc184EzkJLPZCsKdFGrW19+AD
y39Xx8lcFpiPqPIayO3bQ4lPGr1c4juv5Fp3Czc72YJ85Pdb6fXC5C3Y9jvjs0ZJoYu3izIKsGdn
F3XUaWE/Mj15yEwfgr6VQK/l4OhaIbCWq80rEKCstHcwhjKTRIIFG7ptPBLs4KN0v1lSAJL1nBgx
FKfgEOT6XUEbk517oRWlA0JzTrzcFBl1c6UlStkDi07YEgWGHiKk1fgj5mtbwGNxGHz1qP8rRTcE
dZ8Lue0pPy4eCvUpfbREcM12/+yOLu5O9ywB4Hk9eO8J//HheLRMIs5y48LzTCAHbvdCXk6uifGq
6wJw+5BIxFJIGrIyOTgONlUvOa8nwYBtgwxq+tAYFF35rsHoctbLcMGlLykBd/6O/6nPDfOiQKzL
PhNlPfnK9yEbXqiZPUQIbE3XKc79qHKLUm/4F4G3ZUGbAhTllbV6/5fXCmnV9iMTxSbF250SMGa2
PUj8fVN3ybt0YC22vyONUEFh2vatIDwK8Vi1xV8W/GtcXkFCwk1pbO/5I3F897ZhHJcjRjImHsoL
T4wlQm2zzrBopAwiHjXJFFhfRVEo3zOHX+mUcyM2UfTOiwLIHCIs6FZDavroVOuExN8F3s+iGIGq
/91dLu+A74cpBtR5AxbOIS1tvlxvvA00rCJP6v6jV+6oxnVnDP+PrrOlmCrdAWaXnrRdxVxkhZiN
Kq0ZBXUIa8R0XYsG9OZcXsD22WCMVFP1O7T8RydBKsw3H4qQ/VnmFeVKA7CpQCHq3yYmuvf0Bzyn
1lqQI2tXFEZmpQoTFHAXZ6VmTYvMg1y/rPv+uNNEZwxSnDeRtdSFc8XmaY9LGwAFaZDjBvz6ehDd
SYDhwZU0hW0OLSmRboDnsei5uH4ELOagQq5h9Ocjo5H75NYtSXs6Fori9Sq5MGWqv8QMwMT6BQAs
DLciCo5iTzxn6gx5P1slmPN+2WF0LeiZ1vthsbuOqMdJFnMTJBqYNXVK9i/amz/W67NzirwH9gLf
qmILVj+GlgPLEWhElgs8bcd/a9Q0U/rim9TkR54r/fo0Nl5bEsO0Ekka3cqJWhBVmAYUe/4U4HA+
khMmSVdSVQooKyz4coMPp3xRphGLoOr7t/KGSOctIWX+g0NHvSQWgO5+OBITAX5Mx8+z4+0R91nb
hz6iiFduCkRrchv7pEgFOCIZNXxEE3eMfJVYdtq+ciIfBW4ejjkang4fGcjF+MYWZIo7OTNCs/ie
MQbBxm6HRZBGi25bVcs7MdAD28Wl+zx9PwK5EL6g9TphW3tD0zMzoyIuEdcmVqyIuXkmgEU7zwNB
sDq6mc8vIVyTAczSP1ALsUPTks0J0odRBiMMs5BipLuZ2FjaElp6ml5w4agGZUel7UVaMRWsCH8H
T7Yg96ZxJiRAOtbl9Grz07+1+r6u1wJSdhlw/ALjSQ3LX+gbV7TfThbtkp7UXzWDpSNYlkLnsvKJ
I7a5Mke5oTHTj97/QGzgxjKKI38G9KwA/c/s7AOKNUVSuqsWu1hWQ3pOTCeWptipOSA2EnV97CmK
gUPDCwazGzYglwnaht17ZRW6902xvUpuNfLveTrJJJ+R3XzvbQX9/k4t0qmSuP6x/KwDqG1x+81k
5/xZPRByxYjpAPa9vh1r+gwLnawwNL2s4Dti83NA4+DNeplSQkK+7o94Tez0MAYHceZn4YRXmeZf
b0FpQi/TeeQfXgp4p5+IGWfnh0pUkWvvsdfigw1S1hin4xsscKrT1BQ3fuYcNBvibF1iNqSgPcG9
E7hio2frUJjv8BMgIa2GHo7P1am64CxJuHfZMeJRPqoiJsboqOOufN9RDu5a6yc1gkKDIwik6/7+
vN20VsX/mezNL8agnJl+17A48u512X9nuSm+iqdi2APEhfEzm+AZdXcCY4rj/q/0hnDMzzfPZ3y4
TFxZz4OE+EGNoTO/kjq6J1ZIL1qM6ot56WeSmvYpdZ2hTIr0W2LRK0vW/kv9Xe6xJ6Wpu5/xbXJT
HKDytI3kDnH59aO1ADI6TicFHD7ABD05t0BJWQutItP29Vm9G+4zxu0AKY9kLDEeQdMoW1SRUXN/
EJQBMwuPmYn/dHteWAYfwi9mWST9dx9PNnnTofLJ/qMn1pGVFVkDXsjjqa0ShJj4Sh2mzdoo6xx6
AGfFSgpd3MdjJwEeGIE2BIn00LlBCPLM4+iL25kCn4+VBf9x8OxOxWx7btUoicnsBi3YnIrrC9zl
lbKtgu0biZ1aqupJh+uwYSE3uE7F5dGXuYDHo2w7WH02981xwL1uP5YbSC3L8mOZFnDLJm1bKoLV
LKH8di9YYaktHvMmu7uORXRh+vSOxYUywf3au2yXln175sEkkfSqD6nmj4ORX6WCa6BVYeIzbio8
z35uH9diJdnsSvcS2mwUGq7Q+a+/M4zBO/c4bAVOkvKBiNgUm/MB/K/L8LEGHIitDim89bATLqk0
4nvpHOskO/Kt/a9qtxq8Y6fi3oZYPatMeDOulMLzKx+/RSya7irS5VFs/o9zQ9EoJx1Wgd+N3m3q
uTH9zVG7G+5WojM3+tSePDqsUb8dzUXlrsEQzt9B2KNSMQK7y9UdrlV2VfQ+6sfcespDnORT3MJm
EdxeeA90v8SSLhP0Y/McsbhCXdZ4SgA6CEn2DpH0qa8Htcy0ASzOnCtF9HSQL43f6LpXyXtZmcU2
X3+SD+KogWW34iUc12X4cvTwNANsp5T5ImNoFIUWR8OS8P/6hp428q6R0Yl0gvyoo7cnPSP0jquz
KJzIah32exRRBwDZrj52ibIB4LYQ6sBGdwNDwYc9Amr+wUPRZpsWZRUJRmOgZtgnDVeaCIv2XAeb
ypUx6i5VGLb+t5+DbeJHXP0b4uqwYUOXPj1sKJ3CN2cw+hJzVQYD2hPzgoyLx3922G5AoPTJKi3a
hlnDSLkftMG/P79AMGnWsiANK6IqnV/GraQVJYNI/T1rOudl3By7exoyKNmzkgaCljDrk/1Dhln2
13L7gahAGz8zzAGYAiBXACR6QeAtYNGUifhpes41rtwVVg07AairzgwkzVyv/8+BlXMTctOBz5E6
JmQWrTSnbz0bC/F5jCwJAMrqv4G7AVsJbl/Hu3Ps2EVSjdeStqbTMTnELlSUmS1dtfd/bkaHEkgR
qdtGLmmR+HC/+tlxSuBgo3i1MuGI1JZloZCI0UpSJGDbFCtdpQRCrVAwYsEDhJngNsgeKFirEwJG
ed5s8nwTPfZs3QrdXfGUXn/fQSwqR79OK1OEKLVo0bdEigoYLqtWiBfI1QwvkJ+wIT9gp046M+Ld
1yO8duzdWVjssEt6LjQWUbOxde1WWopCPrYwANs82mTOPLPUue+Dp4fOc9vuCc4cYirH7kiPbZPS
5FBI5GG4xdbqhYYYOYWn6YOH6ExEg8j0Ol1F7Emb9Tvemt1LUVJ9vt9/omYgrl7EyakYNQWmsUD8
+73XPLzTgfVSQiJl4YAWvbuKeMc9eLrdqA+66OzrLMGQOl8xsbHz5Ljg1dmHONjGevA94xwQbU7/
BZy4f4M8GtzORHvxMz4dUb9VzZiYqLQC0pSUUiLs5817fmHYgGl4gW3gYXP47rDvwDr0ja06txPD
Mjq1TlATKHQaNVysJMuAnE8BdCn/hUKuxHFDkeC3DDSd4Fwm3Ly6tYrfDIZGPDcYTvuVhmUZ+XPR
KKiaI1P9nnM/27YxFyxkyES9ndmgv0aSfGEDjEI4ud2vXrP8sBAcd/5vWUhk4aLbHDR7Vt04sp9Q
YXkD7tJ7b4l7mGMs6EkWysamGs8ZCH16G+hI1uP2JiwlSire9tVqH0ziDgPEXQfshO8R3d+0cFBd
o3UtVSo9kfwOBlxgosjnj7tIB9Y4iXzveUdnzFPGb3DMshVoWxjOBTE3AR0ZlBXzv/+IpavC5loX
34qFF82L51y9XXvmR7opSpD4WLNB5i/FSWrp2xfsAy4YEgtfU6zArHjZoHj8Wjd7UHy6rDmwsEO7
pq9WpbxIJXCrEZMFOrhK5R4FGWcVoPOqH7YU6N2w1mpdKvfgq69oYVVJl9ksiF+Rk8qJMCC4t0wk
1Coj5MeOgfTHYE4Px64By6ZQjX2BvrKXx3d3aCXmOjc08qvZJw6Rx4JQira0BLJL2d3Or52nlC1y
urqmfF4vs4ny3pXLVfVD2cRIsax+VQkSRL/Hk13tlqymbJ9Di3pJIeeSjvK/6yFZKwJUs/NpiLoq
uQbsYNEUIsbPMbPL9AVwyGak0yz+1AzIC3Wga8VMPLp3081XgZqMOY3KPJRM+KF//X/N6fUpMLtu
5kHQaB0ppbUc8UmCjc55YdTbCiAfTudsZJzDFHr8+8qDws4BBRhGa6e5Yj+0+hgb3hf73k8yHPSk
AFvLS8snsMQJ9KM8mUK9pQMVFLzgpp5G6UhNVxXfbh60GURnfNJ/usDsk19GLcH9Aw1psjLeZSel
YU7z2qp7+YIykjXOnfndiM9ajLKv8jRlyiNrO5VbO46wOi9tfRd4hQskDpH4c8aM4dyg3leJICoY
vzDx1YiQnbrrpqd3/4jw40EjD/rsCnfKoKdzcxSyQ9k5UoEM1AOhEC1bHD4S3wjj104CsFXf7hJN
ly2FCtUTiJcrJQEUPwvtl5n5QNe7vjw4L3Dvs62kAMehAcQI/Q6ACoiw7x7hIiy82MDzQOa2jkZ4
J10yopVyIYVZLybKT/oOReFsk2M7hDZ2MRYcKbHGOg0q0MVzLQnIoY98MprlMFKpDqbOo7Wk/7ZX
WFMqGYCFmtRYhT4fk/yVcI0DRL13CU/UQBiMYP0KWxbkau9vVIqbl/te5QwiqBgIdHbi4+np9Cjl
xbOXMuwVJCLxw8vUbMWqreriioW9QmpQQUxhv91stbSiHuBDPZfBSpzhXx39XaHmFp7Z0BsDkhT0
YHZMMHK47zaKJ8WJa8nNaJ7cTEMcmxKyy2RDj8uvfrT/0qBOrW+vCDLtPbrMip8l7aMCrvCBorGH
hZ8XCVaoJqMvcpkcih7vme0w6L4lbfMW9q366gbkiir9Rv9iQfKKsVUBZhBAJJEmWsxs4VLJGBPT
xdxSImDwNbcRkJLLUOoVfbF+vjnV7n5Q3CBfx+mUrToS63EkxAK4JI5KNaaBPHDn/gzuRFFVK+uF
s/7ofWYBdgY4Wqub+a6cYZiPuE0UgHBxfJCV8eM+ZIGtWG+sE0QcA05rJvsKbd931h+8YkdvshpL
Lvt9M6A4qfb5XiE5NbPSDsJb+F3Z/DANe1jlr+4v9Dw0DjL3zwKDZWucxqp7rEgZt6hLUvBDkJiW
nBF7gIblP6R+esC0DWn67bxcW8fJXBWYGXXU7JZTNa7eHEJK7BWEdyDi9AFM+dFeg+N2lOU8HZtc
hXM3HYplz1jzHF2Rc6MwHHMu0w2XpU+RiSKl9oo7eyL+ruPwZRLS2JM+oS69U8kDtQ6G5Tc999KR
CPmQGhqw+7XwYPleWf4XhYBX/4mEjdoNEFZwMJshdpd3cipWBMmRKY+/0sBKtcPRCsT6dymJin15
t7FFO671VT2JzLsaVv3C9TdFmTibxFENIEixrH8cJkzo5o2nari8xilGfvTshhFrAH38ffv1T5e9
iHPIyVCIfpU89LYSwONbHMbUmZ84P3IWt67ZmCfezq3T59+h2RYp4CgrW8MAWNw3njjTsd/NLZnf
G3PjkaZNqRoL3g1CtqP4jbeWCzwUC7qwgUKekrvBdl+32t7q08dmmH+UzVABkJCzbeljwNHKODtQ
lBhSZV5/izEIDtNsXexIp1cHMLozjaRC3rAV8j0ed/Ch5alVfUqSzy1aK7XRnnn1+u9fKcbPxvlD
3XTDlDKBFkNmEeV1v3CC7xcv2FLI36OHdF5YV3AEGaPW2xRHdfT6oCUhKtRL1skWy/vBJ7WbRbRx
aGwdYteb4294R5XfrHW05Y7YTBYDKUDEgye3BhqDagm+zNtNpXW57F+B/w9JX7AEHFPQoRF6YIbk
iMdcicxA71gMo++p7CEIbBPqXI5zVjozCjH4dyOMtfPxbAp04Yc4XJyqZ4Kbb+zVhlpyAWGy3HLf
NxBt8W4+C5a1OI50UlrUf2F/3gIyCYsGfy9R82BWW34DzUONU9EcCi5VildlVmirw5ZMp1Z6DD+r
Z7qYrsdt4OMqnJ5vcw2KqQTQaLy6TLkfndNjs5VfiyW27jOSukSlvGmGcs1rbXNl2DLuTdanEAbb
tVwwdifzKJZ9WJJe6mzTyJDZ9ThC0TZjlRjIT5/juAaL9MzW9IYK9uB/2OPY0d1y8lRexjEcOjcj
xlE+jg/vyx41Kqx+7JRow3ZxsCsEL6JvgBLc2OazgEYtYZExx/8EbW4+SHie3CaftGiFrkRh31UN
3/PPgzcM6jhfR6aEFz3dDIM+HnYesbUTEeKSHoiNZhs3p8NW6Bu/H1h2R+6sVgKpw3Xl8urUxM5G
yU2DOLQQGv7gnVvh61qF8rfqgodMtTL6FLiyC/oz7BuU+qzWwQunr6j6NN+HcPspUbsKdIQhwi9+
7AdNzD1hr66wZiRzgPSAgLArGU1W675g3ipqoqYV7nD1lj4R+2KmmO3hiw7vMu8RM3zSwvPBZTJ7
x4vyWM6lKjPiZbbfa6qbfWCldIPMxJptjzzpmptAgKj2pi6Ii54a9K2STvy7QBKlrP9eJDJfeVyN
AMIjZSB3D0/pu2JWpYGXFGRvivf1auaI/imRndpjrPOumZlrf+1vjL/bSz2hFt95gHsAAOk0LOj6
B+0PHW/Hzx/6vYoaaxZNAFKUkaszQQNZrMoSAlHF/9zRyDqxqHWn1iRMm4LogspEH9tiTFTyMg3p
h6y28y02p6r/ZprLN1XM16GIZ9lv00TWh1F/xO1VfzFztmgx+Ub7UOfeJtqxbC+IX+gMKjuawHNz
hp7019JGWMoM850jcfzOTxZPc5f0urEVB0WwhjSl7Qt/kJM7IdGV9wC0PBDGQr3WTQigGQH6jnuw
75kPkSqfk7yMkboBggCnPwBEJbWtHGSiSojw379nJkIapf/Qe5dqS99GOlLSZcHrwOExKYeKi1Kd
fS53PNIJlOgf4ytEBIgOaMtiI57ZTc1114f3bYwMvafFgF/m9pZlPvWzUtZLvrZnW5tcuW3u+R9s
jYVpeJJDrwhC6yj2m+RwCtKmbqh7smhayaar9vQHq+IAKxoS3YxITDrcz9re87GSR9Cwv9jKZR8+
S98Fj2a7d6k6SNLN+WPrFv/tyQvJ8DeA+s2GwTMK6RY34MhTZcK8ZSQyHMg04XevBZc8xgbAz3JR
r+wrTy8JGiEowDoIcusW3y+sfGMmydS25D/KMdCuIWMHTnRiGBAVLfjaXFBex/glaS93IDCa5PUU
7DO2xBTFXRj1zfDJ9Yb6KBlRxUF7ute99oZ0uCufkMWxyJ0wy0xIoVsyq/tXLcEXn+lBaDea71M3
DfSkmoXT1C8nmU7EOIQXr0iM3l6G5KcZ4409jKVMMNPpKInrcaZTJ8POwaKJLzAv1Z/jtROnMEXG
5H4RbtA042raLc2GDWwdDTBzLKitnBzeeN/225jDekbJS5trQPnga2/PpRtfWl2wXwZltrL/ubf3
K5BGE9apyyAtYvRDwmaSzLBS9MSwDhJlyOukN07vB05N/gesS+TKD3mG14g594qK2pMAUvbtny82
Yj/BickXBFOOPZ1Bwqqd6bwvPNyIsuqEiWSTrJZ7jcAcGo+SPsf2X9mLjqM6R95TGuTsdYNeBYdK
tbeMZ/iT5blLo4TtTpP9QDnAlzkVvN6EpKrJ19pYBc1l+xBwWTOXsMD7VLM3NS/yRn68kh0FK/4/
1iz6/ho0ukAwBL23ieM0aK7chK0q9k+ZQjSgbPz3sk2LyXNhLM2j7jUZgc3QkS0smzRxGqpWhugx
a7l1AwLWC7XwpLepFlgEBwE6zmtxnV/EGiy02ehLyR7ZLbJl3LoXOIXS6JzVTK44qBeR2xeUTiym
JpFIzJrv0yFpkFliqXloQzDBru8IIRLcAtzF2sllMPcl2RSRYmuysJtn+Miro/QQ/DW4kxKIO7CW
K8+jQkelQYve9hoMKg+VoEWBDqS3sxLvYRS+tuR3k51ACP5lfp961a3H8lQ76K/gh+hDhyl97LB4
/vsMjlVNPbVmDwlNlu/QnhYTtqDVQj8xuaGJ4cX8oWFlFjBD7oahvRtGOHhpW+1nUWPCpfMPRojt
O9liMyREDuGd9pf+w2cCQuSLTCWiX3CV65UIUmj53/AGSeANaZnvKMJl8wNHpQcEdIwmVvnZS5TE
ZcNt4ejXJV6ys4O1JDFYKzCClrDuT3uRuDvgXUh5KgGFjsO0NFvflnSC9Ht8EFQ5VgDNcZmez8Co
hBbbXoxQ35FM4drqVJlnmwkGehde4gbJsuZh3f/Mk7jUuOHmgdHYjQNQKi0JlgccqCTHpwWeIhuR
essQOAyqbOZg+PUos6C6GAtYViLxg9LgHfVAjcp9hDQTv+5GQGP5sNilgfybGQv0Tigunxy+JAVu
WqgeChIkzT38UAK9xbJpF6iIhLdqP/ZIRD3uWlBhNpzf72W7rRtKl8w8itxI1V7DSY3Rxy7r0UPU
wbcqQ/xa4FWGFRcsaOpa5ahYs3dXgCxTUUMwrgk23sgRNZ0zkMVCSIp1zTjjQgdZ7hKeUK4wJ1HX
lK126c4p5c4mlB4/GblpJZMfXBIa+bcCmlaEWoXyai7gb35hyMff3MqfltzhtbZdZQ3RErYzL8xX
R+rsbQVkzMzuauRi59aUIJP8z76vwcRh7Xx6AeaSsgLWxGeC4dZJDK7mlDtQkl+FJ8pTXeK8ZuBu
RvHkCwhuaqFxqD6+i4JJIa23Cqq7ORH+r+rIZT2Vs8KtT6mfWTVmQRaj32yQ5UCS2rWvZZaru7Bi
/ltiau5EYmLNIgklVJieJ+Z4/BHZhP94vjwEvVl/Wxux+T6LPPnjFqEOoXGls1r5wZw7pfI64k+M
cA6T/P+jAuPrkjjHFUj2CpYQclbCR5TrMql3ThuzYpFSyzj1dQbQWaE6VozLeieteBvV7p8WvLCf
cg41x1uiBXKUHwqbr4dCITerFNt12a6DEZkfHVbPktKke06x6Kr6Y+Fzq1H3w/vQO/nTmpYKODiO
HFyj1PL2sNrY0eScu2wVkC1U15D70DI3wV8eVhIcXoyjK/7maKgU5v8HG2jOCbSgY4G1YhEAWpdq
8jeIS+jKrGbXtMNX5nXH93M8H8xOdWLYBGxjrUDZmhbJ+SBqarHT0M9kdpYcFmOJs5BjGKNBiF43
ztID9iyBp/F2LU1FOIkBKwwPlkWGIGkC7wA0l9Ns1SNtS0UxbKffp3Yz1i3Fg0TR9abzgJ3hxH30
SicQhl7h6AqZk70UBUGOKJw7Hpyf8GXj1uABufO1lmSilWu1rf20t1wNDdbKconwsn2wMTyozt7X
bxcPe6QAdh8tClty/5U86yt0f3dh3GJFFhunHh2jDntSRSLdYsT12lpZGdKxQKfPVHmTclr46JQW
avz1/worfUQEIOVCPmUxpJX5im+fEan3mDlGZAVH1ibmZVWL1QGb9LX8cNDE4JS6j8ml2PDlQcrw
7KShZyCkKUaJnrIFZnWEQuNmzQ7U1xECf5TFJavrnsyVyp8xXC46+r7VulhP2LAvxcySRVNp1yPk
M2R+GoZfadJPyfv9ETKxwAZW80LPEIzPdLK4ZzDR5ImOmSwh+hcUbmkglvR4OjB5ZI81Sqji1s+n
5kBYSCGQNi63HqzrJJQGOZJG49UJ8X5pkza2AZOBccII5vtrZCE+BkiEMfJvA87pq1Z0Bw2gwsiF
YaJg4iw97aGHlwpXOZP3qEzsJzrPnLkdekr65vtmDa0SL830AC/YYdg97bx6TmkKFOepkbDh5Fi/
qbhGYTvSOzDBOg+HywqAWTqeGEU4rIKxAdCtVMvjE1BIEBPAHEluXmV7/j5MZR8JJy/swlg0hVF/
TuMq4jbUFCX4KET9GMQ7sHOPisWsJeEuL6VVNNBTH2oC6pocKe5siMYPIcJEZYmCU7P9aambDPVP
vQhFdXfV7CDEGAUxw7CKiSrj0Tc3NBm0ELTD1/4hA4QzFtTuOIepKF/PiIxuT9ivC2++3UgC+/Wa
f2fSIVuhE7HWE0V4EpAi+fXrzmQCeIBW0BWoWZEDededEM/d+SBOZPRsxGzuRs//iHykyz+tsOLV
CZHS7YyRJY0TFA3J3a3oFbCcV6QED28LJHatK8YmqJEldOdnSg3E5QVUpLbGUwyOkuONi4z5QcRG
5qBdEYic2A/zJWpBaoc0QXERxdVuAZhUvcpmtMsLwXh1TzJ7yoVpzhODjnQ7Ly6RA4rKFusZhllM
DdPHS5e1xfQs6If1LHIcoL2EnQjn5kHtNaPZoA88/kdaG95qvQ+nkleZkOHrG+CMzlUcOaKxWnHH
zo9qYhv4w40eDYakX1t3D3whNSwQpkoCllaoJH1XvB27/rlIXI7QY68R8+Eo0XrJIsMOylZa/ZOU
rQdkXqvWqCGjVmY0xsnz4aaid7Lf8hOyPxVOZsljxOCNmmx5ZmH3ppqtDVZ7jHCg5Kf2AAuB4H5E
i2h1fiYO50GgtuvVJSuYeX9Et4QmpsWmROIUNK8pZ5gklHbXlIF4NbpyyrkgvW9juppwGigVuuNd
Ky4jIJbdIFeEn2hAnRKA7ooiS+XMjJ5Ck9zjMF7QGyznfhb3RP2LNY8onswx4yMfCRjYjBIpXojy
pxh01ZsbmeueNp8Yc1eCgVtA8DFuJCFK+i9pfGtUw1srVzint1uZW7mgJKCUKsPW0uytSP7V+/2n
1GcQGPjNrcjFsW0O4Hf/+ZLv2eGMpy1gp8FUVlc9pjUDGlXrAsvfcdTZiX1i3ySoPYniN8YgKYd2
QjkIP+DuhFDJMQ0UwB5Wpx6zab/YPViKm28igu7kWgxe6Rj28/Fv9mhcMVLg4uL0pDR66y7od4DD
GaUJf/DPGTaXkC0XHsyhp8K5/1B04fj52M7+zILFBT5a17fOt4AwGubDI+Ph+6RALtjN7560zzz6
i9St98ssfn+1sDGkLoB3H1Iopl0nJADgZPV6SJkQoKJ1aByrB7bv/k1vieg7tzuP/4RJBkCABil7
tefTzu95fe2ATBiLMuc1Rd+nXBKgTHm4ntFbOZwUN79CgROkPxrs5EVa3JUMnaRGNM85VsW38OdS
SHKJa0tGaioBN6BhD8TkBbphhqeS8oGK2jR/gYVCnQkpGl2VDbq2mqpQGYUWdKFFXWuXMbavP5mv
OpC3ZF5l+DTy8+Jj5bpnMp7rLgoJ3KW+cV+3tKMGaic0CjjqK7Z2COy7DSoT2HmleJxU6kC2/gT0
Kfkv6bXsO5G0p7X6GXTqmEtMD+x6gAJBfON+lF7cw6ewO+ZBUNdbZotCLXxJIPDfCncR+S1U8Bof
vbrNDaetrD7aRkuuxlGoV36Z+0mVpHz9RfFT+8dBKycELreFILt8EIlsZ9HzQpvKZBavo8YQ/ETh
1KdDl2rmBgRLW+joQz/jI4CFqzmylWGGfqUgqp1uhjWuAq+vC9Kc6zJQGdzCTVNgjUJZBALKrbAV
Jv7eqKPqGaJZfRNbiwr0hccdubgTlGXZm3k6qViueFfFeBiZwkWkUcoQck9Z78fgELurnCAR9v0h
17Cw/U10ojaAKHDp+Ru7lbBsEsJKD9gymHUlo9eCHB+y5OyeQas14DH7lkNkPJWLaiQGlliOcQD/
zKIRbj/UaJ9vAPjp9U5FoCQU5PpdY4df47ZRiisHBfEJce0HRq710ZtNDBNneRg390mWpzftVz9+
1OOG0/4uCat0YmVUC0ulmYJHpAFBjAqzinIlzB4DiXIBrklLJ+339kHpT9lIPlsRJVOsvT6VtL03
hBuZCP+Ma7ujcAvI3CA0k0Kb3HNbgk85dKGa6TYdr46UXDgi7grbcE86yjEAm+I3s/YyC6J0WAio
V/lApYhJwiVYkt2FLsrjkDPTqwnnF/ZCyZCBP98WyCoR6SwHxo8ET1iIDVpkjh0SXdTN3akxC9qM
eMgYlV5bMExE1EkV/kaGARMWTa8dzsjIcXML9N/ojyeg3FqqS/UPeR2kBVKP2yyWTA5QHjWBHB0i
G47eMfZ1RaqduudfaVOOkCk4agG3JGOOUBLP+VN1FWUIL4Grxi/iQorSS7DuKzX5LMBjJEQqBVmE
dhFkJ/4Ks3C9HJvYWzVdsCmltveHNr2MK7/2Xerr7ghq/V6QxliKN1kkQSvNg7h4ZJb7aJYB+5jb
yu4dV4SbQbG9oMPZx9aKV8RzHIETyNYGjhAdhx+7YhicjDRNOm5ngA5O9ajqCay1fKsU0Skt+6yF
jH77j4O3VwQ/YHQoTJU+sE92vkM5Jh1E5hvcwc4NXtQxwJpm3HPz7DAYTG9ZmX8Y1gLxx8XnWpb8
TnmrFp49dppA5VILczwGxYBEqlPhjWcolWzLbR8U4zVM2DhJNu/ZFJfnnAN8PmGMY2HnLYxr6hHm
IdrnZ4MEo7n+YVQjM7kRFcI6EGTQH5Ew+7KkhrerWy6hLRxNVx3QRn8XIm2RXBORRu6u/u6omwrx
YYFhYl2ViGdqEeHNGZcvK9C9d6xkJqLB6PhoOEvbyb4pt/jwHMhuGKzXXYqtV7ZgbrvMfTDKy2Il
oTxodKi+x+gS8V4GRQj9aXs1zdSwuKddcWDdTq4eBpNCZO3XKy7WcW/x8RE1/78WMJ4xESWD1lyk
zzaQU4ywAJSCpZDKTqeho6/6QzfFH8V0LVIjC0z12b3R5vYYYHYCtupAzLgPRipZ714ZCulTTQ90
8k707af9EDILDF+3cdWs51D/1IlkGKmjLTpWEjYWek5wmo+UwHjeMU6t8zmGsoweA3CQcCJAeipy
tndAANPx3Y4AIlbGa30E5cX/G8ix5GIkdI9wwkp5JNnapAjYD3tvbhTNMEOEhpfhoQgQ9LI5gWuu
RvpzR+u2OPSifq9RCUTS3QcG6KG7Uyt4Egu+e0cHAsXwW7kil3+Iua8mXLgzRvEB6T3SdJM94mxT
n4KJSEVJ4br3X+Qa7KxBx1HIXfM5uiNsfvLOJu9pRw8WvBm3QrXr4TGExEGdemdGaZoBPkEHCy3S
iF1Og0FSJkeRlBtTlZKKsDTyTqlWHP6U/59yjOBb6kQWbzvfP/e0/CWbrftLQ7f7lliC5wZGpVLf
D9irAZDiPI59bE2dbYvizXAurogysGCToSXO7o2yG2TnkYvXMnmA0AcjJis1hMcvlD7OoFWr1e2m
SOUZtUQfcNg6+h/h4ca8ZjcmSBwnPLrhGnuSSfd4zS/CmKj3MHB6TJRAa5VUYWr8ONzM5hAOmXqN
4a23VlWVYbkN6TsCCmL4o+a6ph7zX5w/8Lg81B64hEdlMTmhtf8hS5MnifOKHV2gvx/o4EkvnidB
Qio9ugMCqd1yMP42y2JKT0xC/NQASzoBECTxMm1QjsdYuT6aXxa1Ze7ibYMMAFfHNnWtA+Z8Dphm
bZIGI2iqbdfBWEHFgrIDssU5xibluxaxICTSsDP9KKrzd4OpXXO+3smikUk1GJatZRocQEtMT6vD
GA1yEisT5zvwKki7Uf7ItjZ+FurBmDPAbc2ZTfQL7a8WfF5zwEzl6P8OhBxMlFaTyi8evA6lMaO9
Zd7oE1+SaSR0OsQ7474E4VEjkkLQ1sQHQK76UrU3x9jpMNOi/9wHF+D7oJ2X9fZGgpvjsdiWlfQ5
FAfCsUdCf+cBlmDhrqGkEhbTnPE/en8Q9AbDlKXJRkpDutTXQUfQksf1cJ8t0ZvOErpb7d/3V3z3
73TwmFaas+Xl3PEs6ZtPxjd62in2SVXFr8CCD9PSgqMK1LU37EMEm744usRD9UlyaPVA35q1euwC
L6Vm3O6jnuX4x4N2MRrCxiOTIZgNB4xVvexx2e3k8G/2s/BNA6HvXgLCB+kNhtpRn5aawhy6z2/r
oGoYnDZz3UfYqmvpBgUVAl7e9Sjn63M5eggW5TxgqvPazlbd/Ez6jW1E+niWooS6auLgOAsJdcnQ
HyYBYwKPA4unOGE5eZeuk7pzyipeiH19JkqpqW+dOd/AVzROC1BYS4Ug3WyOP0wgsp/HDzAvPPVb
hsgUljF7fTTzbKGro4yt5eFvbKNCCh+XCJIBBaqsVrd2zaO4XmSGiZ3wuEcK5LSx9+8k/2sK422+
N6U1trksW0GWV3UpIrc+KV5HhEdU7UjcTRrJiubsFw4jvgEQlsJrDe6YZCMsvon3rzqTC0AvsNzk
fOVKaOdYfaH4K7Kn7kbRvBV50hkdz5nhvQXgkxXddhfRFEs4M8cV4nzN0hUfhhM9rMsDm2W8C1HX
hg5MpeGVzaO0r4h3uLrUsySPk1Jud4KT4L6g0erxGoQXoW2E/uKTOeyyzKZlrlkV60K8/3zKQzWk
lt4hwPNglZ+LC+sN84YNTRbO0nS7pIQUMLPRKsjFF0kvYdpg+1rYEHbb2fi2BwF9kBSpZIBmSstP
eJuWrRDLfKVCGNJ4wh7jsE43+vKJZZOIR9CACNaYm5i/wXUVd+n239FqRd6CVck1NiwCT2YyZ7af
jMhkhZZaisU3cP42SM4hU+O9OFmRewIZAi4paYxxhDxKF92Ak9Nx30fwrhtfP7Ay2ZCIzzf+WTxF
TmzU+cpD504QaBtLzdUuPjJEMY9dqSw80O/JZzpdC5b1WcPyFBF4Rr3YMucxcY/SG/MAlRKTerw8
m2/wQq+dWX8Ml5d3CTK/y0QskckT6OcgjrB5VrH21SxtIlWAPFoh9fC5wTwpPKPctQQQjArrJGRi
G5xD/PwzmRshMX01iHTs/DImIwNCYmAuFwISAuJX7A25vS2sWtQfn8HrJtL1T1UJpfLEuLo2hXQc
2aPMNrJ0xc64l7MEn+fEur+awXokDIiPgelDltlbwscK3RSrEbtSSw9uTGnc7nZKaoXMsKXkHTBA
eprGkDIa7iyTFst3gUP7mUv5sTrtKgo72UlELSsR6Y2QEvu4u7sGNS+W4TZWiAzOzHC86jdELkJ3
XFXfy9x/BmuTqlWjQYtmZr4YFWUp0f0zypxyQCPN0Sb2EwBQxpi8qgQWgCtGQP7o+8qZ7LQClMgo
I4stXXmXfZIF5ZE/ia9JmhaCISAJyJqOxywaZOEMkdK0OXZKiDH5Ssc/yyculPuDRDrFA5MwJBKM
N6IFOYRBysizf1mjnV3kTQnNMNkyJkYSbLfPE01Vp2uvilSkYgwzNiw7stbeAfOcYpEdfnF6xFJA
NsRCGCtC3b2aAIyjSlxnCmjtLI2SEl8HS5T/FPr2lTqw6sgfcpWOOS2yAWfpAeddTcOXF5QLHJZn
V1wA7GPu3hqSKxi1CF339l0Yz9dlrroVwlvNR2ChmrOUgWUBmldiyu+9FAa++GUlN03kZr8dV1ar
jE4swo0W9X+w4xAH6EhLtMpPebsw8r4TaMw+2DxaU0U6z4+ohcyEY9JZMnMzAeiZdqUVre15ydNS
qfDK1Sj5pqDcVfmJPXPVmfZw4m/oPlkimeo31r9WlZ2wy0H9/mwWu0LvtggzDkMvZ6BLNjhiQI4O
G34g26qjRlYlJ5knuqdxynPRYZ39sS4KS99kEbJ1E8JEoQTgS+/N2XnjNukQVXETTFVwtEw1/sJ0
TGd5PkIiqQ9rvrdyQXt8S7o8/xPUk/z88vpLvS4VnqzBmGg9s5vy/LoDqQowfZ6VnJjy7otNd0Je
Gs0DeC4GuRSRJradCTgfkQyaPhonIBxsuA/hUY1a0KRLTiBFcM/UCwIFTAeMRUMA8/uANILbwe3l
dP5YP7Kvl5ql3+D6skGn2fc7Xa6llQWx1Im/+QvJwIpsIEKrz0+46/fp7pvn3RoVJJdN56OlDvoi
SL62PuVj2bPm5e8qGsL1O2qUYhQm6lz1LYiMdWGGbohFtgT6fg+Eo8HnexGvwKsvcGTTuxSGA6Q7
+zMsMYKRb7uW2jrGnGg2z4hSsNDe1w+T1RPEoJMOnPgzNu7mZvtRi4W7ZJYpCRy7BVrwttBLoRfb
Bh2S+Lyb64253Wow5+EFGNBw3QDP8Bt0WnzCO/tc0+HzHd5yA/w2Lrm9dpa8/+uFkGv8grNO7v+G
NwURvn63WUESlaKppgYvuQmppx58j268v11PD73EqGfxTLrbR+OqoDzK6BuirnwdvYhuGxAlr+l2
S/0iSerXqTJeTcwgR+BI381uDh0JtfEnpWwkPeV0ucfaB71s3ZKP21yn8fPAcitEiaLflpZ3YLJD
WHTsH58zqD9IxdHVXeYNrdS0eNST1+87uKOE47vsSlpWLK6Sr0LcXnUdWxKZamMC5+ONWQF++eBn
AzR760yHz9zz5qfhemtFBKGQcugiO9Kxrpo+LUGLAJhhL+6z2YSIBCfgqcN1Qgi8/y35cy0rs7e0
2e/pPjxNPZLvxwSuO3vDEEHuHXlXbzUVrKKKPyOf8tXsSuK1q4QcpUJE+iXefqVyknB7CDGY/aqI
d0cF0wXNKljK1dw0Ptb4KzUUTZWhflvdgrjTzbJoPz1n44/y/B2Bbg9wQiiDPfnlzHkTtZ8Tnt7z
CQeAXaa8uDXd/eO+K/i6yB2+HYC084+2/dr9aQHD7FRmCq+ynTneLvhGFSHO8VKX8hQa7g9HPh92
rnEA2LMQdAv57jjKrHY38SVU030a/ldIPumuWaxaZLXtT0snS9KI8TlPACSjaaWqfX5/lThlcq2e
mRfp5K5KUWo/RpxshsruX9RWDxpC7S5P+05ht0xE6xjHa9RRjRSCO/LiSyXkCDEyln3PpBPPvUi/
TWq+rOEVBYooP5OKcZF0JPyGuEiEfH51N7X7xXgCcydQDzD1UWZqE9pDuDIxOOM+o9yDvcpDhhuo
MkfMzx9Ojbs2r+/xeUQBFnsqAnTFyWK9vEmGDSLvGd8m1+H8C6jXqGDFlr9UzPm+uZYaJcSNzlvm
q+9eLNQ4gTYcnafTMAw+5q89GOPk81bpEaSQYivTHU3GrSkXDng85aGuCrZt1YqfobGGxeXMXJs3
g67AWU+NNuA0OZIvm2SMuXNaYmBs/sgJTEK08ptgXyEMNLCgeVaLCMD1iQyPlIobZCA3K1qa5+DH
D6Zo76PgXVgAD/ZdjcJEsx9MENlWmXV+pFsKIM2TD3TkdinF/VyinFlhTknAXeDd9na7SIOQj5/Q
mILqsiWFz/v52fCyJjkjPscRttEA86iM2VipVWHKQAzdGy/zTwZVYqXji02LM7PGD1nVpGWnzs4O
gJl7wHYbjrGlCP0iBqu83Dacl83oJfemry28L6N7NqmikYuZoumePAxc63AjgJZh+xpNHit+jCNp
fzy5vub52OWEI3jW6fRr1SYTxkDr4yFMzHz/Y9JNTJ1XqnLTO11/Bkmenc0Ha4rP9w/2ALr5zcjp
Cc1TxV8daXUlf/iAPxlf2TlDsX9xdB2w95Ve3NBcgsfjGOzaIOmRJQU91SuCfz2QVrqBLQaAtb0B
gcDZb6C7mrA4EhbSwi6rhyIFJtOf11AVmUbw+HJmdBsqhVys9Va8k7v65ckVcN3VAxtYRDiia05a
+QqXWrk3t1Uj46wPHH0iPqqkxaorhDmGy4BkygkW/+Cl3oroHn5Fy6QW1yCEXHguMmZwRgnMhrDt
qDPEVoCue27CkYw3o6wPTyqgGc0XqJOqZUwOyvp2Wa2iTxS7J+tptWS/cd2rPIgz1aKgybfhxf8c
w9MCRkjEKt/bb5tsQIFqxLQ4etfGQP8DX0ljODO4srs+E28Xn6LCDPAC9O8aTRz1B1SXJlHEIXEV
eahqDI8FbGFdeuvFIfCeyhM6sq0VAxInQaAbBkM64zIcNV2I54ATJ6pwDwORUpT65GX/mr6kGmv8
dZBMB3pexCHUl53nEwZtHoLTKxPeP2YbqrjwyhYmmfZvWEazRzX85T7h9cOSGbhc9/kY4P2LolPA
pa84bF/ThMXC+jfw/nbdKD+R1vdBv/1YpEgXLby9XlqIiCjz/aXLdnay21n7haibwP9iyXrpfOFs
VzbJKn01mhXM6xcC8Se/3VCNKVh++ye7426c4fFeYt0rMlUG9PK+6Z3vjYSXnCpc04BBqxZBJ7KL
I0L6f9B7A1biqtdRIfgPE2XO26HnhXQMlwqV7EAIX9URjT5Dk9t7uSMh+SHbBk2xvt/6FD9OLrQg
EXWHN68WreKKsKAPWeLksrO2lnsPFtJYwe5QsKnLs49AF9zeBVNSirLeJMl/aygEz7Jc+Ep2zi43
o+eq6pW5QtOVD0z6UJpxB2hQErRNM/konh2HLdG90nTutQ4KyOKIMfitOuK/jjq2vL9mHQ9zCXal
yEf9JDB6FvL6f6ojHmZU7U2JPCWCGhMERd13CKAHbOaWctbn5TOI2Wy675wqrJq/3/jOgW3FqGol
iZQATFs+69JERqgGAb7m/8yjKgmwVn/Sx3GiR7E3RxgWGibrU90/eEJdfoayqdJpGi25IAayx5SV
KuUKoeW3ZroMhLTR/6G0+y4cJbt+8/JWbtfLjDrLomTE7EAu33zSiDuAQfvIR1ka9Px+XMR84KQS
tA4vzhAMGTGKWXLYxl9l+AHZ0Dh5i+dO14W8396k0MjpTMfcYBRRSmyL7kCcUqLsw9hrLnrbYgfu
DBPfWsxXi1dpA6q+qSzoGdMXAVyTNZz7xnZZNQJcw6aT0xgtSc1vZ2Ey/JlYG0165d+7SBDTe4lo
jY4DzL/Gav+X51DqitCMpJHZmiMXoDXIqq2gapZxjvSQ+u0s1IvdWM2vnFQFwGIjz2ouMl4ZiI7+
DAxZcIrU/DcSaLXGuuvKsf4IkwYHvI1lbZdN82rXlA5xV3fUMB1hFIjWxQ+k2Ovn2yfO9mqWfZM/
OzM6l/UR5mrsY4a33iO5QDr+uesmLOBwxdm4KQ+rg52pYpMDVcu2FGvmNtftKzN8cBM4LUQTV4Rd
Z2f7XS2MMpwGsqmsqKnY4CWiYzIxWkov0zrys8DoHOnTEtRTICAXKZN91hZGdKc5RgcC0aJNmkIh
SYJ1xJv0Az/BShXlj5rA4p8NiWaZhLTEvnje7TcJjcjDco6yNDl3PMt1Mfm25geKbxBAbwoa3nEu
xKHR8yVcu35gAasWmobCJOvzh/C1Ewi43tnuPL85LDAiX+VZERsuAsAJMoMGUulDB/XpHljeEOLw
UwU8AJ22smc91HN2BONnAnhT1ggLyuCjzxa3SCq/Tw9JybLDk0IsJe1/qGIpYG7jqM+PKUKplayR
ajHfiTgjA12uqnRUERucFSrlL944doAy5EaAaJLgcULFvRaspl01Ib4HcYbJj8xWBSF0S+YZMM+d
/qtm87T6bbmbfCQGfVGIX0yWcNLIH+i21nBTGaTqaNRdjn+O6OAj7p9Ne23aZ1flbETGR6AKyZU/
1kJqcfAsHodHmMETJ7s+pDv4cDHNUd8LvIa4p1e95GpTEojeCwqIlgD+Cp5RkuA9QoyVnK3xEKGl
9sU+45J/th/7ChxLLaYmogI1+ilduoY8Sev3EOuFqPfrDbMWu4vryZIE6pwScoClohrvC4Wg7y2Y
8kzdqcW1QCajIfGpirWdMtv69nrze0DX4UtaLDiQBmiI0GsO739Qley7reUI4thlHpOcdenjlJ9b
sxkd0S4wsUs++xa+NCahi9GcyyA6EJNSM5dwEEbB+aAaQpudsxWoUj93F5OLAltr+4pPFcnFNZpC
m3KUQE9wyUYDUQkNvMJGU+iVnIFHRg0YpG+HUYV1Fx8g4CmlzDqexE0rrRgCGo0UZ73Zj9gxc7T4
0/8CXJQLw9qm/52eJseJXMn9QoVF7AjBx0rQriGBf/FQVNtWBGz9EW+rQavBSXK3yulWUEEMLF43
362DU+lwppTnsik0Pgu3YPKnNvnAcNuQEVGk9Sy+fzgOXqKBf3g8d4tmfddo/gMTyTIMQeLxH9jO
nIKGpOMN/TMo7GHyrkHqh6AJO7L/pD45CZxbM2WxzC1sM1OUsUqL7VtPqQjjU/cEP5THJ/Hc1SdT
hhlPo5C5WBDUCXlUsgZDkf4RqSe/xQykh8BBYS5/EyVvk+O+dBzH5co9dZtdAKkEN1lV85Ok1a7E
z9FceKPZXHFaM95Xx4mJQWL/hzhfgoD7kiPz/A3/SLVcTEF/9kydh6LohP6udHjflomyodOma91L
bRUKH9hrT7sLBD9plJilE9ojm4KE/xYsGXDbyTg5XzkywKzDBfZVhP1xGdlcYZDUQghyIvVSgkmC
FEaYUDwQk0sPm7jQacglxAubheYjZCuPB+NDjMNHnWuS5oqCoD5bUc9ulUo8FBMNfGmXQqsBUSNR
3OWg4aanp6H2+Nxu0xwsHr6quJtRQueWs6EkRDhDLPT3Gebw/aFeDifQxl1c3Lth9yg92l5obEv2
tf5iWZqw0v2GESDi11VyY2u5NtrgjtMFoTbvkkge91nGINurvtsqmE+RMeCNYVThLSTWOk3O+BiW
4qdkpq8wCUelRlyMXF7dFjhBs8HHWQMrG9wYZ4s3qteMH92FdkRlvyCyIYJkUV2fqRWyKjNQByAn
Uhhs20atIfyuDo8iERd9mBQZlODEMhCMjhaTU4H1tcGpLhvYjiUESYfL1IaPXPK2i274zD2AyL8R
ULBvlvorsswAZuB617mFYSwfP8KocUIVv0TjL2RZmZmYmHwSk9CX271hUlFqkrIU/hp3lH8zrT9G
4dTM8kXGY/4ZskauV9idgbl2QS2hRzRQ+lLCtM0klRdDCrhWT+5Ev3zSrolCrhoMS3fEmeXwLqux
HEYtsdPG1J8+H/79jM25gpChEPJyPsnfgnbYiVtby2BLf3zAfDDf2WUtEO4B/5rDqSZYKEFH82CJ
o7couoS6KjIn6dy3iPOmerqqCS5u08U9yGVD2kTbwmwA+jA0t6oMNzgjyhrMdWwAjNLCPADNyVfk
eWnqd73vn2lRHlc9BFDIKqsVy1k4Lcerq1anmizZODcCtu2HQTq+1B+B+tZdfJQ6wuCb+SoDyd3v
Z/BTGbs3prO1G7Dos1chrGBcVWrMvTJUyEcaQF+McTnpNXmvXB6zMn+x/YLE3RI4pBTARBatLE8c
RzfIhobRzKZkRDEALx8C1SFbEXoPHA4r8G2nhUTgTYAwm2vNd9FskMI+ftKKDILJceKNDGhHGJB0
cwRxV23JLL326gOTdHK88IMcbdG/YKUSaUZbqw0EhXydb2wJetjjuVxf4L8BkjJ5MqoaTHTy4V9E
N3wc/+BvCASnvXTp6lZoQzvarlSwLdKYcu6GtmYaCCVrE4tvxfpBnnifPu16+jLcn2l2FCg3BqMa
VOZKKm+XPpc/kME3s6zP7ucVs1xpYnyhzAubgYdzIBqNLFTVRBhXOPGstUli7Cgh2riN3/zug0AT
qLS8xd7+dtxQxh1vkhl7FcBB7v0NlK/RLxDS4FcgAnhZRzkdJKGXNds6Gz4jZyhjAQ7z6otLwJ0U
WJ2bTnPIcNHCgjWuFVy/Ga3U6rJHGoKcRNb9eCDVwIoF8q4Gf77VqFJaY4Bl3Jilk+JkUx2FfHr8
qVGJQ3iRKaSu3rMBHgpx7/OVP1KYdjx7m31GfD/BOY2KggMXILMQl1Vjy85TLggCco6TTGELo0R2
JwM35n0qaHVLF6Vi8Bm9c8NSWnp/3rLQk3RA1lHaDjKODXXMkpJ4LotoEfPE9yF5YZXPJtBDXDKT
zkIxaAK1+GChT9ZC6gHdsQ9Svi6kKNGaxb5X37AT2m8yt6AeKDV4p4CqvXL4c4LLKV3bKgsvgVbD
CY+1TgIwxm9GP/Lyl9RjMMNSYpboc52g8qnOt/pe5lfeOXMKcU+YuwjD6Ljrb4htfpozbQF/fucq
z0aaCwvylJwz9Jsp1DBSZiytiNZ6PjD2BqM0dWFCEws/LKRTHnXsaHOx74r/Q6IrLwgp80ziIjXy
UaIT9xCmRJNziaCEYSmEYnEn6jRLxXWKSoylCiURepVPm+5UvzR4/EyVvrSybIG+j9zhJu8UsjKR
MyQcU23Z0xFc2/MXdVGAjBMAWnYRsthzpOiOndCEd6CG+/8yod3BNN4iECe4zF8y1/0y7Zm2rg81
IVhJVG/jYaz1wW6C+9113d+1J1XQPD7oS2/0tLi0tVHNnB9cjfRyPSu67eyl8038IbqE39PUuQHq
B/xRV3P2tEcrFVafDnQd9ZOshd8g6cuo2IX7lO5QVlYbqPnp705Vy/HdTaNSYk/WNG3m+0ZWnCmY
EvX3yZiJd2s6FEa3MbN8T1b1T98ajGh94iyjb0kzW3LFgB5IUjMftEiMiH/KRaUV8Tc9na/kcxeI
sZaCbzho1k3SfXvpvrVlo9PY4KY6y+1OeMBTDn3OrvR83bZ3lCsR7xFCA+GZtRigkaLjgs2IVsrC
lBM/hx7chz0qGDeuUlBz34hV4dy+zfIVLTnz+AvrStBGxIPVkznYidvQydFDd3D0UOg2xrBb0LW0
elFVxvcVgUSCawygQDvWGrOJuV9m+nWhRDJ7LXPhvpbXiQt50ePEN0g4j/HyBjs3b7IGfjyP1rOf
wblYBKGOp+gOiEcPsmndiOPRlGucNPvzxLVeS1b8A0wDL4L2+I9GOLQWW/g3p0Aw1nflL4BZ98ZZ
sbtTnAzyLMYSxv1Ncjpy9257+9WGUBbIEL5+g0Pkb2aetFYM95g7L5+cAOx3Gz2sXUfkFptxCtBY
TQgXlNT8QeEJ+U73eSyPlC/UGQXEifAOPA8exSDSRv+kQKsJke3YPCALYUy+w/AZi9es+9cz0Ia0
HlRQ39AVn4a6pjCJOnma4qsUsi/k/pO8B+qPn4ZF+8yncIj9Q2WYxsUvaQnPTVcSyyVikTa8sWfl
Kh8cz9obb0mgbgGXv3LoHFQtlb/GlsPrlUzIw9DqWTh6Fj0SsZ5S87cXFNJCYIi0G4r+DE/1v65F
NDkr7Rbo/YiRqqRMxXNcz5PHjQLZ9O4UkwKBuv57eE0VSLs12W5WzSCAN8u1tkkXm7uR6t0L9MSv
ciYrayztTjNx2V/ATcINBgl/yykTCrixEdchexjzsJNtZdnMsut9oSbHYPLCz5M0ixp1UANPeEQ/
0qZ++1+Z92pWoOfCPNcULlYRT6aiFWqwWW0i80pGH81pssCj7c/8cD+4WPklfSSoHEQi6FaDQ0Z5
imbnUI4C33otKJUbZZ2BdjesXTRRkipk4s7bf007gHxXmCnrjXaMsZVeaUA3+X6BnQX7+IkyWyjc
IuGIR0aM8bIsprYuEcD6d2z0eNUPsDPu3iaTo2w8MDYEZbGcR1QoyRF44yeGrq4M2lZAoXATrUkh
h1U/OYzsmRIde0mZ6ve0CiN6xnmcfn78t3MDmR27GY6NvzQW3NhMYGtnlbPRUkKc26YMSuT4mqT0
XIg/zRDAAu0rYWgKdx3iBYq44/6gkg1Fx3c/J/2Rhh+Ht8Md+ywfaYM/YEKxfMxcUzRLbfLpqfqf
uOo909LJnUv1XBzyYqU9b1dTp2F68M4kR0bWHN78hY3xHM/IOJg7Y74p5Cma2UN9YCshHqO6nflV
PSXvF7iIqiU9eAOEH48aeOfzYJUSFIJOtMKYVShoYe8M8x+KyyOp4CIGbhaE8LJ+AkgQDx2FA88T
n9KC6SQMAbsZ9Uq3jept1U4G5tjSyQmLnZqGoXgDY9TaUbfz42cL5wFDgvDxikewV/UsNSzrHFEz
fkT9hU7Vs2fzDKupM1D7gx5oOZ8LacQgXqWKWjUouJtjWnJu/Z6uxdSF87FLZjL6S0AUueEmq3Bp
r45yzrZhnY0mehwGn5kwU0FXeO7lj+nFCaymf3ttzHBbtgKH5AcFiwoEOuy7WIBx3if7emiyU4rF
PZXEw/gKmACYUItvaiK9yMLAOxkOrpv7PhCL737VM6lL3vaZv9HZOXceSsMOZQKYewAQosJpedz8
u7ytAHnCdp4+f3sBYnWs3jPJtDSnB+3a14csbeYWu6bFDkhHk2BH1mgjvVExnXIA82Gk7aNtC7ag
JAv8Taa2AxXnkurmE9Egnwj8ysoiG68jHMowmTd+oZbiahWnX2f3c1YxVfhjrsXLYce94i6g9oYL
l8euBw2ISPOva+WrAK6mOH8GIM+66By1dstLMqG+8J6sIMJcSWbrIITH3SDR0IJs7zSbVzIQMbTL
3R3WMsUR+YPJuu/UPqN0dmyVct02qIkoQz9mYTvB0FBB9fvL93P/GSkCVWbr3fYgjS7T29hA4HrP
ReASh7uyePXrHlLU8i4w8mQ4oZGwX9cY7eWiic+4qM2z83cneIXSBvEEK52OjiIeGycIez0jIF/a
XU/e4Lteq1xu8yjkmsgQEYgVz6g0vf3wqQXE69IuqGqa4EeoxqaWrWSmQwi0lmu/T7/X2YBT6pmL
Dg5//A3onJRH+4OoBIeIhfozaXzgZDcYBFi+zTJu2iFdidrIjLeltKwkEPzmAR0hpvnc4VnLwnq7
37tsLXdFoRo3baVZFgdOmzOQZcovtvEUfNX017MNjUiMcGATRnL/J+lyZaOHMfaxY4eviUVLOmwo
vm5eaB1SNY1cbP+iS8Do/jOl0ngdas3vsopRkwpBqxpBLbXGfrSe3Lc9ZnhQyzEqazdVvqyvyUwI
OjeGawK3jQRry2DOVGkIshaiEsXC1GriaHbd2iAMfvLL1VtU6j1uI2BvcVW8OHQfEC8Qvn1HA6uJ
N8GF7AqKEJUPGjsiPP1H0W9+bBLtSIxDSqDGOEbh02t2atoCjN+XdfloY0Br7+Pmql7LQcnxqZ7Q
vBLtApcZaLSircArKdLLYBXcIkhu7WxT5kav5xNSAh2e4E2jL68vEKGIfxjKpbDwDPxZCce1XqjE
mU0XyBxkaCgVePv3aqh438UNvvWsT3gzYoHj/bVaoHss4ievEFrfIYw4+H2n7NsBxXJcypaElFJJ
BHmAfSDR32JQ36pGAK0LHzSKFDbxK07855uIfr39IE5MDNB1zTU43ejfwkDas2tCryMRJFIiPh+k
LwuMMdO0kFa9H4EsPW+De9VQV5rke/Kl9nwwuVsbpPHYrofjNJgXOoxd9W5vw2jjEUeG1S3x+Sqb
tLDO6QwYWDQSKy6ithEn+GKSRnWlsHxrgLqXNyBB54e6rlZkN4tNQxdosQ0r3vcrHjxYZLNmBN6M
epKM0WNX77rgKS8HjGYNpcBwrLp8/VN+v4fyxmKyz6i38UVlfX94MhifRcHwAeq91Eka9+eizEVn
sQLG61qClIwyU4FEYZ+e1jFBg47o0PTDtEfPzbCyKF10qz508YMdX7ziff7cDMOH956P6zYKkJJl
D1MAtqsf1Idh2a/Y7SiSy4/WkvcuNkmmGr77YTiGgkhVEJJQ3UF2rkRfRrjHHqNRL9GnSo4hrEr+
ocY+UpvvkoEcb+OYq5DDdb9wtIOVZmbL4GxtP4vYh8U0NSP3/jGPp4mRO10CZToTeyN7/uAlLcll
V7Rr11JCHArMBG3s63yNztJgMKFBdUy0QvUxDu+inDYaj50+RTA1slrFIrAtFWnj9CCYMTtZZD4G
fWtZJNtY3QhPZbEyuDOvX987e7YJmR98KQYRzJZeCQ3/GcP3zmIh465Jqbf8ktMYzyUWlCgYMuuC
kGUu1o61K/xleEsZLrhbl0e+y02noHkzd2wux0R8MBYbn7cQMdxv+QtLrRdz9R09e/NKGVf0bYPa
91AOGAkbTN5Idewk+94j4cUfaZvAcuYDrWQpg+RoZ01pv83EJ+WeGNSQ2ZyTN5VHE8WZEuSSR14n
90YSgl0+sr5mQp93W1w313Hi9HwoNoNymtWeweOEMRIwgK1DNu7DmY5R4BslVUSHGUBnFQr1kmXe
UTIT/nRNM1orjsigcECXOhSq9ZpYogwxQBsLE5MsSaR1pIGtoV8GYH6M1xiH4JU9E+fudhEYeY0j
pBaOhXflgAbooK9HPS8KVZaNPkbhjHGRgIkJhEyZoMZ9xeIUFkHFNsAygCPK7Sza2Sm0DuIkll2c
eiB0C9WMrPSpwpl0s4aPn1PTHhrb7w525/JE/Sj+Xxp+9PCRvNaHsAM4dIsnEk55q0HnfOUqLiys
sn0xWd0iFJNiyoeIfAxyPP9+ulMW627VssLzoSXowX6/jRFXXeNojcc0ZXw1QBJJwFV2Uyujxa1I
6bt664xmbV3S9fzHSc6oXxRlfpyEpZ/oVSjD25tatsw3i6fGyZrvqTxluqknwBfuuujB3BTNm5N2
0C15KMZdf/PnDnMkXpXUVIMDPF29PxPeAz8pfug16D1LCM2AvoEcjqO1/nfrRhqVIbwhz0Q8sTNH
td9rgI0184HE3fNvr59Q3OxGgQybt7hliynLUXz7zm1C7xpOEaRPKyf3Ra+bC3Glxe4OAzqc1Kul
dtv1VGHEGg4aahjQOfTAM33v7NoKMNWNLj94E7AOS/KnDmUhdBYRAGxzL7IScQ53ObiBBkNgoLqg
EEPEk2qy6hU7eQN6eTdc/uiAm+ykCaHjNJfy8WYNH7Ba9DhRmVtFcV+oVQXSCU0TZ5tWRpp5ux0U
5h8OdTNVUDg+/WIKtSv7UrV8AE0/fRMUt0kK+XnEG5Ks52/UbotziZGmS0KvzFh7ITUCfUb69inw
8yRGgKxmKDIouytBjGWvFImoDLU3TkZG0D689KOLSodqWpvd2AFMHkI2mh+M9g3P2h+FxuMBR+Kz
EQ+iRf+RZpj2C56IgXc2UtJ+WzZrmDGdSSZ5ZoTlGHP6rniEmFm1isob6wSKWySN46+g019Mx0x1
+549PfyghpRHuDRH80ngbZLEAG2awFWMtqUz6Wq1+giTstXBL+B1Omk0yZhT8pRG3sVu2oucIVwb
oO9WwTAsYEBjf2UmAd7lAym1mBXdjiS6RwGJgX6CK3oXzGuRXfQOylVMViyD3YZMOtW9l/b9/O5c
PmkKx4HA6RvAh4mdmEOv4Q4ICw7xQ1f3ivmS7st0nPRAr2ZG37wJU9b7KQCYJfkMLUCkycvDO0Ff
6Ttyrq2vv/m4oREKpsYtVGUyg65uy0GvBu5IXdA9jTJiaRh4vFqDLWLnNqv0JQCpyntWi9yvHxGj
umaTkRsrTIbB/l2LmcgmsWy/O1lfuMhwECIlKDPhQHu1VmRwQplbsl4ibt3EHE7iFTcBSuNoKqG0
UbJi2c5nJXgFDvtOXZaLlYBcX84FaZ7BiusOu+1xrGsuJrZaVN9A0uAq1+JIw8y0MW/88PZ8Pq1x
ind13rzJuIvCjaLVVBaSY/5MlnOYQ8eHkP8otSn6aY5JSyCMvs/O/K8WcJ07get3ZOW0dt0SXJdu
jjzX4HFIPbQntEkovNgDKYpNK8c6V7z9RtZD7T0lqafWSvC3vCo22MmtFIiouWgzO4mSjSKxD8Qa
8INq/mFKr1HiW1cO7y8OidwL9KNnQdrtUtJSbBoL7kMn4kVQnXekz8A6Jeetnv1iPAiSv752BAwb
+39ULZYFPgRT49mRqX6ugb8i56PHrcLkEMIRt78/4QViS7VW67XA3VoFYb4vgzlgqXyiaSgQD5YM
dJT2JqRgo+TMYAIreDSroJiKoDG9GHihvMXK4ZZqZDbPGhOSPrdQINfiWwtdLSNS2qbdtRLM4akr
2CGMcTd/7cjDQhR+dnnp9lDD/JHUfG0Md7Lf2E7nZV2Eb1l2yRcVuZ43Iimy9mzvcHrTZk5p9eeu
9jEqQBeejH6JImDETbp6S8SGwkSsvLPx3NIv8SiwY5A4wPcAeKcDNg+yM5RLWY76HcFA9AVJkX0D
e0UpRs6CFs5NSVXt623nWP6aBtEKw095f40sChS86pm7LOUIQkY/q06IJaRoki1R2rpSxJGoGMdK
rW3+ttVY/79Y4+rCM3endNjRDVgrKOL6EEJloPd/BZb1tpi8/FYsypvmsoCHKyNRVsZjMG8EW+Jl
/L4BDxeOE5zf2ZvRH+KVGfwP36hUbQi31cAOSRWrLCaf2kpxRU3jaramFLdcfHntAFyTEyS2Kdbx
YtDFrcCMQmVCz0xNDBPoNnT8l/EyCEjWXD4rzzhszdL/zWQjpsliaG1Luh5JbfNFFFvq6ijSWp9F
295/G71b5U18KejpaKYNTKUKMAw0yoWuse8tEqojacGquvTnCeXBR0ON6nfh8ZGbrog0K0qFla+7
M0ppYRTg+j4zFHeWUYyNpr79ISfFEJJUogN/cJCEWnhOVPwHd60sIAzlmKtwnVxWtc1R7Q63/RpN
lcBtD+eXPEplzkD5uYxskn5OFEhn16bcqEVaOzlpaK+vxQzEmOtW+jX3BH4fRRq3yf5ogIJeQ/CE
rSUTpWqbY6sZgYz64AatrI/s3mmAIDhvkj9z6H14Rb8/xQBR+6Qa1MW+PTVGDgmrcZxwpLQLPi7w
XWr/7NLI8TsHkvOxIIjRlzPRe3hBUuvLx9+gC6gxPFBMT0eDyiHNLxkE8s8rMGidFjkpFHm2tlXB
IbApX6uZUJZwstGuy/plOTfw0SMpzWXrpT2kUf5eNgYmk8Z65Da8koBdHxCqoCHk/feNJz6qrTb0
t6ri0GIVMa5bW5QUyV8YRw9W56oo8Qi3bJjpd04IgaAMwBOsR3WLdt4T1i5VglTuPgWqRgyRblwK
jGLgUap9X6b/qAvfUJ+TzV0zAx5KeERppYrdG+ymdWjZtcgb1g+0O/JXQyS4gSCJ3voab1sonDNT
fqO1D0evA/masUmHx0B1LXpb7RHx+eBVnAtcECS08KnJpFBnvVeX+KjSUqQy5hKNIc8bs3HqPWe1
uU8j9fASLjb1fW5FdrsavFWWpH1SFlZJwxNYu16VB4hSDW42yMB7Iorz3bWqUCZSRAOWSLYkmSVV
0b44ZK/tagmED1Ez1DzMN1EIAye9PppjOoR0f2+q0rAFG+ZKYwUhyfX0yRxbjlFkmmJ2sx1Q1bsV
S3Zo2xtmr10PEqOYPJn6fT0h5D5Vjgn5IKKgxRtYwpMKgsVCzPw91bHsDbYChCnMX7wy47UvTljV
Zf8WM6MqaM+CEW0o1EyZoYVXaAsP2EFCZq/t252laQ1vDtnRIvgI/4xND4OkITA1chz6T/c9K+8/
A1uISdiBZdHFf7Hu+nWBjMlJa583xckzRPTSn9yWhrakbj/eUrfhR5XqyxmMtTyKPuWfGoWtGeQf
x0OZJHK2CQdHFOOC/S1V16CfXMSbcHgdFn/bGF5BbFbpZi6L5w7V6C7fGimuBE1VQUek8HBb5tbA
oU7gc9CzXpILBDBzfrB4cRLC2D1REyZHdwdxrmJ1bFLjVeff3dAItkRHddt4Y3LiqF6qNied9sQ7
1TBWw49vAwTe/VjLyYby48GKvmlphaGUQ+eytmgurqjujxhxJPmI78rEyRRgb3UDAjlgw4K/O49P
+zJ4lNkNy2O2lvKmbzwor0lGIhGbNMEO9x09P4Ofu1IbVKj3Y73WX5LGpqEahzyIw33VyCS+/kPc
stJ8v5FmY1xdPFBgN7vsJDTAkPafkc0fpUv2cpopEluvzWKqByYo6al85Am9b+pOIhdvDjUqzr/O
Ut9p2GOFLmZIWEydy5pafY3m69PBZ2tcFRUfaRZ3ypc6jyL34VHOnaXOm9xxfJQezyfqp0NwnPK/
uR58RqohPdVHvE+tUw5Y/BPjz80Szh/3Sjl+r326EkDXH12XNmb80FlhdZEwVMdiA4t1MVDmvdUJ
x1pTQX4u37ysatPQahXofks62gW6pEHSgQvj2CO11s0wpVgBTf29c/5N1S+LhPdFIao6eo9X8ela
Bl37HckTBsw3oJ2zb1W8Lls3Txt+lncuwQGET5l+SCTfCTOYP53EVGsyhw+rhHnx6HMaWV1RauxF
D9M+qiSvbZoaehKKEvWIl9O0Xq5wlluKwvkXN6MHqQ1fBkDZP9GISuR3BLk9Ay5PB/5cwy+wLLH2
1WdgMpn4UV/OCsrt+b8CJwEc1jOOTHNiXy9GfeCiI9bIHNghIMzBMcwlKPJl1QaklHxF1ST+7Lhv
VamrePLa68/atci1M3jZ3pM2hz7zhjdXsuo3MGxzlI11CEnBFh4DZpyRcdsE/jtz0dQU3RS78/NY
MMsLYhAX6aJGjVXcz49FGqKRko11UfXk2PCA1uQw2YHB+C5tgAkQMTENsecYuqblig6t3Y1eRW6c
YThmVLKjVXnqm0gQKcI92+dYh2/p7F/rsOfYLEZd5WPyzVswRBSxsM/1PlS6XGSa/tCI5/DrNcvK
+WFF28w3jIZOh8tnuEtrA6PujYx0UqPSc13ClDhxBMtiGA3YWSz48si0TgqbUA0RTk6PmDQ6H4o1
hhWDJUCdyYXKT2n30Pzc1l+Q/SPC9i7P9twGxNMUHN3RkX4A1LzAmz+K5+4jFqHaRcETyyaaaeN8
UY4cwMGGp5KxMChuJSC7GYQdM/RoeU8GQbuW9yxQUQe5ywgLoiryIeG0b+gFgCSf0EzbOFGr3hKF
sETLx1Gjg+pYu40J5zCfNmWktf7Diis9TEqnIrW/0UUk7Yvh4s5/nhLFbpo6QxRFRPl+ti+fhokp
gfE27psHHllbUDeNmjT+Wu+FNRpHCWl0k5tjtRrwpNVA9sgtEYgbyvMLTTJ2N1R+07ynmWLGGwvf
tQANOlLkIUoU0lMFqIqz3heN5Ied3Kxq9clvUK3ZpiKQX6Zhu6NMWpdjYEobPpwmIfnt9K51tYBD
gfhtUbPssUkc0Dn4MYnXUiGLXqaprskKYLes0TnV8ES3tYki0L1+EXsEGjvEFePeShZmFa4b+fHy
Y42/VgeIPK2qwkFS5cl7PWrL6wI9g2Phl6MdZ0odktE4IYYwcQjq1ck8Ksmeb2aSo4ZzMoS716hN
95cCPoe5Bfac1cxo866UQD/7fP1qoB6D1+W5rOTFtQYL1IC07i+9obqa2TbOs0owYXTVOApjfAm+
/i7ZsR8dPHElRquodmdCJOiw9Lx1d57rCIRnqfEGo/TMK1nu5F3PGqaxoYrtVIiBXhjBVTVkecl8
fa9IfcG8J8KYatRM47V5hFQaO1XYPhZDie/qCtvRxcBkPDATmYYcdZzqkf0w+h6915gQ4QjjcB3H
m21EJWOEGvfvBaxYHEhsBJX+FtICyA/tQ6WXfi7THn55cBjx3DwzXR1/bDoiYWFhDPohyFoqfZ2A
ZX7kabOtKJMSsCFGyFMzDphCEPhRIPCu2qjQVglg30RynZFyL2yreLtKKtd2SutsuR235j9pDFTj
1AHx1rg6kLIoDAo88ysRJKKG1a3xnxsH5jujQLSjHLk3XX6VY33dSiwKAR2rgElESqx8F91ndQiB
Sf1bDjU2I/iwCXGEsyMKmn2vBzizqIyHGcwGt3dNvu5f8T4xEy3K/hq9QT1q3Ajs807etJf3yieb
+l9tk85tfJT9BuBwX5bM9hDqtjj3aQLHDahPVK6helfGHtLJyqQCiTQPunhd3+Y5+N5JxRmoSr0c
L1rbW4/NkghzVccmCJI+LrnHfPPYTQ0/arKZWGOuvyOFY/9ihMQqMtDBpv+BKfR+sEYxw4ARM3dd
7vZD4NbsxSw7c3gWfkvjjAPrioFWupqaUwzexoEeoceK7bZlxsskN02QLfA7LT+BAjpC+dxrLE3L
sGpQQtu3IVduc1e6X0AUJI/XRtiaxTtbNgbShVL30Ix6UtyzL4M28uidGTok3yZTeS8TUEpmPb/U
L/Iq5lD8D/G8cd/VUpo4A0nVMuQ4ILSYI57j1XV66aLoRA2JKtTzrcA9AzU4htIRQ/jT2jaSyvNl
qfwWV55CVwfqTYUjiubeDE914WgY9Oy0bTuyj+s7dfj97PF2gkILzRS+i+BzKQlLgeCl1E09TUXw
owyw2ok42iut/oxZ6UcC1nPIgRqIzZdLfAs9zsy1sW8DtofGdegj3G/bFJBA4X1FvoC0BdgAZjpJ
EHs1tm6asYhIYCFBzxKThKzKdMhvCsCyNoi3jKyuns2k3QC7XjmPLExZ30GMFCnhnXbNjiOTGlCg
wPCurG8mRrdpNsV9WDpjqimj4ZFCB6fs795j34NvpMiZIs0tAh/x7i2a/5zVfnAcjt9rmAZgee3s
MNqUwY3dDVnydZ7qqRXPE6u8gA0YEGEBp3N7yl8i38bpJ5sqrDkuj4ICR6QoIlr9rJyNIAIBboRV
IzXotDN17+lLH0h0jl8JZ9Ebp0DzSVEmw27N8GfhMnlATmZHTykz9INeUq31qgICHmwL2VA8qpEe
31aASKrghDbNCc7Uba+V80nxsuqfxhATuCDQEZwddC7ZCWRwaRRehE0w5YglxJ4LocGD00mO/BpM
LFIo33MS9RfW6CmLCcXtlzxY47RbLzsliR49xApxwwSOmnWFNiLlAKxZQgDCWOro0B8hI08EWGdX
INBmUBYYm7UhPDT9ArKGH7J3YGx7TAqzJqNEfDUo7HsxJAAB7EwTqz0JBpvGSrRmRam+D4kNbrwo
LmJOld6VvBVkfdgzm5Ur5NMDwb+aa1XBL0bnAabDs5zMCvtQSUp8IVjTFxxu97p5gOlpgRKcdX/6
ODDtMMWmWO/KbLCc06fkB3nN3y5TBR0NhM4NCg64dRF+S2OKitLAmSkp+cDzNTPWSqlVihS14LBa
lxRVpzN2StCbFfd8vEsw9CqccQ9jq41aTxz3TDC+YkJPPhM+WRVXuZRSAqdlMEGtX6XwFXS4ZV03
kJ0sRdTaDPzbBsFv7JnPJWBolCWRn3kG3bYSRCk93LwCZeEJPrj48scC0BMJ0CXrNSE8+bFrsoDR
h5Ac4xGdqt44UfHp6WDacb2RBZwZoTVKrSXQcigYid0cgT0fFQiSPDsjLZdVegVIAYW2s4RaViLI
rRtXwDoesx2jdEjeVesOOpJcG+dtRXd7au8PC1cxBbOrPl4n03DVR+Z93iNkS1Nd6ddrPrf0OpoM
w+6r0lvT0K0JY0fCrRqQkTycCjKb5b/gl13nEFjaNBRuN9SIBqMm50lGoU/qpBRnAWvuulF72dn7
alFUvLORFEfMD8+UW0fzVWy5JSwvwaIIb8c0LthWrCCDsnM63ngSV8HZbKWXnRQNmD4Fx0YP2zdi
V/cv5exq01l4v98B4XepExXFytpedQo9m94wTRpzvA0ZeAl880Czu0wLUwXNRivE3qlsVaNRGDLy
sE2hnFEWz98pSRgmvUyTm/C9mBNi9CCgM6I+2N8gsUbrWxC4YVNmNQmCVYg5+sbq310EdSFIbDhe
p+qAJR32Folij83MPmBlbG87BjTuvf/qWK6HPHEa+vQB2I0uGhW6436gP1O+8O1vvOYtI2HdY74M
NRFijwijDuOkw+GrPJJchrMHnWJ1iSve9w6QlJVtjps4cWOg5kFcnRNyn9b8GmyU4XnVqro267lT
SWkAAxBcq/CYoUHh4brB2FKBvnBzLzJTtzAnMmX76UFlYa/szpYKflbTwBeYJoLyaTujaW9sEiKO
ExXiOX1C0Cw07SV+e/UYnLYHXLZfxmv3zTvvM96Adu5DPL180RQptDpxcZKd4cm7c0t8GeCKMHDM
O3x4j4g1pLgSjdyQs/pHuHNFSB3Q/Ryq0lmVtx3ZYZ3a+Y6ksL9X8AHN+6zF2FdeJhxJskwvH4V0
uIyMmCmd8dW6NzYk29AkNShIV8Um5rKiKFAhlQijpSYKGHelv22ib6fJT5h7aMOPQf64uAB3YKP5
XNpXVGo6TRnLd73VJVqh/nMHDQgktGsFnl3grARqSlKcc8WdDzvE0d9RYvu7Xxm0A7S5JmVN0hlZ
rXMyD0nx66C0aeOHJk2D+5FfVMIJSxo4l7vOxnbNS1uSXrlElU615yvYRq6uFXfAloyW7VVPehek
EfJzjjD8mgjLL/MkoGkCs/PmXZhrxcqDkwvDEuwhYgMYfAHHkY+c1g1EdK+4+TDT9/LAlJriFmv4
rBgbdVdkvUfToqq5RyvkWio2wnrkZfhxkQLTRQzvHFNKnuDxpmuP/WHgpaCieJ85f7jcwHyEozhH
e7DDxko5p+XShGvxL86lA4ALaVXSumsgKq0r/hcDYlA3JbrOzPQJNdIiRa/uXQ6vvG6uHHT10B16
Z/1/mNR/rTkwDnQ0ITsKXA0zgjqvTQ97p0yzS6psGuClWx+Pg2ijDznNaeTkj9sKyGi+Dc6/zi2r
SE4jOi9HGHCXCurgQS0xu6bAseb8t88IXzXf1MEdowlsDrOjg0W6HpErnFiArRviJS1fn3ax8scN
7z05qaT21h7v60tBdib61i+VRmQSm4Pu1J83xlNY66NlQykhUxU6rPz7jBiWB5LIh/00lTdCFSs1
mJ2Afjhe1mK8rNqhNLt9iASmMIWD4aWM/z98wv3qTfM/2ecKfPiJk7PUjG0KrDAnI2mc82xMheCx
Iuad88KkBigBPwfk2HnHEPX/fiG04ouABuH9iH0xv2dJq+1XzSXKZSqGvef0+qaBGJCZyx5JRr0I
JBRkwXvIx10i3guq2aGeuFO1V3lP5XGL6EN58pYj/q2q6WyqiWdrQ2Q7erjWYUrSti6pAtut+fg8
IuBcnrGkbsFAeO8xqxmmDuv2UsfOKKQoLajgkX0Enx2syyCdPu1CFFXlmF/BB7R/6yPxsiOqtg+2
7TRDo/D76Bj3IoFBzxIBw+GhrQNhqyZaeAof/mkE+v/Kov+aQjvD9JVOSNTcPWffkLTXmY3fgM/5
1qXeCe+5/Fg1Jm6z3B7Dw+YmyEBi+1hc8h/tcaZBJAEhh8y57GUj4LynIx0H1ydHnPydoH5H1Z+f
4L1EZZXD07dX6UzkzBaYhfUO3/ihHl3ilnjs9ccqFJ9O8yz2XTE9sDwsyx++xCB38QrUbpd3eEWj
XzujDhT5oVh4UkGr9HS7xtqWXPwo1pLZHX7Kccx9EfJ6QpQIuOxv9fft106lgiek8/NumgX0B/52
v3xiFB6N6CIJuljyRNNtN/7inPul6iz5XPq6ylf4KACwXl+JpKDa8ZD8sRQjeLwxQmyGVThyAmF0
UqzE8m6g0LTr7729f5XoRBA+AAIFpF8f5ILe0YDusAsSgKx+Z3djtVd1bciucr1bVOGw9HmSTi1G
qgw7ypzXJRRJoHJypv+/cTtANv3uj1Xfo5y4n/3ZeYB4dD9hBMOKkWlsIvK/wQxVezhmix5/U8+X
74dCAZt4G47aqTGK2W3qbjV8C9DklS5XtKXZVQZ3PiFaAickEolYCCdJ8KJoRZJN3S0tBxpnJHGF
MzjTm/6lezpS8oKHh8rtyinK04XTm0hvRxqEzGYE/C2m27WZJmyd91AMRKrllVqSdmnPT5ivrLx/
GHc6olVHuRrUTfTAgEawFZyw+3KZaqul6DbDuGh4A2cvltywjiounl4VTqbuim+8ULINd2mpXk4A
ZXLEftR0AbU2LdkP1bGHCdZfqypCt1YkPyuiDlE49d0ClnPcklhq5eZiichTtmBrpzlVBfjmKXXB
ztaUTEEhrLmy/rXWLkzg5vXbgeunaqVVQIBsrRiMmEbBj5TDMQo/GYGWaLgmxWGy7PpKee4m2nkF
UwUcYSk3ggrv3R4M+erGGMKerBZRgiPAXsoT+NgeSXU6Ls7ACtr8JJPMHWeXUsgKtu2BC9Yr24FX
VABT/VxPAlYCOLgZUfb1oWjXJaRUjOwZp95CRwFkUUjM5iUSimOLfTIQU/yWtkfOXRwH5VpS+TGe
e0lR9r+ftKf8KqxacnonJFmmv36QI+Iq9CDT3gYkCNc66TAlJSjqcTlJYeMwEU8IFz0sXp4O9JBy
gP8BDNSXeE5YjDtuJfEukqCjJibWNXydjCnyc+2uXBStU7dXxFAGFasUpce46ZMSn34uXxKbxJDJ
+/+vBRCrITm3lFAR3T62RSaeFtrUrIx4JmKsI9sQjtqeovJswevW/+hFsemRyBYk0RDF1NnMlFcz
QiGRtAyjVyD5hWWshDz7OzbJFCd0mjSNtPu+zYel99Qsq+I38wN7V3M4vnA1G5T6R+uVdYwORwLx
NbrDwjBDa/Rpp7CZl1t2DSdsl3XapQWv5Va+xitbYByVDdscL0YmZvKsKcFTDr+6zUzD95KSQ7oF
Zxcy3EVxbWNJkrkxDsm8yrOr4Bu6R8MUtTk5GQYmYY0/0L8oarISCX0LiXXj4VZXAExs9hpsxcdG
3NxTpS45jEROJdc5pXHou+hE/8ZMddsY3hHNtbeAO14asijRtNfhTy5+/6dc5ZMui1AotALUsyJk
eLdxmPrV339w0N5muhr9ZwfgKnRZVqutf0e885rlYZ71FfMpgBTUxo3AgfQvXMP2IBrJ7x441oS0
JMKBagldMUoZLtCXm5FG374D3X/YE8bYivmz+8HWAC0bkTgItGrl4e0Iy3wyf2ivoFJTmGQD4JF5
VJHDrpVt3y/oXCUdU5ynXCUbRSC/tr+UqNfIxUm5iGQ0hy1KzUBHn/3hhJc3aTfyMBQyKvTnUeKW
aXMrPc9Rt+FUTdPlwUmUb1PPCJfcAa6eKki7LDJHAfu88+XE0z/aHztBaIdjhO1062cljbSB3a4k
S7yv9OM1xPqDj9jAOe5WHGeOQUM7yge+A/w1zTeu55m/39rBuPFUd9xPR0I6LxAwbK9lWjlfWM5l
ww+p0o2ZMMKXnK+rww9yhk0jQuS9PMWxjdsMaJUWESvU+JJi9B8BdqXWYYnE7N0CAl+t2a1KMhvo
CiM5rzMXW3xNCjcHsNvI+M8Kimu9c9409bXBT+Il3Vt3VcSY+YHKIlyTSKt0wgf6Dae+QrIJFD5r
Oo6J86AxfTTPm8wSG5Guk/guMm5cXebf/sIBYkpd/EuJzgxLlC5gQt9mKjAV1LgaPwHgiMt4Hvs8
tdhuyCafDTToxDv2J74qhI6R22NPFqTODFqb9vKjAg/LTxpaV9H9AEEr9K6CSCZdlMAtFrIOupFO
cN1VOjWZZ6C8DWMIJ0qDAWhltZJ3R2o06OYi4//2UKlV7ABF3sGrf4vP9uJoZfKeP2DG7mvb91nd
cuwMwc5gW407L1x4NvRNz2/NsmEdcvLjS1SBhHJerpG9QAsUbiGcFjjanEbeNAij1A2rr8Vb+Zq0
WWYnKGBdZKf/zzDyxSYsEngWDKvwrD+4QQOujCvtu5yK8NbP7pPqOyBjLASJ9FidcURd+BnDfO/R
yrgIG1EzNFf99YaxZ9z4c/EcFSNLeR3WN9kRcpvpW9pg/S2GHYoiCWgpfOjaqmMrLb9ZL3f3j4BN
cPusHwCiM9LB581Rx3u0dbuEwhekoXsNblhfGFsb4FzzMHVQnST9mPdaK1SnqFPmd7IJBtQZt8d+
fnRkZCFMuB4KU8z302BZhCpBX210eppcD1/UYnWHpE2FSC/b3nATt/UiLIrNVoiyd5QTNoLYvhSM
ixHEjXbeEJZMnLjoExZT2ZqLo/9bXn2HLt9HjWFC5IMOKSvGtu0Mb99jvG8jgvfEASg+ErvxycJK
HefezFarTWTUJqjXjs7Im2mL+bO+M8IAR9xE0HiCYng3GUdRA2XUpx0wPTYR2BLN1kicPy+fENhg
0XhXFi9xfiTcvMtoSiSdVZE/7p7nvo/wmPJOVwIsdS012e9IKns5K+ejGAKhCgZIo+F/glMQ2FRz
ZFeQg9J5wSG/XPlOJIW4NkOIFbrjBVCgzROvMbNQoYYitZgPK4Aml70MbU/kNxRv6oczWfFGPpxe
XwTctOX4EKmmP94u1LmXBCnGPO22NscbTOKA5uVaZdNLHe6y3wUk9slH//UuQpbWJ5/v6xivX4Mb
A659Twq1v2vXARqRhvV8WyecfLyhgMkRLVox5TGxrhxugTp5I/JmLYt17uvun/PBrwG/0ATK+uPa
fUouj+N4jNj13wbTfWWTfiL2c3Ck8921OLJiNYCXArzzeRAmw90rxH7wMOGmSZtNsDuKeRTgbDLA
VU+zvng4/sFu54H8+RWjQDnXlCP9fLh2uv4muqDRyPM2+HwQUP66ExzyUW4bDxWxV8z58EaXUbOG
/XaX8F9dWsqq9NrXTDVjg/MZoTVqaMsZaG35IbwlLZy/iAGD8JJ2zhy024miIVMCvHOWohftcuoa
ecdqxVWtSnvkkaf0hXJDfYgEWD1ziXu+/ysuO2hjVnlBn+EeAg9/cfjs2Prk/TI8TOPBZBq8Tctb
mNJnIPkUcGL21rIZKPB//QxZrMIdomeqrEzK6bf8hCdctGnpBru2PTwGGXxo2dP6A8JWR0259+IA
IoVJBIzeTgg0KlVgVmhXGMJkcHoO6p36HRvd9J5QJ1iL6UT3HCbBeELzeC5Zz2qtQoqzLAgKdgeL
SmrQsGUBz5BSIQ9FAp0n0Yt3/lwPk8drBhpM6juBKZXZMelPVjQAEPtQohO/RRECBZtC7sVKkilX
a+LW/BKU1yQTay4AlHN6+TXfe2Th3J3D4bB1O3eCaem9QQmQJwFG7ozkaOx4X3yh/lyyq3+WuEDx
0ulrdNEqkI8uZ2s+gEhSzHo/KBFOxQiuf9ln5zSWxSDD60Fw7xpVVg9YtHMa32N/mZ5RvodBYsIC
8lEhrSkTZwds4OEdmX4ShY808tT3TpBsgG6oZRU3iCkbLHFdQ5olFo9PzRYiIbrs/cic2wGKbxt3
T7Sf5b8hi4nCn1eU9C9eoWjzHGm4KOmWiI/lpaYnl5mohKeEHijI8dF4iC2ymVy9quZHrTTQlEkV
hB0M6kGw+5fziw87oIsvmtXqBKcQl3+qvlNOMsZeGT4OXBudpozeDonRk8i4eq4pBNM758qOhKca
f4jpR966p2leabU1UYq0MpncwZed4PwcWf4FFRf+kDj4qjwrUNPTGB425kPSGEwVy+8W3VWt5HUr
u6P0hDvAGezIGxj3QW4gD+DpTedWMNKA7pW9fAPg5Jvc3ozqjduDNhp0MSx5je+G6O98MDMtzWsm
7stzY7alrGTbA1Hd5MKTBPTgQOaIEvITR2y2prEF/kGT+QRgTFjlO32CVnRqZoXiNYLjCGeZjkW7
CHXlqAO+SICo8L0sTebUAWMlClk+/vX8hBsANTLo5p+k/+Ec3A/YCCM5q8+fzXafQEtz2X2PUNo/
EZhfFnYHEaGWqsD1MsH2gkTKkcdNxW75WJIfWeDwPz8Vg/8eGlDHZaPk5HgZj3lCqMBAdT0VS33Y
bia6+3LbQ3loYLghCTLj5laQzZFSWUB86f7lCBHPkAd4c65I+WVQGMZNDgMpwmpbcEyuTl5Jppgn
YeDroZqXO5wnh1FYF2+mvvCIUcofVWlznTqW+lqM7LkXitfHUfxc+MPXvUTuon3atIXivyzvRFMg
NU24/Wrdm9WEFznZfJvHfGTv4xSM5qiLIiKeYFCk9qFytnJwembnWZdUZEb9Cz6dD3CU0yKUwAbb
jHmI3gcMv7PCi/z2gwzYVGhJ4hQIpstAPd5LQXjwFGzY/RsPioafnXIkzxAVrXUcVxvxeHsDgr12
86w22kn2/tfyUCuFX4aPcvwoJlkmE5SeuASpCNR+qdoUS1lUvq0zfSV/+AIHNJm43IzpSRPpjKKK
rXlpU+uNgPYD4Mcsc0BdB9Wc9E2oXueEso6rQAey3HVSDcM1osudqVWiEMGOULHqZJJc3bRWhYRt
sP3g1rCEuQK0DW3TQnbrHh9GKer+uAJ6OFYzrim+oS8eeNxQgwoPmTWRI9yeErD0JSdPDqqfZqsI
Z2T4mPL9wply1BiG2XuQ1/+IPEMkPs+qer3fZxC4FLloPq8Ofg/JCSZRZbiZEvOL6EdwNXtR2wNS
jnw+lgkMLPdtSdzJfTnzJRTGt5xZJcKvLvtnZv/oSILz17qRSbN5BzIat5rp7hOGdZNI4+RklCG7
Qs78mYKZjkZlNHIFxjGC0p4doZW/f7hK9imXo5xd73tL68Q9pk03rMySI5EzOlYz9xvYTqh+unmD
P+Bcy7mzlISOoTU3FWpYOqYbQlFQRG5LizpOh7gI3QPCqwxEiigYD04XhgFmAup+BeZydBXv8Qqq
7ZskQpvWxVm7xEy3dUH6+eyW/yXvJ2T1eHS1dTyKuUG303reLCCsc7J/8CsLMJbVuPW5NHF2P3Dd
5cET+78OBl5a5E+7tly9575XBjOonZS12CYFg8OsZl87c4uvr6opCjuF2JMFg15gj8iPp2Yeb+SN
zCgSl7XwydfBIPcEanTFq/VT5iSSFxuMen+zDXy0aIMLIfmGjj1p6C8lR4ZQjKN62ua3JurIHl9y
8wb1GIPXAoaGsf/op2Fw0SCpy2brrb4WV6O/+q7bJbjFk+ffLL2KnKum3/DvM7PRTOVFBnSWVkzY
5FOR0Fx8GHroOnJjW/5QT4kjlP4KabCi43apjgFHeadHVAegI6+6zVN85N2dTO8okkdkxrfx7bux
kdugAHMfoVHs9aIKkBzfteABVP6uno5fDMxCzNrzsnyLXb3KXQMr8Ar43ZqHKCR/vp+hC39teruh
1m95lfVEXbQCwq1d9tXKpD69tqzNatRZH/YaEDGGbcM+84CPHDowwKeW3YPXZLY3j8UD5bl2Pv9h
m25UptxS0/4ti36rFKXXxCTomSwvU/ynd7SjSt2PFwx0btmbEvBJ+RvVXFcOYf9nS73ZkimZ3idL
hKPJ36lAbHkT00Pq65ou+v7TCzwYSryzaSJQc8SB5wDbdz6DgKF6vCwdDfZ2R0yCpTYlXcKpclda
8ZZyobPQb6OUkJBTsPOpNlyFjYfk3iqX5q/MpC/ZvayZ9O/WZsL1TI2rC6DonbCL7pGuQA91qGGw
aBQPORs/AaI6sD5yp5nBmMOM0ZzETYqbiMhy8BoAS7XCw3NSNi7oe33FqJfrlqJjMHPRrtnYH8PS
k2J28aqO7MsokM19GTGWtUySyeydIYLExqx0Sw+JXeSOcU0Z9Nv+mWevuxp6HSzYyzy1RwxQZU9P
T1PyLv/wMHn7VTHmjnWE7G9IDqHEGdcwn1qQHbi8foiHoHGa+YS/jIIKM8EH3x/dTR6krxvW26Ac
UpQfCaUvOzPTnAPmbY3Ps3mWioEHjsYyE+qRscp+T2FSZ1NajE+ylxF5aYsrFJxryFjZ7Q0wKwvM
COA9vgdVCE9sUcNkbyRYXdZntY2cfpN9s9ix9uBP/LzmQmQAj5UI5F2EqyCk8zH2s+kkAYZg8yTk
DOfFtm1vW2m9wSjCPjPnOLoNGB/1wKnp7/vSjs0qeZWbWRyxNdsFJJ8zxB73SKpn8txY/K2DMq08
DE9Ka1/HlUGS3U9KMVou95FnTDlbFq4udklhAwUIMIjcHYZZr5NkWbVDfIcG8g8wt4X/g87Po6p6
cOkrbeQfwFI90r/EpGMAwODh1Xl0QthVBB6qMYzqPZs8h5lOrJrtimZ58MsJCVbOaNKMBDJt7+g4
bXrhAsUUChS7CkO+d7oB+ifFd4yoTbaavwAACSFP5PDSrzkJsI8LGABipDs3MeGpwVrwCz9nRtwq
dgo/MWnqg5pamroXHYJ4nAdvwxu25i0C4Zl3u0/p0mSwYx1cX18XspWTDWS4tUz6rDPFbzOn9bic
tybeuI4KztxaaIOn2MYK7tYtNWeHgQCkSOs7VHJYbgPCrxYXfANoO/6rpGwGX7iJk37oPTPY5YF0
JmT5IekKDTWSkRkRdfvTZRKNAowchuJ8AP+sSqLtjyY/1qwKSU0BAsdaAO3/m1vuZ0rHV7TXBECK
/mNkSCG0Fd5xI9YoAiYYPGji0WXspB/EPLGODhwdLSmm5lG9i9K3+uWFxa8OemE+mIDFFdaYYjiU
scBnDn4yXcZI9B7qr37NaNgbeRDie5055raM9gm0CPQ7+Sb64//qn4NHJC7s3P4FUYx11cX6ewWx
ytXSyHhTOf90awBad8/svAr62zaG7UZyk/duMYzicIgvxfhTPId8fiENlJ0QAqDywLydYzYMHC1p
hj3rNqdZoiXD2uDKt5flMOlfAB4b5tDdNIilrAyrfqzST4zeMwYtRFR9+Pk/qJovjrg9i/uvZCFn
DcMrsGVdYUqxfxY5wZ+rlnxylWDbGzK1HKsTjBVCXqi1Xz/06dkYg3mJTeEu0fGtHT6dy+ZC/iT6
QioRf+Cwzf7GiwKhTHXby5S8NUlAmhffooFfyRehGfOfz+DOiNtZUTEM3nmVRu0cs9iVb7brNPQ2
2iwPKDDTxNwWVmYQEu7sPoBGWApyElnh4BHcAMSzSf4R348Nt72ykeipK3AIaQlxQHXhi0iEjUtK
WPR002pdl+yivTZ/tMElhBjhncuzXcDFs/FsigozG+sp+5sxPviY6/x34P7/SMXScK6MV5UWKj9G
3TvmSMd0hErWq6JwFMHEVGFXuJVW7S2xs+batPSQMiY6yKAmwWlhDojczHeMMiiJYLg7BIqrH6tw
G3YDR2q8yooOkQRQnPfpUR99ctWc90GLdLsMESk/du4KiKA1E6wY23xYO2fRJIoFCsaeQkZm2MLW
Tkm2V0mbaKyZ2dgZb8oQimPRS8U+X0h4TslatMs0QYiz6haHDa0rt7tja0GU/g1yyMDK3Zsb3Yai
TtOcjLOdvZkAzt7zHDmeQLBRym6iDjx6bx8SCHpO4eZUZW0wc+oasxIcnfkqTqziN9o6qK8OKDYl
KwPhwwGL/nVq+/YriLYXqAy/3clbVdy/HSkU6KfGxrjDvAs2eHEbwnpP5K7RyzJ8BVpR+GxMLYzX
hnXm9COu8Ji5ejMMKx0CQitJdMnqFt31CTHp4y12WB8FjlBSpbQhwi402cTA3vactQG+E+2zvBNJ
WuzsI1wZnAMn/RSY+nBjcKsGwNnbutZ0WduGOJQrBCH2pjpwvgaXtYZ7DQ758mZhtHZNolTkYkRc
Ypxr94I56rEnGEGosKABko3PGQnIyEGvMy6MUYGP+QloS/sOOh9g/S/rlOEUBXKvme1Yd10ESwAG
BFjHl126VxKanLFBYdQt7LO7Ggc5RPS86mfrD7dyyRWxz6NIhxMIrIIbUC2XdB2iznmVIu4XFiYn
6ltePT52OtfEa8CrUYR98J2OYlhEy06YZrupZAWXEaY/qaG85pVDATxsxTTzKeHiIIU04oex67C8
+Xi7iT4coQR/ehFm8+4sEIgljjfMyonto89uwQD1Y9xnAhQFSTU3zVuwrKhTJREMK8NKuFONQwHc
ojIW8yk+qFyqDlAMxbCkfqKMoGc0htIH0fskei3eo7CcvBCm6LNomu5jY1pH0gbthHx404TFrQrm
es8+avQ5DTpcjAiTL/5Z3dW9KcTpVMVmbE5aSHw9xHlgOhrHdhBFtu8fFXcc5BrJNBE8WuLINxCO
2WCnQGopuraL2L6Iw55Y1IevJdcU9rZKXBu11NwHfhFul7wkRED0Jn3VKBnpDkohZma0YMgysfUM
Q3bRGWyKejC6kjEQQynyEfHuWN0KzQtO77O27OfrAQ8OpLeR+W4yNfwi8K34kfALQOKic9jsyWnU
hqMHp1uwiwby7Qa9OL2p4VFwSUJQK0W2mraNYZe6xmcG962ELd9i5Rd2OVkvvQDMEvzvQkq0EhmN
w+t4KpwiAa4h3ZUeykZlg1hYWIsKjQ+n2necUQAo5d/nJgoEZdKx4Mmoso3M1WVWjOvaOT51PK0U
edbGuMTWZ7kaOmYzCX9O5GBTHjGq6KbIocTCYGl1+kkAijIGflmc0HZYsR15lA6prLVFIx/E0NBQ
tRFxNM+Pp6evltck01epMpyaBGheD0POzezUpxwizIW7YJrje740GyVUvbS70kfDBdDZD3qNflYX
aqL0XrUJ4q7std20GmqczLUwtL+dHlHHIIIIg1hF4slDUjPWa9CZioEEIY/MXrD9yWKLIbfWV9bs
uLImYSpXhloKdRVwHRuIbSmkjci4DWAoAiHX9kmtT1G4tkP209ILIWF8HsGRlN7Arv96oqKgp7Zn
31e53CZ3T2HtZTVJ78HBxR+Ph7/J8nKqzVdPV03tjf1/Si61GxXMdjfaIJzRyWD2ooidrcL22fqd
BSAFUdhxXm6pey00Oi5F/WHkSRa0ZcaaEUYznZWReh9v9BVV7a22ehjoO2v2OhtlokwAlsAl7t7t
ZJY0S7T7PI+1h7hNidV1/1O7/HXWDAsOtipKYfnN61RfVhl13krqN7ZAhyWoiwP0cueRUIzMDJqG
a7H/Gbd0jOPP2erPOpqvT2NM4YsVVVUz1IQ+/c9Ur9hGe/hryLwI497Z38pDmSjvOEzbIiQGTrzZ
j5gsJjzH3KGXcXjiE5BVnLh7cplTvWsSnS7dYCWrWBQoWuHZqW7/JQKlnkfxBZxPZSLYakujN6op
JpklwYcSM798Ksa6ZBl2AirHhxtsLDM5peFV27NkQmj2KHzHoroMMDIbOF6XU3n+Qyi11obhVZxN
IRvquqbV5/6Kr9jrjha5rzVQGz/E+64cnUK1Tpk22bQC+RuElfCq5Y0QatyBk4BHCmzogU1JFn6h
GihleTFVQeGR4okpzg9gZbQMpe5uGgiP+CAsRJC9ydLbfq/fnyg6R2iYXICxk7ktj2iUsfAbKrQA
HIc3gIfaqaaDkxJcCKy8ZEXhwS1fxylPGCllXBDtS+WE7IaNWDBJKTATNgRMxtlEBQoGCBNXjiPw
e+9ZtSD098H9zZcr4+hvDSR+xCVxrYDM6bLLfohl1kWDQtThj98fLIFsixazK6wj2EqrnrOiTJEQ
1CY+GPlgMO5NHHsTiHdwSCvV4q4WCIv+ILxInMqAxDlendzHa4zWD95w5ytmkS0DNsjPc1b/TTKO
Yn4TBWGDsyXnL39sSzjEOCIN88L+atjD4efBnH1Uzoiqdn179DXRAdZ3Owgrk1TLjLQE4cI8WDoU
j7fcm4rs0zdxF8eluJ9fKKGvYOLn9z1Ef/4vrZ+sfI4QiCeyvF6Asz5vII57DAaCZAu7gq83zrXg
ie50i1L6lDnDpem/ljlgjgIU2PFmJTL2hoE=
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw1n;
use gw1n.components.all;

entity PSRAM_Memory_Interface_HS_Top is
port(
  clk :  in std_logic;
  memory_clk :  in std_logic;
  pll_lock :  in std_logic;
  rst_n :  in std_logic;
  O_psram_ck :  out std_logic_vector(1 downto 0);
  O_psram_ck_n :  out std_logic_vector(1 downto 0);
  IO_psram_dq :  inout std_logic_vector(15 downto 0);
  IO_psram_rwds :  inout std_logic_vector(1 downto 0);
  O_psram_cs_n :  out std_logic_vector(1 downto 0);
  O_psram_reset_n :  out std_logic_vector(1 downto 0);
  wr_data :  in std_logic_vector(63 downto 0);
  rd_data :  out std_logic_vector(63 downto 0);
  rd_data_valid :  out std_logic;
  addr :  in std_logic_vector(20 downto 0);
  cmd :  in std_logic;
  cmd_en :  in std_logic;
  init_calib :  out std_logic;
  clk_out :  out std_logic;
  data_mask :  in std_logic_vector(7 downto 0));
end PSRAM_Memory_Interface_HS_Top;
architecture beh of PSRAM_Memory_Interface_HS_Top is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
  signal NN_0 : std_logic;
  signal NN_1 : std_logic;
component \~psram_top.PSRAM_Memory_Interface_HS_Top\
port(
  memory_clk: in std_logic;
  GND_0: in std_logic;
  rst_n: in std_logic;
  pll_lock: in std_logic;
  VCC_0: in std_logic;
  cmd: in std_logic;
  cmd_en: in std_logic;
  clk: in std_logic;
  wr_data : in std_logic_vector(63 downto 0);
  addr : in std_logic_vector(20 downto 0);
  data_mask : in std_logic_vector(7 downto 0);
  clk_out: out std_logic;
  rd_data_valid: out std_logic;
  init_calib: out std_logic;
  rd_data : out std_logic_vector(63 downto 0);
  O_psram_ck : out std_logic_vector(1 downto 0);
  O_psram_ck_n : out std_logic_vector(1 downto 0);
  O_psram_cs_n : out std_logic_vector(1 downto 0);
  O_psram_reset_n : out std_logic_vector(1 downto 1);
  IO_psram_dq : inout std_logic_vector(15 downto 0);
  IO_psram_rwds : inout std_logic_vector(1 downto 0));
end component;
begin
GND_s5: GND
port map (
  G => GND_0);
VCC_s4: VCC
port map (
  V => VCC_0);
GSR_30: GSR
port map (
  GSRI => VCC_0);
u_psram_top: \~psram_top.PSRAM_Memory_Interface_HS_Top\
port map(
  memory_clk => memory_clk,
  GND_0 => GND_0,
  rst_n => rst_n,
  pll_lock => pll_lock,
  VCC_0 => VCC_0,
  cmd => cmd,
  cmd_en => cmd_en,
  clk => clk,
  wr_data(63 downto 0) => wr_data(63 downto 0),
  addr(20 downto 0) => addr(20 downto 0),
  data_mask(7 downto 0) => data_mask(7 downto 0),
  clk_out => NN_0,
  rd_data_valid => rd_data_valid,
  init_calib => NN_1,
  rd_data(63 downto 0) => rd_data(63 downto 0),
  O_psram_ck(1 downto 0) => O_psram_ck(1 downto 0),
  O_psram_ck_n(1 downto 0) => O_psram_ck_n(1 downto 0),
  O_psram_cs_n(1 downto 0) => O_psram_cs_n(1 downto 0),
  O_psram_reset_n(1) => NN,
  IO_psram_dq(15 downto 0) => IO_psram_dq(15 downto 0),
  IO_psram_rwds(1 downto 0) => IO_psram_rwds(1 downto 0));
  O_psram_reset_n(0) <= NN;
  O_psram_reset_n(1) <= NN;
  clk_out <= NN_0;
  init_calib <= NN_1;
end beh;
